magic
tech sky130A
magscale 1 2
timestamp 1629190088
<< nwell >>
rect 40625 13166 43821 17512
rect 39137 10778 51261 12888
rect 39137 6977 51261 9087
rect 40625 2353 43821 6699
<< pwell >>
rect 40625 17860 49773 19734
rect 45789 15322 46191 16618
rect 39339 4710 40059 6906
rect 44495 4070 45215 6266
rect 45789 3247 46191 4543
rect 40625 131 49773 2005
<< pmoslvt >>
rect 40821 16493 41021 17293
rect 41193 16493 41393 17293
rect 41565 16493 41765 17293
rect 41937 16493 42137 17293
rect 42309 16493 42509 17293
rect 42681 16493 42881 17293
rect 43053 16493 43253 17293
rect 43425 16493 43625 17293
rect 40821 15457 41021 16257
rect 41193 15457 41393 16257
rect 41565 15457 41765 16257
rect 41937 15457 42137 16257
rect 42309 15457 42509 16257
rect 42681 15457 42881 16257
rect 43053 15457 43253 16257
rect 43425 15457 43625 16257
rect 40821 14421 41021 15221
rect 41193 14421 41393 15221
rect 41565 14421 41765 15221
rect 41937 14421 42137 15221
rect 42309 14421 42509 15221
rect 42681 14421 42881 15221
rect 43053 14421 43253 15221
rect 43425 14421 43625 15221
rect 40821 13385 41021 14185
rect 41193 13385 41393 14185
rect 41565 13385 41765 14185
rect 41937 13385 42137 14185
rect 42309 13385 42509 14185
rect 42681 13385 42881 14185
rect 43053 13385 43253 14185
rect 43425 13385 43625 14185
rect 39333 12269 39533 12669
rect 39705 12269 39905 12669
rect 40077 12269 40277 12669
rect 40449 12269 40649 12669
rect 40821 12269 41021 12669
rect 41193 12269 41393 12669
rect 41565 12269 41765 12669
rect 41937 12269 42137 12669
rect 42309 12269 42509 12669
rect 42681 12269 42881 12669
rect 43053 12269 43253 12669
rect 43425 12269 43625 12669
rect 43797 12269 43997 12669
rect 44169 12269 44369 12669
rect 44541 12269 44741 12669
rect 44913 12269 45113 12669
rect 45285 12269 45485 12669
rect 45657 12269 45857 12669
rect 46029 12269 46229 12669
rect 46401 12269 46601 12669
rect 46773 12269 46973 12669
rect 47145 12269 47345 12669
rect 47517 12269 47717 12669
rect 47889 12269 48089 12669
rect 48261 12269 48461 12669
rect 48633 12269 48833 12669
rect 49005 12269 49205 12669
rect 49377 12269 49577 12669
rect 49749 12269 49949 12669
rect 50121 12269 50321 12669
rect 50493 12269 50693 12669
rect 50865 12269 51065 12669
rect 39333 11633 39533 12033
rect 39705 11633 39905 12033
rect 40077 11633 40277 12033
rect 40449 11633 40649 12033
rect 40821 11633 41021 12033
rect 41193 11633 41393 12033
rect 41565 11633 41765 12033
rect 41937 11633 42137 12033
rect 42309 11633 42509 12033
rect 42681 11633 42881 12033
rect 43053 11633 43253 12033
rect 43425 11633 43625 12033
rect 43797 11633 43997 12033
rect 44169 11633 44369 12033
rect 44541 11633 44741 12033
rect 44913 11633 45113 12033
rect 45285 11633 45485 12033
rect 45657 11633 45857 12033
rect 46029 11633 46229 12033
rect 46401 11633 46601 12033
rect 46773 11633 46973 12033
rect 47145 11633 47345 12033
rect 47517 11633 47717 12033
rect 47889 11633 48089 12033
rect 48261 11633 48461 12033
rect 48633 11633 48833 12033
rect 49005 11633 49205 12033
rect 49377 11633 49577 12033
rect 49749 11633 49949 12033
rect 50121 11633 50321 12033
rect 50493 11633 50693 12033
rect 50865 11633 51065 12033
rect 39333 10997 39533 11397
rect 39705 10997 39905 11397
rect 40077 10997 40277 11397
rect 40449 10997 40649 11397
rect 40821 10997 41021 11397
rect 41193 10997 41393 11397
rect 41565 10997 41765 11397
rect 41937 10997 42137 11397
rect 42309 10997 42509 11397
rect 42681 10997 42881 11397
rect 43053 10997 43253 11397
rect 43425 10997 43625 11397
rect 43797 10997 43997 11397
rect 44169 10997 44369 11397
rect 44541 10997 44741 11397
rect 44913 10997 45113 11397
rect 45285 10997 45485 11397
rect 45657 10997 45857 11397
rect 46029 10997 46229 11397
rect 46401 10997 46601 11397
rect 46773 10997 46973 11397
rect 47145 10997 47345 11397
rect 47517 10997 47717 11397
rect 47889 10997 48089 11397
rect 48261 10997 48461 11397
rect 48633 10997 48833 11397
rect 49005 10997 49205 11397
rect 49377 10997 49577 11397
rect 49749 10997 49949 11397
rect 50121 10997 50321 11397
rect 50493 10997 50693 11397
rect 50865 10997 51065 11397
rect 39333 8468 39533 8868
rect 39705 8468 39905 8868
rect 40077 8468 40277 8868
rect 40449 8468 40649 8868
rect 40821 8468 41021 8868
rect 41193 8468 41393 8868
rect 41565 8468 41765 8868
rect 41937 8468 42137 8868
rect 42309 8468 42509 8868
rect 42681 8468 42881 8868
rect 43053 8468 43253 8868
rect 43425 8468 43625 8868
rect 43797 8468 43997 8868
rect 44169 8468 44369 8868
rect 44541 8468 44741 8868
rect 44913 8468 45113 8868
rect 45285 8468 45485 8868
rect 45657 8468 45857 8868
rect 46029 8468 46229 8868
rect 46401 8468 46601 8868
rect 46773 8468 46973 8868
rect 47145 8468 47345 8868
rect 47517 8468 47717 8868
rect 47889 8468 48089 8868
rect 48261 8468 48461 8868
rect 48633 8468 48833 8868
rect 49005 8468 49205 8868
rect 49377 8468 49577 8868
rect 49749 8468 49949 8868
rect 50121 8468 50321 8868
rect 50493 8468 50693 8868
rect 50865 8468 51065 8868
rect 39333 7832 39533 8232
rect 39705 7832 39905 8232
rect 40077 7832 40277 8232
rect 40449 7832 40649 8232
rect 40821 7832 41021 8232
rect 41193 7832 41393 8232
rect 41565 7832 41765 8232
rect 41937 7832 42137 8232
rect 42309 7832 42509 8232
rect 42681 7832 42881 8232
rect 43053 7832 43253 8232
rect 43425 7832 43625 8232
rect 43797 7832 43997 8232
rect 44169 7832 44369 8232
rect 44541 7832 44741 8232
rect 44913 7832 45113 8232
rect 45285 7832 45485 8232
rect 45657 7832 45857 8232
rect 46029 7832 46229 8232
rect 46401 7832 46601 8232
rect 46773 7832 46973 8232
rect 47145 7832 47345 8232
rect 47517 7832 47717 8232
rect 47889 7832 48089 8232
rect 48261 7832 48461 8232
rect 48633 7832 48833 8232
rect 49005 7832 49205 8232
rect 49377 7832 49577 8232
rect 49749 7832 49949 8232
rect 50121 7832 50321 8232
rect 50493 7832 50693 8232
rect 50865 7832 51065 8232
rect 39333 7196 39533 7596
rect 39705 7196 39905 7596
rect 40077 7196 40277 7596
rect 40449 7196 40649 7596
rect 40821 7196 41021 7596
rect 41193 7196 41393 7596
rect 41565 7196 41765 7596
rect 41937 7196 42137 7596
rect 42309 7196 42509 7596
rect 42681 7196 42881 7596
rect 43053 7196 43253 7596
rect 43425 7196 43625 7596
rect 43797 7196 43997 7596
rect 44169 7196 44369 7596
rect 44541 7196 44741 7596
rect 44913 7196 45113 7596
rect 45285 7196 45485 7596
rect 45657 7196 45857 7596
rect 46029 7196 46229 7596
rect 46401 7196 46601 7596
rect 46773 7196 46973 7596
rect 47145 7196 47345 7596
rect 47517 7196 47717 7596
rect 47889 7196 48089 7596
rect 48261 7196 48461 7596
rect 48633 7196 48833 7596
rect 49005 7196 49205 7596
rect 49377 7196 49577 7596
rect 49749 7196 49949 7596
rect 50121 7196 50321 7596
rect 50493 7196 50693 7596
rect 50865 7196 51065 7596
rect 40821 5680 41021 6480
rect 41193 5680 41393 6480
rect 41565 5680 41765 6480
rect 41937 5680 42137 6480
rect 42309 5680 42509 6480
rect 42681 5680 42881 6480
rect 43053 5680 43253 6480
rect 43425 5680 43625 6480
rect 40821 4644 41021 5444
rect 41193 4644 41393 5444
rect 41565 4644 41765 5444
rect 41937 4644 42137 5444
rect 42309 4644 42509 5444
rect 42681 4644 42881 5444
rect 43053 4644 43253 5444
rect 43425 4644 43625 5444
rect 40821 3608 41021 4408
rect 41193 3608 41393 4408
rect 41565 3608 41765 4408
rect 41937 3608 42137 4408
rect 42309 3608 42509 4408
rect 42681 3608 42881 4408
rect 43053 3608 43253 4408
rect 43425 3608 43625 4408
rect 40821 2572 41021 3372
rect 41193 2572 41393 3372
rect 41565 2572 41765 3372
rect 41937 2572 42137 3372
rect 42309 2572 42509 3372
rect 42681 2572 42881 3372
rect 43053 2572 43253 3372
rect 43425 2572 43625 3372
<< nmoslvt >>
rect 40821 19324 41021 19524
rect 41193 19324 41393 19524
rect 41565 19324 41765 19524
rect 41937 19324 42137 19524
rect 42309 19324 42509 19524
rect 42681 19324 42881 19524
rect 43053 19324 43253 19524
rect 43425 19324 43625 19524
rect 43797 19324 43997 19524
rect 44169 19324 44369 19524
rect 44541 19324 44741 19524
rect 44913 19324 45113 19524
rect 45285 19324 45485 19524
rect 45657 19324 45857 19524
rect 46029 19324 46229 19524
rect 46401 19324 46601 19524
rect 46773 19324 46973 19524
rect 47145 19324 47345 19524
rect 47517 19324 47717 19524
rect 47889 19324 48089 19524
rect 48261 19324 48461 19524
rect 48633 19324 48833 19524
rect 49005 19324 49205 19524
rect 49377 19324 49577 19524
rect 40821 18906 41021 19106
rect 41193 18906 41393 19106
rect 41565 18906 41765 19106
rect 41937 18906 42137 19106
rect 42309 18906 42509 19106
rect 42681 18906 42881 19106
rect 43053 18906 43253 19106
rect 43425 18906 43625 19106
rect 43797 18906 43997 19106
rect 44169 18906 44369 19106
rect 44541 18906 44741 19106
rect 44913 18906 45113 19106
rect 45285 18906 45485 19106
rect 45657 18906 45857 19106
rect 46029 18906 46229 19106
rect 46401 18906 46601 19106
rect 46773 18906 46973 19106
rect 47145 18906 47345 19106
rect 47517 18906 47717 19106
rect 47889 18906 48089 19106
rect 48261 18906 48461 19106
rect 48633 18906 48833 19106
rect 49005 18906 49205 19106
rect 49377 18906 49577 19106
rect 40821 18488 41021 18688
rect 41193 18488 41393 18688
rect 41565 18488 41765 18688
rect 41937 18488 42137 18688
rect 42309 18488 42509 18688
rect 42681 18488 42881 18688
rect 43053 18488 43253 18688
rect 43425 18488 43625 18688
rect 43797 18488 43997 18688
rect 44169 18488 44369 18688
rect 44541 18488 44741 18688
rect 44913 18488 45113 18688
rect 45285 18488 45485 18688
rect 45657 18488 45857 18688
rect 46029 18488 46229 18688
rect 46401 18488 46601 18688
rect 46773 18488 46973 18688
rect 47145 18488 47345 18688
rect 47517 18488 47717 18688
rect 47889 18488 48089 18688
rect 48261 18488 48461 18688
rect 48633 18488 48833 18688
rect 49005 18488 49205 18688
rect 49377 18488 49577 18688
rect 40821 18070 41021 18270
rect 41193 18070 41393 18270
rect 41565 18070 41765 18270
rect 41937 18070 42137 18270
rect 42309 18070 42509 18270
rect 42681 18070 42881 18270
rect 43053 18070 43253 18270
rect 43425 18070 43625 18270
rect 43797 18070 43997 18270
rect 44169 18070 44369 18270
rect 44541 18070 44741 18270
rect 44913 18070 45113 18270
rect 45285 18070 45485 18270
rect 45657 18070 45857 18270
rect 46029 18070 46229 18270
rect 46401 18070 46601 18270
rect 46773 18070 46973 18270
rect 47145 18070 47345 18270
rect 47517 18070 47717 18270
rect 47889 18070 48089 18270
rect 48261 18070 48461 18270
rect 48633 18070 48833 18270
rect 49005 18070 49205 18270
rect 49377 18070 49577 18270
rect 40821 1595 41021 1795
rect 41193 1595 41393 1795
rect 41565 1595 41765 1795
rect 41937 1595 42137 1795
rect 42309 1595 42509 1795
rect 42681 1595 42881 1795
rect 43053 1595 43253 1795
rect 43425 1595 43625 1795
rect 43797 1595 43997 1795
rect 44169 1595 44369 1795
rect 44541 1595 44741 1795
rect 44913 1595 45113 1795
rect 45285 1595 45485 1795
rect 45657 1595 45857 1795
rect 46029 1595 46229 1795
rect 46401 1595 46601 1795
rect 46773 1595 46973 1795
rect 47145 1595 47345 1795
rect 47517 1595 47717 1795
rect 47889 1595 48089 1795
rect 48261 1595 48461 1795
rect 48633 1595 48833 1795
rect 49005 1595 49205 1795
rect 49377 1595 49577 1795
rect 40821 1177 41021 1377
rect 41193 1177 41393 1377
rect 41565 1177 41765 1377
rect 41937 1177 42137 1377
rect 42309 1177 42509 1377
rect 42681 1177 42881 1377
rect 43053 1177 43253 1377
rect 43425 1177 43625 1377
rect 43797 1177 43997 1377
rect 44169 1177 44369 1377
rect 44541 1177 44741 1377
rect 44913 1177 45113 1377
rect 45285 1177 45485 1377
rect 45657 1177 45857 1377
rect 46029 1177 46229 1377
rect 46401 1177 46601 1377
rect 46773 1177 46973 1377
rect 47145 1177 47345 1377
rect 47517 1177 47717 1377
rect 47889 1177 48089 1377
rect 48261 1177 48461 1377
rect 48633 1177 48833 1377
rect 49005 1177 49205 1377
rect 49377 1177 49577 1377
rect 40821 759 41021 959
rect 41193 759 41393 959
rect 41565 759 41765 959
rect 41937 759 42137 959
rect 42309 759 42509 959
rect 42681 759 42881 959
rect 43053 759 43253 959
rect 43425 759 43625 959
rect 43797 759 43997 959
rect 44169 759 44369 959
rect 44541 759 44741 959
rect 44913 759 45113 959
rect 45285 759 45485 959
rect 45657 759 45857 959
rect 46029 759 46229 959
rect 46401 759 46601 959
rect 46773 759 46973 959
rect 47145 759 47345 959
rect 47517 759 47717 959
rect 47889 759 48089 959
rect 48261 759 48461 959
rect 48633 759 48833 959
rect 49005 759 49205 959
rect 49377 759 49577 959
rect 40821 341 41021 541
rect 41193 341 41393 541
rect 41565 341 41765 541
rect 41937 341 42137 541
rect 42309 341 42509 541
rect 42681 341 42881 541
rect 43053 341 43253 541
rect 43425 341 43625 541
rect 43797 341 43997 541
rect 44169 341 44369 541
rect 44541 341 44741 541
rect 44913 341 45113 541
rect 45285 341 45485 541
rect 45657 341 45857 541
rect 46029 341 46229 541
rect 46401 341 46601 541
rect 46773 341 46973 541
rect 47145 341 47345 541
rect 47517 341 47717 541
rect 47889 341 48089 541
rect 48261 341 48461 541
rect 48633 341 48833 541
rect 49005 341 49205 541
rect 49377 341 49577 541
<< ndiff >>
rect 40763 19512 40821 19524
rect 40763 19336 40775 19512
rect 40809 19336 40821 19512
rect 40763 19324 40821 19336
rect 41021 19512 41079 19524
rect 41021 19336 41033 19512
rect 41067 19336 41079 19512
rect 41021 19324 41079 19336
rect 41135 19512 41193 19524
rect 41135 19336 41147 19512
rect 41181 19336 41193 19512
rect 41135 19324 41193 19336
rect 41393 19512 41451 19524
rect 41393 19336 41405 19512
rect 41439 19336 41451 19512
rect 41393 19324 41451 19336
rect 41507 19512 41565 19524
rect 41507 19336 41519 19512
rect 41553 19336 41565 19512
rect 41507 19324 41565 19336
rect 41765 19512 41823 19524
rect 41765 19336 41777 19512
rect 41811 19336 41823 19512
rect 41765 19324 41823 19336
rect 41879 19512 41937 19524
rect 41879 19336 41891 19512
rect 41925 19336 41937 19512
rect 41879 19324 41937 19336
rect 42137 19512 42195 19524
rect 42137 19336 42149 19512
rect 42183 19336 42195 19512
rect 42137 19324 42195 19336
rect 42251 19512 42309 19524
rect 42251 19336 42263 19512
rect 42297 19336 42309 19512
rect 42251 19324 42309 19336
rect 42509 19512 42567 19524
rect 42509 19336 42521 19512
rect 42555 19336 42567 19512
rect 42509 19324 42567 19336
rect 42623 19512 42681 19524
rect 42623 19336 42635 19512
rect 42669 19336 42681 19512
rect 42623 19324 42681 19336
rect 42881 19512 42939 19524
rect 42881 19336 42893 19512
rect 42927 19336 42939 19512
rect 42881 19324 42939 19336
rect 42995 19512 43053 19524
rect 42995 19336 43007 19512
rect 43041 19336 43053 19512
rect 42995 19324 43053 19336
rect 43253 19512 43311 19524
rect 43253 19336 43265 19512
rect 43299 19336 43311 19512
rect 43253 19324 43311 19336
rect 43367 19512 43425 19524
rect 43367 19336 43379 19512
rect 43413 19336 43425 19512
rect 43367 19324 43425 19336
rect 43625 19512 43683 19524
rect 43625 19336 43637 19512
rect 43671 19336 43683 19512
rect 43625 19324 43683 19336
rect 43739 19512 43797 19524
rect 43739 19336 43751 19512
rect 43785 19336 43797 19512
rect 43739 19324 43797 19336
rect 43997 19512 44055 19524
rect 43997 19336 44009 19512
rect 44043 19336 44055 19512
rect 43997 19324 44055 19336
rect 44111 19512 44169 19524
rect 44111 19336 44123 19512
rect 44157 19336 44169 19512
rect 44111 19324 44169 19336
rect 44369 19512 44427 19524
rect 44369 19336 44381 19512
rect 44415 19336 44427 19512
rect 44369 19324 44427 19336
rect 44483 19512 44541 19524
rect 44483 19336 44495 19512
rect 44529 19336 44541 19512
rect 44483 19324 44541 19336
rect 44741 19512 44799 19524
rect 44741 19336 44753 19512
rect 44787 19336 44799 19512
rect 44741 19324 44799 19336
rect 44855 19512 44913 19524
rect 44855 19336 44867 19512
rect 44901 19336 44913 19512
rect 44855 19324 44913 19336
rect 45113 19512 45171 19524
rect 45113 19336 45125 19512
rect 45159 19336 45171 19512
rect 45113 19324 45171 19336
rect 45227 19512 45285 19524
rect 45227 19336 45239 19512
rect 45273 19336 45285 19512
rect 45227 19324 45285 19336
rect 45485 19512 45543 19524
rect 45485 19336 45497 19512
rect 45531 19336 45543 19512
rect 45485 19324 45543 19336
rect 45599 19512 45657 19524
rect 45599 19336 45611 19512
rect 45645 19336 45657 19512
rect 45599 19324 45657 19336
rect 45857 19512 45915 19524
rect 45857 19336 45869 19512
rect 45903 19336 45915 19512
rect 45857 19324 45915 19336
rect 45971 19512 46029 19524
rect 45971 19336 45983 19512
rect 46017 19336 46029 19512
rect 45971 19324 46029 19336
rect 46229 19512 46287 19524
rect 46229 19336 46241 19512
rect 46275 19336 46287 19512
rect 46229 19324 46287 19336
rect 46343 19512 46401 19524
rect 46343 19336 46355 19512
rect 46389 19336 46401 19512
rect 46343 19324 46401 19336
rect 46601 19512 46659 19524
rect 46601 19336 46613 19512
rect 46647 19336 46659 19512
rect 46601 19324 46659 19336
rect 46715 19512 46773 19524
rect 46715 19336 46727 19512
rect 46761 19336 46773 19512
rect 46715 19324 46773 19336
rect 46973 19512 47031 19524
rect 46973 19336 46985 19512
rect 47019 19336 47031 19512
rect 46973 19324 47031 19336
rect 47087 19512 47145 19524
rect 47087 19336 47099 19512
rect 47133 19336 47145 19512
rect 47087 19324 47145 19336
rect 47345 19512 47403 19524
rect 47345 19336 47357 19512
rect 47391 19336 47403 19512
rect 47345 19324 47403 19336
rect 47459 19512 47517 19524
rect 47459 19336 47471 19512
rect 47505 19336 47517 19512
rect 47459 19324 47517 19336
rect 47717 19512 47775 19524
rect 47717 19336 47729 19512
rect 47763 19336 47775 19512
rect 47717 19324 47775 19336
rect 47831 19512 47889 19524
rect 47831 19336 47843 19512
rect 47877 19336 47889 19512
rect 47831 19324 47889 19336
rect 48089 19512 48147 19524
rect 48089 19336 48101 19512
rect 48135 19336 48147 19512
rect 48089 19324 48147 19336
rect 48203 19512 48261 19524
rect 48203 19336 48215 19512
rect 48249 19336 48261 19512
rect 48203 19324 48261 19336
rect 48461 19512 48519 19524
rect 48461 19336 48473 19512
rect 48507 19336 48519 19512
rect 48461 19324 48519 19336
rect 48575 19512 48633 19524
rect 48575 19336 48587 19512
rect 48621 19336 48633 19512
rect 48575 19324 48633 19336
rect 48833 19512 48891 19524
rect 48833 19336 48845 19512
rect 48879 19336 48891 19512
rect 48833 19324 48891 19336
rect 48947 19512 49005 19524
rect 48947 19336 48959 19512
rect 48993 19336 49005 19512
rect 48947 19324 49005 19336
rect 49205 19512 49263 19524
rect 49205 19336 49217 19512
rect 49251 19336 49263 19512
rect 49205 19324 49263 19336
rect 49319 19512 49377 19524
rect 49319 19336 49331 19512
rect 49365 19336 49377 19512
rect 49319 19324 49377 19336
rect 49577 19512 49635 19524
rect 49577 19336 49589 19512
rect 49623 19336 49635 19512
rect 49577 19324 49635 19336
rect 40763 19094 40821 19106
rect 40763 18918 40775 19094
rect 40809 18918 40821 19094
rect 40763 18906 40821 18918
rect 41021 19094 41079 19106
rect 41021 18918 41033 19094
rect 41067 18918 41079 19094
rect 41021 18906 41079 18918
rect 41135 19094 41193 19106
rect 41135 18918 41147 19094
rect 41181 18918 41193 19094
rect 41135 18906 41193 18918
rect 41393 19094 41451 19106
rect 41393 18918 41405 19094
rect 41439 18918 41451 19094
rect 41393 18906 41451 18918
rect 41507 19094 41565 19106
rect 41507 18918 41519 19094
rect 41553 18918 41565 19094
rect 41507 18906 41565 18918
rect 41765 19094 41823 19106
rect 41765 18918 41777 19094
rect 41811 18918 41823 19094
rect 41765 18906 41823 18918
rect 41879 19094 41937 19106
rect 41879 18918 41891 19094
rect 41925 18918 41937 19094
rect 41879 18906 41937 18918
rect 42137 19094 42195 19106
rect 42137 18918 42149 19094
rect 42183 18918 42195 19094
rect 42137 18906 42195 18918
rect 42251 19094 42309 19106
rect 42251 18918 42263 19094
rect 42297 18918 42309 19094
rect 42251 18906 42309 18918
rect 42509 19094 42567 19106
rect 42509 18918 42521 19094
rect 42555 18918 42567 19094
rect 42509 18906 42567 18918
rect 42623 19094 42681 19106
rect 42623 18918 42635 19094
rect 42669 18918 42681 19094
rect 42623 18906 42681 18918
rect 42881 19094 42939 19106
rect 42881 18918 42893 19094
rect 42927 18918 42939 19094
rect 42881 18906 42939 18918
rect 42995 19094 43053 19106
rect 42995 18918 43007 19094
rect 43041 18918 43053 19094
rect 42995 18906 43053 18918
rect 43253 19094 43311 19106
rect 43253 18918 43265 19094
rect 43299 18918 43311 19094
rect 43253 18906 43311 18918
rect 43367 19094 43425 19106
rect 43367 18918 43379 19094
rect 43413 18918 43425 19094
rect 43367 18906 43425 18918
rect 43625 19094 43683 19106
rect 43625 18918 43637 19094
rect 43671 18918 43683 19094
rect 43625 18906 43683 18918
rect 43739 19094 43797 19106
rect 43739 18918 43751 19094
rect 43785 18918 43797 19094
rect 43739 18906 43797 18918
rect 43997 19094 44055 19106
rect 43997 18918 44009 19094
rect 44043 18918 44055 19094
rect 43997 18906 44055 18918
rect 44111 19094 44169 19106
rect 44111 18918 44123 19094
rect 44157 18918 44169 19094
rect 44111 18906 44169 18918
rect 44369 19094 44427 19106
rect 44369 18918 44381 19094
rect 44415 18918 44427 19094
rect 44369 18906 44427 18918
rect 44483 19094 44541 19106
rect 44483 18918 44495 19094
rect 44529 18918 44541 19094
rect 44483 18906 44541 18918
rect 44741 19094 44799 19106
rect 44741 18918 44753 19094
rect 44787 18918 44799 19094
rect 44741 18906 44799 18918
rect 44855 19094 44913 19106
rect 44855 18918 44867 19094
rect 44901 18918 44913 19094
rect 44855 18906 44913 18918
rect 45113 19094 45171 19106
rect 45113 18918 45125 19094
rect 45159 18918 45171 19094
rect 45113 18906 45171 18918
rect 45227 19094 45285 19106
rect 45227 18918 45239 19094
rect 45273 18918 45285 19094
rect 45227 18906 45285 18918
rect 45485 19094 45543 19106
rect 45485 18918 45497 19094
rect 45531 18918 45543 19094
rect 45485 18906 45543 18918
rect 45599 19094 45657 19106
rect 45599 18918 45611 19094
rect 45645 18918 45657 19094
rect 45599 18906 45657 18918
rect 45857 19094 45915 19106
rect 45857 18918 45869 19094
rect 45903 18918 45915 19094
rect 45857 18906 45915 18918
rect 45971 19094 46029 19106
rect 45971 18918 45983 19094
rect 46017 18918 46029 19094
rect 45971 18906 46029 18918
rect 46229 19094 46287 19106
rect 46229 18918 46241 19094
rect 46275 18918 46287 19094
rect 46229 18906 46287 18918
rect 46343 19094 46401 19106
rect 46343 18918 46355 19094
rect 46389 18918 46401 19094
rect 46343 18906 46401 18918
rect 46601 19094 46659 19106
rect 46601 18918 46613 19094
rect 46647 18918 46659 19094
rect 46601 18906 46659 18918
rect 46715 19094 46773 19106
rect 46715 18918 46727 19094
rect 46761 18918 46773 19094
rect 46715 18906 46773 18918
rect 46973 19094 47031 19106
rect 46973 18918 46985 19094
rect 47019 18918 47031 19094
rect 46973 18906 47031 18918
rect 47087 19094 47145 19106
rect 47087 18918 47099 19094
rect 47133 18918 47145 19094
rect 47087 18906 47145 18918
rect 47345 19094 47403 19106
rect 47345 18918 47357 19094
rect 47391 18918 47403 19094
rect 47345 18906 47403 18918
rect 47459 19094 47517 19106
rect 47459 18918 47471 19094
rect 47505 18918 47517 19094
rect 47459 18906 47517 18918
rect 47717 19094 47775 19106
rect 47717 18918 47729 19094
rect 47763 18918 47775 19094
rect 47717 18906 47775 18918
rect 47831 19094 47889 19106
rect 47831 18918 47843 19094
rect 47877 18918 47889 19094
rect 47831 18906 47889 18918
rect 48089 19094 48147 19106
rect 48089 18918 48101 19094
rect 48135 18918 48147 19094
rect 48089 18906 48147 18918
rect 48203 19094 48261 19106
rect 48203 18918 48215 19094
rect 48249 18918 48261 19094
rect 48203 18906 48261 18918
rect 48461 19094 48519 19106
rect 48461 18918 48473 19094
rect 48507 18918 48519 19094
rect 48461 18906 48519 18918
rect 48575 19094 48633 19106
rect 48575 18918 48587 19094
rect 48621 18918 48633 19094
rect 48575 18906 48633 18918
rect 48833 19094 48891 19106
rect 48833 18918 48845 19094
rect 48879 18918 48891 19094
rect 48833 18906 48891 18918
rect 48947 19094 49005 19106
rect 48947 18918 48959 19094
rect 48993 18918 49005 19094
rect 48947 18906 49005 18918
rect 49205 19094 49263 19106
rect 49205 18918 49217 19094
rect 49251 18918 49263 19094
rect 49205 18906 49263 18918
rect 49319 19094 49377 19106
rect 49319 18918 49331 19094
rect 49365 18918 49377 19094
rect 49319 18906 49377 18918
rect 49577 19094 49635 19106
rect 49577 18918 49589 19094
rect 49623 18918 49635 19094
rect 49577 18906 49635 18918
rect 40763 18676 40821 18688
rect 40763 18500 40775 18676
rect 40809 18500 40821 18676
rect 40763 18488 40821 18500
rect 41021 18676 41079 18688
rect 41021 18500 41033 18676
rect 41067 18500 41079 18676
rect 41021 18488 41079 18500
rect 41135 18676 41193 18688
rect 41135 18500 41147 18676
rect 41181 18500 41193 18676
rect 41135 18488 41193 18500
rect 41393 18676 41451 18688
rect 41393 18500 41405 18676
rect 41439 18500 41451 18676
rect 41393 18488 41451 18500
rect 41507 18676 41565 18688
rect 41507 18500 41519 18676
rect 41553 18500 41565 18676
rect 41507 18488 41565 18500
rect 41765 18676 41823 18688
rect 41765 18500 41777 18676
rect 41811 18500 41823 18676
rect 41765 18488 41823 18500
rect 41879 18676 41937 18688
rect 41879 18500 41891 18676
rect 41925 18500 41937 18676
rect 41879 18488 41937 18500
rect 42137 18676 42195 18688
rect 42137 18500 42149 18676
rect 42183 18500 42195 18676
rect 42137 18488 42195 18500
rect 42251 18676 42309 18688
rect 42251 18500 42263 18676
rect 42297 18500 42309 18676
rect 42251 18488 42309 18500
rect 42509 18676 42567 18688
rect 42509 18500 42521 18676
rect 42555 18500 42567 18676
rect 42509 18488 42567 18500
rect 42623 18676 42681 18688
rect 42623 18500 42635 18676
rect 42669 18500 42681 18676
rect 42623 18488 42681 18500
rect 42881 18676 42939 18688
rect 42881 18500 42893 18676
rect 42927 18500 42939 18676
rect 42881 18488 42939 18500
rect 42995 18676 43053 18688
rect 42995 18500 43007 18676
rect 43041 18500 43053 18676
rect 42995 18488 43053 18500
rect 43253 18676 43311 18688
rect 43253 18500 43265 18676
rect 43299 18500 43311 18676
rect 43253 18488 43311 18500
rect 43367 18676 43425 18688
rect 43367 18500 43379 18676
rect 43413 18500 43425 18676
rect 43367 18488 43425 18500
rect 43625 18676 43683 18688
rect 43625 18500 43637 18676
rect 43671 18500 43683 18676
rect 43625 18488 43683 18500
rect 43739 18676 43797 18688
rect 43739 18500 43751 18676
rect 43785 18500 43797 18676
rect 43739 18488 43797 18500
rect 43997 18676 44055 18688
rect 43997 18500 44009 18676
rect 44043 18500 44055 18676
rect 43997 18488 44055 18500
rect 44111 18676 44169 18688
rect 44111 18500 44123 18676
rect 44157 18500 44169 18676
rect 44111 18488 44169 18500
rect 44369 18676 44427 18688
rect 44369 18500 44381 18676
rect 44415 18500 44427 18676
rect 44369 18488 44427 18500
rect 44483 18676 44541 18688
rect 44483 18500 44495 18676
rect 44529 18500 44541 18676
rect 44483 18488 44541 18500
rect 44741 18676 44799 18688
rect 44741 18500 44753 18676
rect 44787 18500 44799 18676
rect 44741 18488 44799 18500
rect 44855 18676 44913 18688
rect 44855 18500 44867 18676
rect 44901 18500 44913 18676
rect 44855 18488 44913 18500
rect 45113 18676 45171 18688
rect 45113 18500 45125 18676
rect 45159 18500 45171 18676
rect 45113 18488 45171 18500
rect 45227 18676 45285 18688
rect 45227 18500 45239 18676
rect 45273 18500 45285 18676
rect 45227 18488 45285 18500
rect 45485 18676 45543 18688
rect 45485 18500 45497 18676
rect 45531 18500 45543 18676
rect 45485 18488 45543 18500
rect 45599 18676 45657 18688
rect 45599 18500 45611 18676
rect 45645 18500 45657 18676
rect 45599 18488 45657 18500
rect 45857 18676 45915 18688
rect 45857 18500 45869 18676
rect 45903 18500 45915 18676
rect 45857 18488 45915 18500
rect 45971 18676 46029 18688
rect 45971 18500 45983 18676
rect 46017 18500 46029 18676
rect 45971 18488 46029 18500
rect 46229 18676 46287 18688
rect 46229 18500 46241 18676
rect 46275 18500 46287 18676
rect 46229 18488 46287 18500
rect 46343 18676 46401 18688
rect 46343 18500 46355 18676
rect 46389 18500 46401 18676
rect 46343 18488 46401 18500
rect 46601 18676 46659 18688
rect 46601 18500 46613 18676
rect 46647 18500 46659 18676
rect 46601 18488 46659 18500
rect 46715 18676 46773 18688
rect 46715 18500 46727 18676
rect 46761 18500 46773 18676
rect 46715 18488 46773 18500
rect 46973 18676 47031 18688
rect 46973 18500 46985 18676
rect 47019 18500 47031 18676
rect 46973 18488 47031 18500
rect 47087 18676 47145 18688
rect 47087 18500 47099 18676
rect 47133 18500 47145 18676
rect 47087 18488 47145 18500
rect 47345 18676 47403 18688
rect 47345 18500 47357 18676
rect 47391 18500 47403 18676
rect 47345 18488 47403 18500
rect 47459 18676 47517 18688
rect 47459 18500 47471 18676
rect 47505 18500 47517 18676
rect 47459 18488 47517 18500
rect 47717 18676 47775 18688
rect 47717 18500 47729 18676
rect 47763 18500 47775 18676
rect 47717 18488 47775 18500
rect 47831 18676 47889 18688
rect 47831 18500 47843 18676
rect 47877 18500 47889 18676
rect 47831 18488 47889 18500
rect 48089 18676 48147 18688
rect 48089 18500 48101 18676
rect 48135 18500 48147 18676
rect 48089 18488 48147 18500
rect 48203 18676 48261 18688
rect 48203 18500 48215 18676
rect 48249 18500 48261 18676
rect 48203 18488 48261 18500
rect 48461 18676 48519 18688
rect 48461 18500 48473 18676
rect 48507 18500 48519 18676
rect 48461 18488 48519 18500
rect 48575 18676 48633 18688
rect 48575 18500 48587 18676
rect 48621 18500 48633 18676
rect 48575 18488 48633 18500
rect 48833 18676 48891 18688
rect 48833 18500 48845 18676
rect 48879 18500 48891 18676
rect 48833 18488 48891 18500
rect 48947 18676 49005 18688
rect 48947 18500 48959 18676
rect 48993 18500 49005 18676
rect 48947 18488 49005 18500
rect 49205 18676 49263 18688
rect 49205 18500 49217 18676
rect 49251 18500 49263 18676
rect 49205 18488 49263 18500
rect 49319 18676 49377 18688
rect 49319 18500 49331 18676
rect 49365 18500 49377 18676
rect 49319 18488 49377 18500
rect 49577 18676 49635 18688
rect 49577 18500 49589 18676
rect 49623 18500 49635 18676
rect 49577 18488 49635 18500
rect 40763 18258 40821 18270
rect 40763 18082 40775 18258
rect 40809 18082 40821 18258
rect 40763 18070 40821 18082
rect 41021 18258 41079 18270
rect 41021 18082 41033 18258
rect 41067 18082 41079 18258
rect 41021 18070 41079 18082
rect 41135 18258 41193 18270
rect 41135 18082 41147 18258
rect 41181 18082 41193 18258
rect 41135 18070 41193 18082
rect 41393 18258 41451 18270
rect 41393 18082 41405 18258
rect 41439 18082 41451 18258
rect 41393 18070 41451 18082
rect 41507 18258 41565 18270
rect 41507 18082 41519 18258
rect 41553 18082 41565 18258
rect 41507 18070 41565 18082
rect 41765 18258 41823 18270
rect 41765 18082 41777 18258
rect 41811 18082 41823 18258
rect 41765 18070 41823 18082
rect 41879 18258 41937 18270
rect 41879 18082 41891 18258
rect 41925 18082 41937 18258
rect 41879 18070 41937 18082
rect 42137 18258 42195 18270
rect 42137 18082 42149 18258
rect 42183 18082 42195 18258
rect 42137 18070 42195 18082
rect 42251 18258 42309 18270
rect 42251 18082 42263 18258
rect 42297 18082 42309 18258
rect 42251 18070 42309 18082
rect 42509 18258 42567 18270
rect 42509 18082 42521 18258
rect 42555 18082 42567 18258
rect 42509 18070 42567 18082
rect 42623 18258 42681 18270
rect 42623 18082 42635 18258
rect 42669 18082 42681 18258
rect 42623 18070 42681 18082
rect 42881 18258 42939 18270
rect 42881 18082 42893 18258
rect 42927 18082 42939 18258
rect 42881 18070 42939 18082
rect 42995 18258 43053 18270
rect 42995 18082 43007 18258
rect 43041 18082 43053 18258
rect 42995 18070 43053 18082
rect 43253 18258 43311 18270
rect 43253 18082 43265 18258
rect 43299 18082 43311 18258
rect 43253 18070 43311 18082
rect 43367 18258 43425 18270
rect 43367 18082 43379 18258
rect 43413 18082 43425 18258
rect 43367 18070 43425 18082
rect 43625 18258 43683 18270
rect 43625 18082 43637 18258
rect 43671 18082 43683 18258
rect 43625 18070 43683 18082
rect 43739 18258 43797 18270
rect 43739 18082 43751 18258
rect 43785 18082 43797 18258
rect 43739 18070 43797 18082
rect 43997 18258 44055 18270
rect 43997 18082 44009 18258
rect 44043 18082 44055 18258
rect 43997 18070 44055 18082
rect 44111 18258 44169 18270
rect 44111 18082 44123 18258
rect 44157 18082 44169 18258
rect 44111 18070 44169 18082
rect 44369 18258 44427 18270
rect 44369 18082 44381 18258
rect 44415 18082 44427 18258
rect 44369 18070 44427 18082
rect 44483 18258 44541 18270
rect 44483 18082 44495 18258
rect 44529 18082 44541 18258
rect 44483 18070 44541 18082
rect 44741 18258 44799 18270
rect 44741 18082 44753 18258
rect 44787 18082 44799 18258
rect 44741 18070 44799 18082
rect 44855 18258 44913 18270
rect 44855 18082 44867 18258
rect 44901 18082 44913 18258
rect 44855 18070 44913 18082
rect 45113 18258 45171 18270
rect 45113 18082 45125 18258
rect 45159 18082 45171 18258
rect 45113 18070 45171 18082
rect 45227 18258 45285 18270
rect 45227 18082 45239 18258
rect 45273 18082 45285 18258
rect 45227 18070 45285 18082
rect 45485 18258 45543 18270
rect 45485 18082 45497 18258
rect 45531 18082 45543 18258
rect 45485 18070 45543 18082
rect 45599 18258 45657 18270
rect 45599 18082 45611 18258
rect 45645 18082 45657 18258
rect 45599 18070 45657 18082
rect 45857 18258 45915 18270
rect 45857 18082 45869 18258
rect 45903 18082 45915 18258
rect 45857 18070 45915 18082
rect 45971 18258 46029 18270
rect 45971 18082 45983 18258
rect 46017 18082 46029 18258
rect 45971 18070 46029 18082
rect 46229 18258 46287 18270
rect 46229 18082 46241 18258
rect 46275 18082 46287 18258
rect 46229 18070 46287 18082
rect 46343 18258 46401 18270
rect 46343 18082 46355 18258
rect 46389 18082 46401 18258
rect 46343 18070 46401 18082
rect 46601 18258 46659 18270
rect 46601 18082 46613 18258
rect 46647 18082 46659 18258
rect 46601 18070 46659 18082
rect 46715 18258 46773 18270
rect 46715 18082 46727 18258
rect 46761 18082 46773 18258
rect 46715 18070 46773 18082
rect 46973 18258 47031 18270
rect 46973 18082 46985 18258
rect 47019 18082 47031 18258
rect 46973 18070 47031 18082
rect 47087 18258 47145 18270
rect 47087 18082 47099 18258
rect 47133 18082 47145 18258
rect 47087 18070 47145 18082
rect 47345 18258 47403 18270
rect 47345 18082 47357 18258
rect 47391 18082 47403 18258
rect 47345 18070 47403 18082
rect 47459 18258 47517 18270
rect 47459 18082 47471 18258
rect 47505 18082 47517 18258
rect 47459 18070 47517 18082
rect 47717 18258 47775 18270
rect 47717 18082 47729 18258
rect 47763 18082 47775 18258
rect 47717 18070 47775 18082
rect 47831 18258 47889 18270
rect 47831 18082 47843 18258
rect 47877 18082 47889 18258
rect 47831 18070 47889 18082
rect 48089 18258 48147 18270
rect 48089 18082 48101 18258
rect 48135 18082 48147 18258
rect 48089 18070 48147 18082
rect 48203 18258 48261 18270
rect 48203 18082 48215 18258
rect 48249 18082 48261 18258
rect 48203 18070 48261 18082
rect 48461 18258 48519 18270
rect 48461 18082 48473 18258
rect 48507 18082 48519 18258
rect 48461 18070 48519 18082
rect 48575 18258 48633 18270
rect 48575 18082 48587 18258
rect 48621 18082 48633 18258
rect 48575 18070 48633 18082
rect 48833 18258 48891 18270
rect 48833 18082 48845 18258
rect 48879 18082 48891 18258
rect 48833 18070 48891 18082
rect 48947 18258 49005 18270
rect 48947 18082 48959 18258
rect 48993 18082 49005 18258
rect 48947 18070 49005 18082
rect 49205 18258 49263 18270
rect 49205 18082 49217 18258
rect 49251 18082 49263 18258
rect 49205 18070 49263 18082
rect 49319 18258 49377 18270
rect 49319 18082 49331 18258
rect 49365 18082 49377 18258
rect 49319 18070 49377 18082
rect 49577 18258 49635 18270
rect 49577 18082 49589 18258
rect 49623 18082 49635 18258
rect 49577 18070 49635 18082
rect 40763 1783 40821 1795
rect 40763 1607 40775 1783
rect 40809 1607 40821 1783
rect 40763 1595 40821 1607
rect 41021 1783 41079 1795
rect 41021 1607 41033 1783
rect 41067 1607 41079 1783
rect 41021 1595 41079 1607
rect 41135 1783 41193 1795
rect 41135 1607 41147 1783
rect 41181 1607 41193 1783
rect 41135 1595 41193 1607
rect 41393 1783 41451 1795
rect 41393 1607 41405 1783
rect 41439 1607 41451 1783
rect 41393 1595 41451 1607
rect 41507 1783 41565 1795
rect 41507 1607 41519 1783
rect 41553 1607 41565 1783
rect 41507 1595 41565 1607
rect 41765 1783 41823 1795
rect 41765 1607 41777 1783
rect 41811 1607 41823 1783
rect 41765 1595 41823 1607
rect 41879 1783 41937 1795
rect 41879 1607 41891 1783
rect 41925 1607 41937 1783
rect 41879 1595 41937 1607
rect 42137 1783 42195 1795
rect 42137 1607 42149 1783
rect 42183 1607 42195 1783
rect 42137 1595 42195 1607
rect 42251 1783 42309 1795
rect 42251 1607 42263 1783
rect 42297 1607 42309 1783
rect 42251 1595 42309 1607
rect 42509 1783 42567 1795
rect 42509 1607 42521 1783
rect 42555 1607 42567 1783
rect 42509 1595 42567 1607
rect 42623 1783 42681 1795
rect 42623 1607 42635 1783
rect 42669 1607 42681 1783
rect 42623 1595 42681 1607
rect 42881 1783 42939 1795
rect 42881 1607 42893 1783
rect 42927 1607 42939 1783
rect 42881 1595 42939 1607
rect 42995 1783 43053 1795
rect 42995 1607 43007 1783
rect 43041 1607 43053 1783
rect 42995 1595 43053 1607
rect 43253 1783 43311 1795
rect 43253 1607 43265 1783
rect 43299 1607 43311 1783
rect 43253 1595 43311 1607
rect 43367 1783 43425 1795
rect 43367 1607 43379 1783
rect 43413 1607 43425 1783
rect 43367 1595 43425 1607
rect 43625 1783 43683 1795
rect 43625 1607 43637 1783
rect 43671 1607 43683 1783
rect 43625 1595 43683 1607
rect 43739 1783 43797 1795
rect 43739 1607 43751 1783
rect 43785 1607 43797 1783
rect 43739 1595 43797 1607
rect 43997 1783 44055 1795
rect 43997 1607 44009 1783
rect 44043 1607 44055 1783
rect 43997 1595 44055 1607
rect 44111 1783 44169 1795
rect 44111 1607 44123 1783
rect 44157 1607 44169 1783
rect 44111 1595 44169 1607
rect 44369 1783 44427 1795
rect 44369 1607 44381 1783
rect 44415 1607 44427 1783
rect 44369 1595 44427 1607
rect 44483 1783 44541 1795
rect 44483 1607 44495 1783
rect 44529 1607 44541 1783
rect 44483 1595 44541 1607
rect 44741 1783 44799 1795
rect 44741 1607 44753 1783
rect 44787 1607 44799 1783
rect 44741 1595 44799 1607
rect 44855 1783 44913 1795
rect 44855 1607 44867 1783
rect 44901 1607 44913 1783
rect 44855 1595 44913 1607
rect 45113 1783 45171 1795
rect 45113 1607 45125 1783
rect 45159 1607 45171 1783
rect 45113 1595 45171 1607
rect 45227 1783 45285 1795
rect 45227 1607 45239 1783
rect 45273 1607 45285 1783
rect 45227 1595 45285 1607
rect 45485 1783 45543 1795
rect 45485 1607 45497 1783
rect 45531 1607 45543 1783
rect 45485 1595 45543 1607
rect 45599 1783 45657 1795
rect 45599 1607 45611 1783
rect 45645 1607 45657 1783
rect 45599 1595 45657 1607
rect 45857 1783 45915 1795
rect 45857 1607 45869 1783
rect 45903 1607 45915 1783
rect 45857 1595 45915 1607
rect 45971 1783 46029 1795
rect 45971 1607 45983 1783
rect 46017 1607 46029 1783
rect 45971 1595 46029 1607
rect 46229 1783 46287 1795
rect 46229 1607 46241 1783
rect 46275 1607 46287 1783
rect 46229 1595 46287 1607
rect 46343 1783 46401 1795
rect 46343 1607 46355 1783
rect 46389 1607 46401 1783
rect 46343 1595 46401 1607
rect 46601 1783 46659 1795
rect 46601 1607 46613 1783
rect 46647 1607 46659 1783
rect 46601 1595 46659 1607
rect 46715 1783 46773 1795
rect 46715 1607 46727 1783
rect 46761 1607 46773 1783
rect 46715 1595 46773 1607
rect 46973 1783 47031 1795
rect 46973 1607 46985 1783
rect 47019 1607 47031 1783
rect 46973 1595 47031 1607
rect 47087 1783 47145 1795
rect 47087 1607 47099 1783
rect 47133 1607 47145 1783
rect 47087 1595 47145 1607
rect 47345 1783 47403 1795
rect 47345 1607 47357 1783
rect 47391 1607 47403 1783
rect 47345 1595 47403 1607
rect 47459 1783 47517 1795
rect 47459 1607 47471 1783
rect 47505 1607 47517 1783
rect 47459 1595 47517 1607
rect 47717 1783 47775 1795
rect 47717 1607 47729 1783
rect 47763 1607 47775 1783
rect 47717 1595 47775 1607
rect 47831 1783 47889 1795
rect 47831 1607 47843 1783
rect 47877 1607 47889 1783
rect 47831 1595 47889 1607
rect 48089 1783 48147 1795
rect 48089 1607 48101 1783
rect 48135 1607 48147 1783
rect 48089 1595 48147 1607
rect 48203 1783 48261 1795
rect 48203 1607 48215 1783
rect 48249 1607 48261 1783
rect 48203 1595 48261 1607
rect 48461 1783 48519 1795
rect 48461 1607 48473 1783
rect 48507 1607 48519 1783
rect 48461 1595 48519 1607
rect 48575 1783 48633 1795
rect 48575 1607 48587 1783
rect 48621 1607 48633 1783
rect 48575 1595 48633 1607
rect 48833 1783 48891 1795
rect 48833 1607 48845 1783
rect 48879 1607 48891 1783
rect 48833 1595 48891 1607
rect 48947 1783 49005 1795
rect 48947 1607 48959 1783
rect 48993 1607 49005 1783
rect 48947 1595 49005 1607
rect 49205 1783 49263 1795
rect 49205 1607 49217 1783
rect 49251 1607 49263 1783
rect 49205 1595 49263 1607
rect 49319 1783 49377 1795
rect 49319 1607 49331 1783
rect 49365 1607 49377 1783
rect 49319 1595 49377 1607
rect 49577 1783 49635 1795
rect 49577 1607 49589 1783
rect 49623 1607 49635 1783
rect 49577 1595 49635 1607
rect 40763 1365 40821 1377
rect 40763 1189 40775 1365
rect 40809 1189 40821 1365
rect 40763 1177 40821 1189
rect 41021 1365 41079 1377
rect 41021 1189 41033 1365
rect 41067 1189 41079 1365
rect 41021 1177 41079 1189
rect 41135 1365 41193 1377
rect 41135 1189 41147 1365
rect 41181 1189 41193 1365
rect 41135 1177 41193 1189
rect 41393 1365 41451 1377
rect 41393 1189 41405 1365
rect 41439 1189 41451 1365
rect 41393 1177 41451 1189
rect 41507 1365 41565 1377
rect 41507 1189 41519 1365
rect 41553 1189 41565 1365
rect 41507 1177 41565 1189
rect 41765 1365 41823 1377
rect 41765 1189 41777 1365
rect 41811 1189 41823 1365
rect 41765 1177 41823 1189
rect 41879 1365 41937 1377
rect 41879 1189 41891 1365
rect 41925 1189 41937 1365
rect 41879 1177 41937 1189
rect 42137 1365 42195 1377
rect 42137 1189 42149 1365
rect 42183 1189 42195 1365
rect 42137 1177 42195 1189
rect 42251 1365 42309 1377
rect 42251 1189 42263 1365
rect 42297 1189 42309 1365
rect 42251 1177 42309 1189
rect 42509 1365 42567 1377
rect 42509 1189 42521 1365
rect 42555 1189 42567 1365
rect 42509 1177 42567 1189
rect 42623 1365 42681 1377
rect 42623 1189 42635 1365
rect 42669 1189 42681 1365
rect 42623 1177 42681 1189
rect 42881 1365 42939 1377
rect 42881 1189 42893 1365
rect 42927 1189 42939 1365
rect 42881 1177 42939 1189
rect 42995 1365 43053 1377
rect 42995 1189 43007 1365
rect 43041 1189 43053 1365
rect 42995 1177 43053 1189
rect 43253 1365 43311 1377
rect 43253 1189 43265 1365
rect 43299 1189 43311 1365
rect 43253 1177 43311 1189
rect 43367 1365 43425 1377
rect 43367 1189 43379 1365
rect 43413 1189 43425 1365
rect 43367 1177 43425 1189
rect 43625 1365 43683 1377
rect 43625 1189 43637 1365
rect 43671 1189 43683 1365
rect 43625 1177 43683 1189
rect 43739 1365 43797 1377
rect 43739 1189 43751 1365
rect 43785 1189 43797 1365
rect 43739 1177 43797 1189
rect 43997 1365 44055 1377
rect 43997 1189 44009 1365
rect 44043 1189 44055 1365
rect 43997 1177 44055 1189
rect 44111 1365 44169 1377
rect 44111 1189 44123 1365
rect 44157 1189 44169 1365
rect 44111 1177 44169 1189
rect 44369 1365 44427 1377
rect 44369 1189 44381 1365
rect 44415 1189 44427 1365
rect 44369 1177 44427 1189
rect 44483 1365 44541 1377
rect 44483 1189 44495 1365
rect 44529 1189 44541 1365
rect 44483 1177 44541 1189
rect 44741 1365 44799 1377
rect 44741 1189 44753 1365
rect 44787 1189 44799 1365
rect 44741 1177 44799 1189
rect 44855 1365 44913 1377
rect 44855 1189 44867 1365
rect 44901 1189 44913 1365
rect 44855 1177 44913 1189
rect 45113 1365 45171 1377
rect 45113 1189 45125 1365
rect 45159 1189 45171 1365
rect 45113 1177 45171 1189
rect 45227 1365 45285 1377
rect 45227 1189 45239 1365
rect 45273 1189 45285 1365
rect 45227 1177 45285 1189
rect 45485 1365 45543 1377
rect 45485 1189 45497 1365
rect 45531 1189 45543 1365
rect 45485 1177 45543 1189
rect 45599 1365 45657 1377
rect 45599 1189 45611 1365
rect 45645 1189 45657 1365
rect 45599 1177 45657 1189
rect 45857 1365 45915 1377
rect 45857 1189 45869 1365
rect 45903 1189 45915 1365
rect 45857 1177 45915 1189
rect 45971 1365 46029 1377
rect 45971 1189 45983 1365
rect 46017 1189 46029 1365
rect 45971 1177 46029 1189
rect 46229 1365 46287 1377
rect 46229 1189 46241 1365
rect 46275 1189 46287 1365
rect 46229 1177 46287 1189
rect 46343 1365 46401 1377
rect 46343 1189 46355 1365
rect 46389 1189 46401 1365
rect 46343 1177 46401 1189
rect 46601 1365 46659 1377
rect 46601 1189 46613 1365
rect 46647 1189 46659 1365
rect 46601 1177 46659 1189
rect 46715 1365 46773 1377
rect 46715 1189 46727 1365
rect 46761 1189 46773 1365
rect 46715 1177 46773 1189
rect 46973 1365 47031 1377
rect 46973 1189 46985 1365
rect 47019 1189 47031 1365
rect 46973 1177 47031 1189
rect 47087 1365 47145 1377
rect 47087 1189 47099 1365
rect 47133 1189 47145 1365
rect 47087 1177 47145 1189
rect 47345 1365 47403 1377
rect 47345 1189 47357 1365
rect 47391 1189 47403 1365
rect 47345 1177 47403 1189
rect 47459 1365 47517 1377
rect 47459 1189 47471 1365
rect 47505 1189 47517 1365
rect 47459 1177 47517 1189
rect 47717 1365 47775 1377
rect 47717 1189 47729 1365
rect 47763 1189 47775 1365
rect 47717 1177 47775 1189
rect 47831 1365 47889 1377
rect 47831 1189 47843 1365
rect 47877 1189 47889 1365
rect 47831 1177 47889 1189
rect 48089 1365 48147 1377
rect 48089 1189 48101 1365
rect 48135 1189 48147 1365
rect 48089 1177 48147 1189
rect 48203 1365 48261 1377
rect 48203 1189 48215 1365
rect 48249 1189 48261 1365
rect 48203 1177 48261 1189
rect 48461 1365 48519 1377
rect 48461 1189 48473 1365
rect 48507 1189 48519 1365
rect 48461 1177 48519 1189
rect 48575 1365 48633 1377
rect 48575 1189 48587 1365
rect 48621 1189 48633 1365
rect 48575 1177 48633 1189
rect 48833 1365 48891 1377
rect 48833 1189 48845 1365
rect 48879 1189 48891 1365
rect 48833 1177 48891 1189
rect 48947 1365 49005 1377
rect 48947 1189 48959 1365
rect 48993 1189 49005 1365
rect 48947 1177 49005 1189
rect 49205 1365 49263 1377
rect 49205 1189 49217 1365
rect 49251 1189 49263 1365
rect 49205 1177 49263 1189
rect 49319 1365 49377 1377
rect 49319 1189 49331 1365
rect 49365 1189 49377 1365
rect 49319 1177 49377 1189
rect 49577 1365 49635 1377
rect 49577 1189 49589 1365
rect 49623 1189 49635 1365
rect 49577 1177 49635 1189
rect 40763 947 40821 959
rect 40763 771 40775 947
rect 40809 771 40821 947
rect 40763 759 40821 771
rect 41021 947 41079 959
rect 41021 771 41033 947
rect 41067 771 41079 947
rect 41021 759 41079 771
rect 41135 947 41193 959
rect 41135 771 41147 947
rect 41181 771 41193 947
rect 41135 759 41193 771
rect 41393 947 41451 959
rect 41393 771 41405 947
rect 41439 771 41451 947
rect 41393 759 41451 771
rect 41507 947 41565 959
rect 41507 771 41519 947
rect 41553 771 41565 947
rect 41507 759 41565 771
rect 41765 947 41823 959
rect 41765 771 41777 947
rect 41811 771 41823 947
rect 41765 759 41823 771
rect 41879 947 41937 959
rect 41879 771 41891 947
rect 41925 771 41937 947
rect 41879 759 41937 771
rect 42137 947 42195 959
rect 42137 771 42149 947
rect 42183 771 42195 947
rect 42137 759 42195 771
rect 42251 947 42309 959
rect 42251 771 42263 947
rect 42297 771 42309 947
rect 42251 759 42309 771
rect 42509 947 42567 959
rect 42509 771 42521 947
rect 42555 771 42567 947
rect 42509 759 42567 771
rect 42623 947 42681 959
rect 42623 771 42635 947
rect 42669 771 42681 947
rect 42623 759 42681 771
rect 42881 947 42939 959
rect 42881 771 42893 947
rect 42927 771 42939 947
rect 42881 759 42939 771
rect 42995 947 43053 959
rect 42995 771 43007 947
rect 43041 771 43053 947
rect 42995 759 43053 771
rect 43253 947 43311 959
rect 43253 771 43265 947
rect 43299 771 43311 947
rect 43253 759 43311 771
rect 43367 947 43425 959
rect 43367 771 43379 947
rect 43413 771 43425 947
rect 43367 759 43425 771
rect 43625 947 43683 959
rect 43625 771 43637 947
rect 43671 771 43683 947
rect 43625 759 43683 771
rect 43739 947 43797 959
rect 43739 771 43751 947
rect 43785 771 43797 947
rect 43739 759 43797 771
rect 43997 947 44055 959
rect 43997 771 44009 947
rect 44043 771 44055 947
rect 43997 759 44055 771
rect 44111 947 44169 959
rect 44111 771 44123 947
rect 44157 771 44169 947
rect 44111 759 44169 771
rect 44369 947 44427 959
rect 44369 771 44381 947
rect 44415 771 44427 947
rect 44369 759 44427 771
rect 44483 947 44541 959
rect 44483 771 44495 947
rect 44529 771 44541 947
rect 44483 759 44541 771
rect 44741 947 44799 959
rect 44741 771 44753 947
rect 44787 771 44799 947
rect 44741 759 44799 771
rect 44855 947 44913 959
rect 44855 771 44867 947
rect 44901 771 44913 947
rect 44855 759 44913 771
rect 45113 947 45171 959
rect 45113 771 45125 947
rect 45159 771 45171 947
rect 45113 759 45171 771
rect 45227 947 45285 959
rect 45227 771 45239 947
rect 45273 771 45285 947
rect 45227 759 45285 771
rect 45485 947 45543 959
rect 45485 771 45497 947
rect 45531 771 45543 947
rect 45485 759 45543 771
rect 45599 947 45657 959
rect 45599 771 45611 947
rect 45645 771 45657 947
rect 45599 759 45657 771
rect 45857 947 45915 959
rect 45857 771 45869 947
rect 45903 771 45915 947
rect 45857 759 45915 771
rect 45971 947 46029 959
rect 45971 771 45983 947
rect 46017 771 46029 947
rect 45971 759 46029 771
rect 46229 947 46287 959
rect 46229 771 46241 947
rect 46275 771 46287 947
rect 46229 759 46287 771
rect 46343 947 46401 959
rect 46343 771 46355 947
rect 46389 771 46401 947
rect 46343 759 46401 771
rect 46601 947 46659 959
rect 46601 771 46613 947
rect 46647 771 46659 947
rect 46601 759 46659 771
rect 46715 947 46773 959
rect 46715 771 46727 947
rect 46761 771 46773 947
rect 46715 759 46773 771
rect 46973 947 47031 959
rect 46973 771 46985 947
rect 47019 771 47031 947
rect 46973 759 47031 771
rect 47087 947 47145 959
rect 47087 771 47099 947
rect 47133 771 47145 947
rect 47087 759 47145 771
rect 47345 947 47403 959
rect 47345 771 47357 947
rect 47391 771 47403 947
rect 47345 759 47403 771
rect 47459 947 47517 959
rect 47459 771 47471 947
rect 47505 771 47517 947
rect 47459 759 47517 771
rect 47717 947 47775 959
rect 47717 771 47729 947
rect 47763 771 47775 947
rect 47717 759 47775 771
rect 47831 947 47889 959
rect 47831 771 47843 947
rect 47877 771 47889 947
rect 47831 759 47889 771
rect 48089 947 48147 959
rect 48089 771 48101 947
rect 48135 771 48147 947
rect 48089 759 48147 771
rect 48203 947 48261 959
rect 48203 771 48215 947
rect 48249 771 48261 947
rect 48203 759 48261 771
rect 48461 947 48519 959
rect 48461 771 48473 947
rect 48507 771 48519 947
rect 48461 759 48519 771
rect 48575 947 48633 959
rect 48575 771 48587 947
rect 48621 771 48633 947
rect 48575 759 48633 771
rect 48833 947 48891 959
rect 48833 771 48845 947
rect 48879 771 48891 947
rect 48833 759 48891 771
rect 48947 947 49005 959
rect 48947 771 48959 947
rect 48993 771 49005 947
rect 48947 759 49005 771
rect 49205 947 49263 959
rect 49205 771 49217 947
rect 49251 771 49263 947
rect 49205 759 49263 771
rect 49319 947 49377 959
rect 49319 771 49331 947
rect 49365 771 49377 947
rect 49319 759 49377 771
rect 49577 947 49635 959
rect 49577 771 49589 947
rect 49623 771 49635 947
rect 49577 759 49635 771
rect 40763 529 40821 541
rect 40763 353 40775 529
rect 40809 353 40821 529
rect 40763 341 40821 353
rect 41021 529 41079 541
rect 41021 353 41033 529
rect 41067 353 41079 529
rect 41021 341 41079 353
rect 41135 529 41193 541
rect 41135 353 41147 529
rect 41181 353 41193 529
rect 41135 341 41193 353
rect 41393 529 41451 541
rect 41393 353 41405 529
rect 41439 353 41451 529
rect 41393 341 41451 353
rect 41507 529 41565 541
rect 41507 353 41519 529
rect 41553 353 41565 529
rect 41507 341 41565 353
rect 41765 529 41823 541
rect 41765 353 41777 529
rect 41811 353 41823 529
rect 41765 341 41823 353
rect 41879 529 41937 541
rect 41879 353 41891 529
rect 41925 353 41937 529
rect 41879 341 41937 353
rect 42137 529 42195 541
rect 42137 353 42149 529
rect 42183 353 42195 529
rect 42137 341 42195 353
rect 42251 529 42309 541
rect 42251 353 42263 529
rect 42297 353 42309 529
rect 42251 341 42309 353
rect 42509 529 42567 541
rect 42509 353 42521 529
rect 42555 353 42567 529
rect 42509 341 42567 353
rect 42623 529 42681 541
rect 42623 353 42635 529
rect 42669 353 42681 529
rect 42623 341 42681 353
rect 42881 529 42939 541
rect 42881 353 42893 529
rect 42927 353 42939 529
rect 42881 341 42939 353
rect 42995 529 43053 541
rect 42995 353 43007 529
rect 43041 353 43053 529
rect 42995 341 43053 353
rect 43253 529 43311 541
rect 43253 353 43265 529
rect 43299 353 43311 529
rect 43253 341 43311 353
rect 43367 529 43425 541
rect 43367 353 43379 529
rect 43413 353 43425 529
rect 43367 341 43425 353
rect 43625 529 43683 541
rect 43625 353 43637 529
rect 43671 353 43683 529
rect 43625 341 43683 353
rect 43739 529 43797 541
rect 43739 353 43751 529
rect 43785 353 43797 529
rect 43739 341 43797 353
rect 43997 529 44055 541
rect 43997 353 44009 529
rect 44043 353 44055 529
rect 43997 341 44055 353
rect 44111 529 44169 541
rect 44111 353 44123 529
rect 44157 353 44169 529
rect 44111 341 44169 353
rect 44369 529 44427 541
rect 44369 353 44381 529
rect 44415 353 44427 529
rect 44369 341 44427 353
rect 44483 529 44541 541
rect 44483 353 44495 529
rect 44529 353 44541 529
rect 44483 341 44541 353
rect 44741 529 44799 541
rect 44741 353 44753 529
rect 44787 353 44799 529
rect 44741 341 44799 353
rect 44855 529 44913 541
rect 44855 353 44867 529
rect 44901 353 44913 529
rect 44855 341 44913 353
rect 45113 529 45171 541
rect 45113 353 45125 529
rect 45159 353 45171 529
rect 45113 341 45171 353
rect 45227 529 45285 541
rect 45227 353 45239 529
rect 45273 353 45285 529
rect 45227 341 45285 353
rect 45485 529 45543 541
rect 45485 353 45497 529
rect 45531 353 45543 529
rect 45485 341 45543 353
rect 45599 529 45657 541
rect 45599 353 45611 529
rect 45645 353 45657 529
rect 45599 341 45657 353
rect 45857 529 45915 541
rect 45857 353 45869 529
rect 45903 353 45915 529
rect 45857 341 45915 353
rect 45971 529 46029 541
rect 45971 353 45983 529
rect 46017 353 46029 529
rect 45971 341 46029 353
rect 46229 529 46287 541
rect 46229 353 46241 529
rect 46275 353 46287 529
rect 46229 341 46287 353
rect 46343 529 46401 541
rect 46343 353 46355 529
rect 46389 353 46401 529
rect 46343 341 46401 353
rect 46601 529 46659 541
rect 46601 353 46613 529
rect 46647 353 46659 529
rect 46601 341 46659 353
rect 46715 529 46773 541
rect 46715 353 46727 529
rect 46761 353 46773 529
rect 46715 341 46773 353
rect 46973 529 47031 541
rect 46973 353 46985 529
rect 47019 353 47031 529
rect 46973 341 47031 353
rect 47087 529 47145 541
rect 47087 353 47099 529
rect 47133 353 47145 529
rect 47087 341 47145 353
rect 47345 529 47403 541
rect 47345 353 47357 529
rect 47391 353 47403 529
rect 47345 341 47403 353
rect 47459 529 47517 541
rect 47459 353 47471 529
rect 47505 353 47517 529
rect 47459 341 47517 353
rect 47717 529 47775 541
rect 47717 353 47729 529
rect 47763 353 47775 529
rect 47717 341 47775 353
rect 47831 529 47889 541
rect 47831 353 47843 529
rect 47877 353 47889 529
rect 47831 341 47889 353
rect 48089 529 48147 541
rect 48089 353 48101 529
rect 48135 353 48147 529
rect 48089 341 48147 353
rect 48203 529 48261 541
rect 48203 353 48215 529
rect 48249 353 48261 529
rect 48203 341 48261 353
rect 48461 529 48519 541
rect 48461 353 48473 529
rect 48507 353 48519 529
rect 48461 341 48519 353
rect 48575 529 48633 541
rect 48575 353 48587 529
rect 48621 353 48633 529
rect 48575 341 48633 353
rect 48833 529 48891 541
rect 48833 353 48845 529
rect 48879 353 48891 529
rect 48833 341 48891 353
rect 48947 529 49005 541
rect 48947 353 48959 529
rect 48993 353 49005 529
rect 48947 341 49005 353
rect 49205 529 49263 541
rect 49205 353 49217 529
rect 49251 353 49263 529
rect 49205 341 49263 353
rect 49319 529 49377 541
rect 49319 353 49331 529
rect 49365 353 49377 529
rect 49319 341 49377 353
rect 49577 529 49635 541
rect 49577 353 49589 529
rect 49623 353 49635 529
rect 49577 341 49635 353
<< pdiff >>
rect 40763 17281 40821 17293
rect 40763 16505 40775 17281
rect 40809 16505 40821 17281
rect 40763 16493 40821 16505
rect 41021 17281 41079 17293
rect 41021 16505 41033 17281
rect 41067 16505 41079 17281
rect 41021 16493 41079 16505
rect 41135 17281 41193 17293
rect 41135 16505 41147 17281
rect 41181 16505 41193 17281
rect 41135 16493 41193 16505
rect 41393 17281 41451 17293
rect 41393 16505 41405 17281
rect 41439 16505 41451 17281
rect 41393 16493 41451 16505
rect 41507 17281 41565 17293
rect 41507 16505 41519 17281
rect 41553 16505 41565 17281
rect 41507 16493 41565 16505
rect 41765 17281 41823 17293
rect 41765 16505 41777 17281
rect 41811 16505 41823 17281
rect 41765 16493 41823 16505
rect 41879 17281 41937 17293
rect 41879 16505 41891 17281
rect 41925 16505 41937 17281
rect 41879 16493 41937 16505
rect 42137 17281 42195 17293
rect 42137 16505 42149 17281
rect 42183 16505 42195 17281
rect 42137 16493 42195 16505
rect 42251 17281 42309 17293
rect 42251 16505 42263 17281
rect 42297 16505 42309 17281
rect 42251 16493 42309 16505
rect 42509 17281 42567 17293
rect 42509 16505 42521 17281
rect 42555 16505 42567 17281
rect 42509 16493 42567 16505
rect 42623 17281 42681 17293
rect 42623 16505 42635 17281
rect 42669 16505 42681 17281
rect 42623 16493 42681 16505
rect 42881 17281 42939 17293
rect 42881 16505 42893 17281
rect 42927 16505 42939 17281
rect 42881 16493 42939 16505
rect 42995 17281 43053 17293
rect 42995 16505 43007 17281
rect 43041 16505 43053 17281
rect 42995 16493 43053 16505
rect 43253 17281 43311 17293
rect 43253 16505 43265 17281
rect 43299 16505 43311 17281
rect 43253 16493 43311 16505
rect 43367 17281 43425 17293
rect 43367 16505 43379 17281
rect 43413 16505 43425 17281
rect 43367 16493 43425 16505
rect 43625 17281 43683 17293
rect 43625 16505 43637 17281
rect 43671 16505 43683 17281
rect 43625 16493 43683 16505
rect 40763 16245 40821 16257
rect 40763 15469 40775 16245
rect 40809 15469 40821 16245
rect 40763 15457 40821 15469
rect 41021 16245 41079 16257
rect 41021 15469 41033 16245
rect 41067 15469 41079 16245
rect 41021 15457 41079 15469
rect 41135 16245 41193 16257
rect 41135 15469 41147 16245
rect 41181 15469 41193 16245
rect 41135 15457 41193 15469
rect 41393 16245 41451 16257
rect 41393 15469 41405 16245
rect 41439 15469 41451 16245
rect 41393 15457 41451 15469
rect 41507 16245 41565 16257
rect 41507 15469 41519 16245
rect 41553 15469 41565 16245
rect 41507 15457 41565 15469
rect 41765 16245 41823 16257
rect 41765 15469 41777 16245
rect 41811 15469 41823 16245
rect 41765 15457 41823 15469
rect 41879 16245 41937 16257
rect 41879 15469 41891 16245
rect 41925 15469 41937 16245
rect 41879 15457 41937 15469
rect 42137 16245 42195 16257
rect 42137 15469 42149 16245
rect 42183 15469 42195 16245
rect 42137 15457 42195 15469
rect 42251 16245 42309 16257
rect 42251 15469 42263 16245
rect 42297 15469 42309 16245
rect 42251 15457 42309 15469
rect 42509 16245 42567 16257
rect 42509 15469 42521 16245
rect 42555 15469 42567 16245
rect 42509 15457 42567 15469
rect 42623 16245 42681 16257
rect 42623 15469 42635 16245
rect 42669 15469 42681 16245
rect 42623 15457 42681 15469
rect 42881 16245 42939 16257
rect 42881 15469 42893 16245
rect 42927 15469 42939 16245
rect 42881 15457 42939 15469
rect 42995 16245 43053 16257
rect 42995 15469 43007 16245
rect 43041 15469 43053 16245
rect 42995 15457 43053 15469
rect 43253 16245 43311 16257
rect 43253 15469 43265 16245
rect 43299 15469 43311 16245
rect 43253 15457 43311 15469
rect 43367 16245 43425 16257
rect 43367 15469 43379 16245
rect 43413 15469 43425 16245
rect 43367 15457 43425 15469
rect 43625 16245 43683 16257
rect 43625 15469 43637 16245
rect 43671 15469 43683 16245
rect 43625 15457 43683 15469
rect 40763 15209 40821 15221
rect 40763 14433 40775 15209
rect 40809 14433 40821 15209
rect 40763 14421 40821 14433
rect 41021 15209 41079 15221
rect 41021 14433 41033 15209
rect 41067 14433 41079 15209
rect 41021 14421 41079 14433
rect 41135 15209 41193 15221
rect 41135 14433 41147 15209
rect 41181 14433 41193 15209
rect 41135 14421 41193 14433
rect 41393 15209 41451 15221
rect 41393 14433 41405 15209
rect 41439 14433 41451 15209
rect 41393 14421 41451 14433
rect 41507 15209 41565 15221
rect 41507 14433 41519 15209
rect 41553 14433 41565 15209
rect 41507 14421 41565 14433
rect 41765 15209 41823 15221
rect 41765 14433 41777 15209
rect 41811 14433 41823 15209
rect 41765 14421 41823 14433
rect 41879 15209 41937 15221
rect 41879 14433 41891 15209
rect 41925 14433 41937 15209
rect 41879 14421 41937 14433
rect 42137 15209 42195 15221
rect 42137 14433 42149 15209
rect 42183 14433 42195 15209
rect 42137 14421 42195 14433
rect 42251 15209 42309 15221
rect 42251 14433 42263 15209
rect 42297 14433 42309 15209
rect 42251 14421 42309 14433
rect 42509 15209 42567 15221
rect 42509 14433 42521 15209
rect 42555 14433 42567 15209
rect 42509 14421 42567 14433
rect 42623 15209 42681 15221
rect 42623 14433 42635 15209
rect 42669 14433 42681 15209
rect 42623 14421 42681 14433
rect 42881 15209 42939 15221
rect 42881 14433 42893 15209
rect 42927 14433 42939 15209
rect 42881 14421 42939 14433
rect 42995 15209 43053 15221
rect 42995 14433 43007 15209
rect 43041 14433 43053 15209
rect 42995 14421 43053 14433
rect 43253 15209 43311 15221
rect 43253 14433 43265 15209
rect 43299 14433 43311 15209
rect 43253 14421 43311 14433
rect 43367 15209 43425 15221
rect 43367 14433 43379 15209
rect 43413 14433 43425 15209
rect 43367 14421 43425 14433
rect 43625 15209 43683 15221
rect 43625 14433 43637 15209
rect 43671 14433 43683 15209
rect 43625 14421 43683 14433
rect 40763 14173 40821 14185
rect 40763 13397 40775 14173
rect 40809 13397 40821 14173
rect 40763 13385 40821 13397
rect 41021 14173 41079 14185
rect 41021 13397 41033 14173
rect 41067 13397 41079 14173
rect 41021 13385 41079 13397
rect 41135 14173 41193 14185
rect 41135 13397 41147 14173
rect 41181 13397 41193 14173
rect 41135 13385 41193 13397
rect 41393 14173 41451 14185
rect 41393 13397 41405 14173
rect 41439 13397 41451 14173
rect 41393 13385 41451 13397
rect 41507 14173 41565 14185
rect 41507 13397 41519 14173
rect 41553 13397 41565 14173
rect 41507 13385 41565 13397
rect 41765 14173 41823 14185
rect 41765 13397 41777 14173
rect 41811 13397 41823 14173
rect 41765 13385 41823 13397
rect 41879 14173 41937 14185
rect 41879 13397 41891 14173
rect 41925 13397 41937 14173
rect 41879 13385 41937 13397
rect 42137 14173 42195 14185
rect 42137 13397 42149 14173
rect 42183 13397 42195 14173
rect 42137 13385 42195 13397
rect 42251 14173 42309 14185
rect 42251 13397 42263 14173
rect 42297 13397 42309 14173
rect 42251 13385 42309 13397
rect 42509 14173 42567 14185
rect 42509 13397 42521 14173
rect 42555 13397 42567 14173
rect 42509 13385 42567 13397
rect 42623 14173 42681 14185
rect 42623 13397 42635 14173
rect 42669 13397 42681 14173
rect 42623 13385 42681 13397
rect 42881 14173 42939 14185
rect 42881 13397 42893 14173
rect 42927 13397 42939 14173
rect 42881 13385 42939 13397
rect 42995 14173 43053 14185
rect 42995 13397 43007 14173
rect 43041 13397 43053 14173
rect 42995 13385 43053 13397
rect 43253 14173 43311 14185
rect 43253 13397 43265 14173
rect 43299 13397 43311 14173
rect 43253 13385 43311 13397
rect 43367 14173 43425 14185
rect 43367 13397 43379 14173
rect 43413 13397 43425 14173
rect 43367 13385 43425 13397
rect 43625 14173 43683 14185
rect 43625 13397 43637 14173
rect 43671 13397 43683 14173
rect 43625 13385 43683 13397
rect 39275 12657 39333 12669
rect 39275 12281 39287 12657
rect 39321 12281 39333 12657
rect 39275 12269 39333 12281
rect 39533 12657 39591 12669
rect 39533 12281 39545 12657
rect 39579 12281 39591 12657
rect 39533 12269 39591 12281
rect 39647 12657 39705 12669
rect 39647 12281 39659 12657
rect 39693 12281 39705 12657
rect 39647 12269 39705 12281
rect 39905 12657 39963 12669
rect 39905 12281 39917 12657
rect 39951 12281 39963 12657
rect 39905 12269 39963 12281
rect 40019 12657 40077 12669
rect 40019 12281 40031 12657
rect 40065 12281 40077 12657
rect 40019 12269 40077 12281
rect 40277 12657 40335 12669
rect 40277 12281 40289 12657
rect 40323 12281 40335 12657
rect 40277 12269 40335 12281
rect 40391 12657 40449 12669
rect 40391 12281 40403 12657
rect 40437 12281 40449 12657
rect 40391 12269 40449 12281
rect 40649 12657 40707 12669
rect 40649 12281 40661 12657
rect 40695 12281 40707 12657
rect 40649 12269 40707 12281
rect 40763 12657 40821 12669
rect 40763 12281 40775 12657
rect 40809 12281 40821 12657
rect 40763 12269 40821 12281
rect 41021 12657 41079 12669
rect 41021 12281 41033 12657
rect 41067 12281 41079 12657
rect 41021 12269 41079 12281
rect 41135 12657 41193 12669
rect 41135 12281 41147 12657
rect 41181 12281 41193 12657
rect 41135 12269 41193 12281
rect 41393 12657 41451 12669
rect 41393 12281 41405 12657
rect 41439 12281 41451 12657
rect 41393 12269 41451 12281
rect 41507 12657 41565 12669
rect 41507 12281 41519 12657
rect 41553 12281 41565 12657
rect 41507 12269 41565 12281
rect 41765 12657 41823 12669
rect 41765 12281 41777 12657
rect 41811 12281 41823 12657
rect 41765 12269 41823 12281
rect 41879 12657 41937 12669
rect 41879 12281 41891 12657
rect 41925 12281 41937 12657
rect 41879 12269 41937 12281
rect 42137 12657 42195 12669
rect 42137 12281 42149 12657
rect 42183 12281 42195 12657
rect 42137 12269 42195 12281
rect 42251 12657 42309 12669
rect 42251 12281 42263 12657
rect 42297 12281 42309 12657
rect 42251 12269 42309 12281
rect 42509 12657 42567 12669
rect 42509 12281 42521 12657
rect 42555 12281 42567 12657
rect 42509 12269 42567 12281
rect 42623 12657 42681 12669
rect 42623 12281 42635 12657
rect 42669 12281 42681 12657
rect 42623 12269 42681 12281
rect 42881 12657 42939 12669
rect 42881 12281 42893 12657
rect 42927 12281 42939 12657
rect 42881 12269 42939 12281
rect 42995 12657 43053 12669
rect 42995 12281 43007 12657
rect 43041 12281 43053 12657
rect 42995 12269 43053 12281
rect 43253 12657 43311 12669
rect 43253 12281 43265 12657
rect 43299 12281 43311 12657
rect 43253 12269 43311 12281
rect 43367 12657 43425 12669
rect 43367 12281 43379 12657
rect 43413 12281 43425 12657
rect 43367 12269 43425 12281
rect 43625 12657 43683 12669
rect 43625 12281 43637 12657
rect 43671 12281 43683 12657
rect 43625 12269 43683 12281
rect 43739 12657 43797 12669
rect 43739 12281 43751 12657
rect 43785 12281 43797 12657
rect 43739 12269 43797 12281
rect 43997 12657 44055 12669
rect 43997 12281 44009 12657
rect 44043 12281 44055 12657
rect 43997 12269 44055 12281
rect 44111 12657 44169 12669
rect 44111 12281 44123 12657
rect 44157 12281 44169 12657
rect 44111 12269 44169 12281
rect 44369 12657 44427 12669
rect 44369 12281 44381 12657
rect 44415 12281 44427 12657
rect 44369 12269 44427 12281
rect 44483 12657 44541 12669
rect 44483 12281 44495 12657
rect 44529 12281 44541 12657
rect 44483 12269 44541 12281
rect 44741 12657 44799 12669
rect 44741 12281 44753 12657
rect 44787 12281 44799 12657
rect 44741 12269 44799 12281
rect 44855 12657 44913 12669
rect 44855 12281 44867 12657
rect 44901 12281 44913 12657
rect 44855 12269 44913 12281
rect 45113 12657 45171 12669
rect 45113 12281 45125 12657
rect 45159 12281 45171 12657
rect 45113 12269 45171 12281
rect 45227 12657 45285 12669
rect 45227 12281 45239 12657
rect 45273 12281 45285 12657
rect 45227 12269 45285 12281
rect 45485 12657 45543 12669
rect 45485 12281 45497 12657
rect 45531 12281 45543 12657
rect 45485 12269 45543 12281
rect 45599 12657 45657 12669
rect 45599 12281 45611 12657
rect 45645 12281 45657 12657
rect 45599 12269 45657 12281
rect 45857 12657 45915 12669
rect 45857 12281 45869 12657
rect 45903 12281 45915 12657
rect 45857 12269 45915 12281
rect 45971 12657 46029 12669
rect 45971 12281 45983 12657
rect 46017 12281 46029 12657
rect 45971 12269 46029 12281
rect 46229 12657 46287 12669
rect 46229 12281 46241 12657
rect 46275 12281 46287 12657
rect 46229 12269 46287 12281
rect 46343 12657 46401 12669
rect 46343 12281 46355 12657
rect 46389 12281 46401 12657
rect 46343 12269 46401 12281
rect 46601 12657 46659 12669
rect 46601 12281 46613 12657
rect 46647 12281 46659 12657
rect 46601 12269 46659 12281
rect 46715 12657 46773 12669
rect 46715 12281 46727 12657
rect 46761 12281 46773 12657
rect 46715 12269 46773 12281
rect 46973 12657 47031 12669
rect 46973 12281 46985 12657
rect 47019 12281 47031 12657
rect 46973 12269 47031 12281
rect 47087 12657 47145 12669
rect 47087 12281 47099 12657
rect 47133 12281 47145 12657
rect 47087 12269 47145 12281
rect 47345 12657 47403 12669
rect 47345 12281 47357 12657
rect 47391 12281 47403 12657
rect 47345 12269 47403 12281
rect 47459 12657 47517 12669
rect 47459 12281 47471 12657
rect 47505 12281 47517 12657
rect 47459 12269 47517 12281
rect 47717 12657 47775 12669
rect 47717 12281 47729 12657
rect 47763 12281 47775 12657
rect 47717 12269 47775 12281
rect 47831 12657 47889 12669
rect 47831 12281 47843 12657
rect 47877 12281 47889 12657
rect 47831 12269 47889 12281
rect 48089 12657 48147 12669
rect 48089 12281 48101 12657
rect 48135 12281 48147 12657
rect 48089 12269 48147 12281
rect 48203 12657 48261 12669
rect 48203 12281 48215 12657
rect 48249 12281 48261 12657
rect 48203 12269 48261 12281
rect 48461 12657 48519 12669
rect 48461 12281 48473 12657
rect 48507 12281 48519 12657
rect 48461 12269 48519 12281
rect 48575 12657 48633 12669
rect 48575 12281 48587 12657
rect 48621 12281 48633 12657
rect 48575 12269 48633 12281
rect 48833 12657 48891 12669
rect 48833 12281 48845 12657
rect 48879 12281 48891 12657
rect 48833 12269 48891 12281
rect 48947 12657 49005 12669
rect 48947 12281 48959 12657
rect 48993 12281 49005 12657
rect 48947 12269 49005 12281
rect 49205 12657 49263 12669
rect 49205 12281 49217 12657
rect 49251 12281 49263 12657
rect 49205 12269 49263 12281
rect 49319 12657 49377 12669
rect 49319 12281 49331 12657
rect 49365 12281 49377 12657
rect 49319 12269 49377 12281
rect 49577 12657 49635 12669
rect 49577 12281 49589 12657
rect 49623 12281 49635 12657
rect 49577 12269 49635 12281
rect 49691 12657 49749 12669
rect 49691 12281 49703 12657
rect 49737 12281 49749 12657
rect 49691 12269 49749 12281
rect 49949 12657 50007 12669
rect 49949 12281 49961 12657
rect 49995 12281 50007 12657
rect 49949 12269 50007 12281
rect 50063 12657 50121 12669
rect 50063 12281 50075 12657
rect 50109 12281 50121 12657
rect 50063 12269 50121 12281
rect 50321 12657 50379 12669
rect 50321 12281 50333 12657
rect 50367 12281 50379 12657
rect 50321 12269 50379 12281
rect 50435 12657 50493 12669
rect 50435 12281 50447 12657
rect 50481 12281 50493 12657
rect 50435 12269 50493 12281
rect 50693 12657 50751 12669
rect 50693 12281 50705 12657
rect 50739 12281 50751 12657
rect 50693 12269 50751 12281
rect 50807 12657 50865 12669
rect 50807 12281 50819 12657
rect 50853 12281 50865 12657
rect 50807 12269 50865 12281
rect 51065 12657 51123 12669
rect 51065 12281 51077 12657
rect 51111 12281 51123 12657
rect 51065 12269 51123 12281
rect 39275 12021 39333 12033
rect 39275 11645 39287 12021
rect 39321 11645 39333 12021
rect 39275 11633 39333 11645
rect 39533 12021 39591 12033
rect 39533 11645 39545 12021
rect 39579 11645 39591 12021
rect 39533 11633 39591 11645
rect 39647 12021 39705 12033
rect 39647 11645 39659 12021
rect 39693 11645 39705 12021
rect 39647 11633 39705 11645
rect 39905 12021 39963 12033
rect 39905 11645 39917 12021
rect 39951 11645 39963 12021
rect 39905 11633 39963 11645
rect 40019 12021 40077 12033
rect 40019 11645 40031 12021
rect 40065 11645 40077 12021
rect 40019 11633 40077 11645
rect 40277 12021 40335 12033
rect 40277 11645 40289 12021
rect 40323 11645 40335 12021
rect 40277 11633 40335 11645
rect 40391 12021 40449 12033
rect 40391 11645 40403 12021
rect 40437 11645 40449 12021
rect 40391 11633 40449 11645
rect 40649 12021 40707 12033
rect 40649 11645 40661 12021
rect 40695 11645 40707 12021
rect 40649 11633 40707 11645
rect 40763 12021 40821 12033
rect 40763 11645 40775 12021
rect 40809 11645 40821 12021
rect 40763 11633 40821 11645
rect 41021 12021 41079 12033
rect 41021 11645 41033 12021
rect 41067 11645 41079 12021
rect 41021 11633 41079 11645
rect 41135 12021 41193 12033
rect 41135 11645 41147 12021
rect 41181 11645 41193 12021
rect 41135 11633 41193 11645
rect 41393 12021 41451 12033
rect 41393 11645 41405 12021
rect 41439 11645 41451 12021
rect 41393 11633 41451 11645
rect 41507 12021 41565 12033
rect 41507 11645 41519 12021
rect 41553 11645 41565 12021
rect 41507 11633 41565 11645
rect 41765 12021 41823 12033
rect 41765 11645 41777 12021
rect 41811 11645 41823 12021
rect 41765 11633 41823 11645
rect 41879 12021 41937 12033
rect 41879 11645 41891 12021
rect 41925 11645 41937 12021
rect 41879 11633 41937 11645
rect 42137 12021 42195 12033
rect 42137 11645 42149 12021
rect 42183 11645 42195 12021
rect 42137 11633 42195 11645
rect 42251 12021 42309 12033
rect 42251 11645 42263 12021
rect 42297 11645 42309 12021
rect 42251 11633 42309 11645
rect 42509 12021 42567 12033
rect 42509 11645 42521 12021
rect 42555 11645 42567 12021
rect 42509 11633 42567 11645
rect 42623 12021 42681 12033
rect 42623 11645 42635 12021
rect 42669 11645 42681 12021
rect 42623 11633 42681 11645
rect 42881 12021 42939 12033
rect 42881 11645 42893 12021
rect 42927 11645 42939 12021
rect 42881 11633 42939 11645
rect 42995 12021 43053 12033
rect 42995 11645 43007 12021
rect 43041 11645 43053 12021
rect 42995 11633 43053 11645
rect 43253 12021 43311 12033
rect 43253 11645 43265 12021
rect 43299 11645 43311 12021
rect 43253 11633 43311 11645
rect 43367 12021 43425 12033
rect 43367 11645 43379 12021
rect 43413 11645 43425 12021
rect 43367 11633 43425 11645
rect 43625 12021 43683 12033
rect 43625 11645 43637 12021
rect 43671 11645 43683 12021
rect 43625 11633 43683 11645
rect 43739 12021 43797 12033
rect 43739 11645 43751 12021
rect 43785 11645 43797 12021
rect 43739 11633 43797 11645
rect 43997 12021 44055 12033
rect 43997 11645 44009 12021
rect 44043 11645 44055 12021
rect 43997 11633 44055 11645
rect 44111 12021 44169 12033
rect 44111 11645 44123 12021
rect 44157 11645 44169 12021
rect 44111 11633 44169 11645
rect 44369 12021 44427 12033
rect 44369 11645 44381 12021
rect 44415 11645 44427 12021
rect 44369 11633 44427 11645
rect 44483 12021 44541 12033
rect 44483 11645 44495 12021
rect 44529 11645 44541 12021
rect 44483 11633 44541 11645
rect 44741 12021 44799 12033
rect 44741 11645 44753 12021
rect 44787 11645 44799 12021
rect 44741 11633 44799 11645
rect 44855 12021 44913 12033
rect 44855 11645 44867 12021
rect 44901 11645 44913 12021
rect 44855 11633 44913 11645
rect 45113 12021 45171 12033
rect 45113 11645 45125 12021
rect 45159 11645 45171 12021
rect 45113 11633 45171 11645
rect 45227 12021 45285 12033
rect 45227 11645 45239 12021
rect 45273 11645 45285 12021
rect 45227 11633 45285 11645
rect 45485 12021 45543 12033
rect 45485 11645 45497 12021
rect 45531 11645 45543 12021
rect 45485 11633 45543 11645
rect 45599 12021 45657 12033
rect 45599 11645 45611 12021
rect 45645 11645 45657 12021
rect 45599 11633 45657 11645
rect 45857 12021 45915 12033
rect 45857 11645 45869 12021
rect 45903 11645 45915 12021
rect 45857 11633 45915 11645
rect 45971 12021 46029 12033
rect 45971 11645 45983 12021
rect 46017 11645 46029 12021
rect 45971 11633 46029 11645
rect 46229 12021 46287 12033
rect 46229 11645 46241 12021
rect 46275 11645 46287 12021
rect 46229 11633 46287 11645
rect 46343 12021 46401 12033
rect 46343 11645 46355 12021
rect 46389 11645 46401 12021
rect 46343 11633 46401 11645
rect 46601 12021 46659 12033
rect 46601 11645 46613 12021
rect 46647 11645 46659 12021
rect 46601 11633 46659 11645
rect 46715 12021 46773 12033
rect 46715 11645 46727 12021
rect 46761 11645 46773 12021
rect 46715 11633 46773 11645
rect 46973 12021 47031 12033
rect 46973 11645 46985 12021
rect 47019 11645 47031 12021
rect 46973 11633 47031 11645
rect 47087 12021 47145 12033
rect 47087 11645 47099 12021
rect 47133 11645 47145 12021
rect 47087 11633 47145 11645
rect 47345 12021 47403 12033
rect 47345 11645 47357 12021
rect 47391 11645 47403 12021
rect 47345 11633 47403 11645
rect 47459 12021 47517 12033
rect 47459 11645 47471 12021
rect 47505 11645 47517 12021
rect 47459 11633 47517 11645
rect 47717 12021 47775 12033
rect 47717 11645 47729 12021
rect 47763 11645 47775 12021
rect 47717 11633 47775 11645
rect 47831 12021 47889 12033
rect 47831 11645 47843 12021
rect 47877 11645 47889 12021
rect 47831 11633 47889 11645
rect 48089 12021 48147 12033
rect 48089 11645 48101 12021
rect 48135 11645 48147 12021
rect 48089 11633 48147 11645
rect 48203 12021 48261 12033
rect 48203 11645 48215 12021
rect 48249 11645 48261 12021
rect 48203 11633 48261 11645
rect 48461 12021 48519 12033
rect 48461 11645 48473 12021
rect 48507 11645 48519 12021
rect 48461 11633 48519 11645
rect 48575 12021 48633 12033
rect 48575 11645 48587 12021
rect 48621 11645 48633 12021
rect 48575 11633 48633 11645
rect 48833 12021 48891 12033
rect 48833 11645 48845 12021
rect 48879 11645 48891 12021
rect 48833 11633 48891 11645
rect 48947 12021 49005 12033
rect 48947 11645 48959 12021
rect 48993 11645 49005 12021
rect 48947 11633 49005 11645
rect 49205 12021 49263 12033
rect 49205 11645 49217 12021
rect 49251 11645 49263 12021
rect 49205 11633 49263 11645
rect 49319 12021 49377 12033
rect 49319 11645 49331 12021
rect 49365 11645 49377 12021
rect 49319 11633 49377 11645
rect 49577 12021 49635 12033
rect 49577 11645 49589 12021
rect 49623 11645 49635 12021
rect 49577 11633 49635 11645
rect 49691 12021 49749 12033
rect 49691 11645 49703 12021
rect 49737 11645 49749 12021
rect 49691 11633 49749 11645
rect 49949 12021 50007 12033
rect 49949 11645 49961 12021
rect 49995 11645 50007 12021
rect 49949 11633 50007 11645
rect 50063 12021 50121 12033
rect 50063 11645 50075 12021
rect 50109 11645 50121 12021
rect 50063 11633 50121 11645
rect 50321 12021 50379 12033
rect 50321 11645 50333 12021
rect 50367 11645 50379 12021
rect 50321 11633 50379 11645
rect 50435 12021 50493 12033
rect 50435 11645 50447 12021
rect 50481 11645 50493 12021
rect 50435 11633 50493 11645
rect 50693 12021 50751 12033
rect 50693 11645 50705 12021
rect 50739 11645 50751 12021
rect 50693 11633 50751 11645
rect 50807 12021 50865 12033
rect 50807 11645 50819 12021
rect 50853 11645 50865 12021
rect 50807 11633 50865 11645
rect 51065 12021 51123 12033
rect 51065 11645 51077 12021
rect 51111 11645 51123 12021
rect 51065 11633 51123 11645
rect 39275 11385 39333 11397
rect 39275 11009 39287 11385
rect 39321 11009 39333 11385
rect 39275 10997 39333 11009
rect 39533 11385 39591 11397
rect 39533 11009 39545 11385
rect 39579 11009 39591 11385
rect 39533 10997 39591 11009
rect 39647 11385 39705 11397
rect 39647 11009 39659 11385
rect 39693 11009 39705 11385
rect 39647 10997 39705 11009
rect 39905 11385 39963 11397
rect 39905 11009 39917 11385
rect 39951 11009 39963 11385
rect 39905 10997 39963 11009
rect 40019 11385 40077 11397
rect 40019 11009 40031 11385
rect 40065 11009 40077 11385
rect 40019 10997 40077 11009
rect 40277 11385 40335 11397
rect 40277 11009 40289 11385
rect 40323 11009 40335 11385
rect 40277 10997 40335 11009
rect 40391 11385 40449 11397
rect 40391 11009 40403 11385
rect 40437 11009 40449 11385
rect 40391 10997 40449 11009
rect 40649 11385 40707 11397
rect 40649 11009 40661 11385
rect 40695 11009 40707 11385
rect 40649 10997 40707 11009
rect 40763 11385 40821 11397
rect 40763 11009 40775 11385
rect 40809 11009 40821 11385
rect 40763 10997 40821 11009
rect 41021 11385 41079 11397
rect 41021 11009 41033 11385
rect 41067 11009 41079 11385
rect 41021 10997 41079 11009
rect 41135 11385 41193 11397
rect 41135 11009 41147 11385
rect 41181 11009 41193 11385
rect 41135 10997 41193 11009
rect 41393 11385 41451 11397
rect 41393 11009 41405 11385
rect 41439 11009 41451 11385
rect 41393 10997 41451 11009
rect 41507 11385 41565 11397
rect 41507 11009 41519 11385
rect 41553 11009 41565 11385
rect 41507 10997 41565 11009
rect 41765 11385 41823 11397
rect 41765 11009 41777 11385
rect 41811 11009 41823 11385
rect 41765 10997 41823 11009
rect 41879 11385 41937 11397
rect 41879 11009 41891 11385
rect 41925 11009 41937 11385
rect 41879 10997 41937 11009
rect 42137 11385 42195 11397
rect 42137 11009 42149 11385
rect 42183 11009 42195 11385
rect 42137 10997 42195 11009
rect 42251 11385 42309 11397
rect 42251 11009 42263 11385
rect 42297 11009 42309 11385
rect 42251 10997 42309 11009
rect 42509 11385 42567 11397
rect 42509 11009 42521 11385
rect 42555 11009 42567 11385
rect 42509 10997 42567 11009
rect 42623 11385 42681 11397
rect 42623 11009 42635 11385
rect 42669 11009 42681 11385
rect 42623 10997 42681 11009
rect 42881 11385 42939 11397
rect 42881 11009 42893 11385
rect 42927 11009 42939 11385
rect 42881 10997 42939 11009
rect 42995 11385 43053 11397
rect 42995 11009 43007 11385
rect 43041 11009 43053 11385
rect 42995 10997 43053 11009
rect 43253 11385 43311 11397
rect 43253 11009 43265 11385
rect 43299 11009 43311 11385
rect 43253 10997 43311 11009
rect 43367 11385 43425 11397
rect 43367 11009 43379 11385
rect 43413 11009 43425 11385
rect 43367 10997 43425 11009
rect 43625 11385 43683 11397
rect 43625 11009 43637 11385
rect 43671 11009 43683 11385
rect 43625 10997 43683 11009
rect 43739 11385 43797 11397
rect 43739 11009 43751 11385
rect 43785 11009 43797 11385
rect 43739 10997 43797 11009
rect 43997 11385 44055 11397
rect 43997 11009 44009 11385
rect 44043 11009 44055 11385
rect 43997 10997 44055 11009
rect 44111 11385 44169 11397
rect 44111 11009 44123 11385
rect 44157 11009 44169 11385
rect 44111 10997 44169 11009
rect 44369 11385 44427 11397
rect 44369 11009 44381 11385
rect 44415 11009 44427 11385
rect 44369 10997 44427 11009
rect 44483 11385 44541 11397
rect 44483 11009 44495 11385
rect 44529 11009 44541 11385
rect 44483 10997 44541 11009
rect 44741 11385 44799 11397
rect 44741 11009 44753 11385
rect 44787 11009 44799 11385
rect 44741 10997 44799 11009
rect 44855 11385 44913 11397
rect 44855 11009 44867 11385
rect 44901 11009 44913 11385
rect 44855 10997 44913 11009
rect 45113 11385 45171 11397
rect 45113 11009 45125 11385
rect 45159 11009 45171 11385
rect 45113 10997 45171 11009
rect 45227 11385 45285 11397
rect 45227 11009 45239 11385
rect 45273 11009 45285 11385
rect 45227 10997 45285 11009
rect 45485 11385 45543 11397
rect 45485 11009 45497 11385
rect 45531 11009 45543 11385
rect 45485 10997 45543 11009
rect 45599 11385 45657 11397
rect 45599 11009 45611 11385
rect 45645 11009 45657 11385
rect 45599 10997 45657 11009
rect 45857 11385 45915 11397
rect 45857 11009 45869 11385
rect 45903 11009 45915 11385
rect 45857 10997 45915 11009
rect 45971 11385 46029 11397
rect 45971 11009 45983 11385
rect 46017 11009 46029 11385
rect 45971 10997 46029 11009
rect 46229 11385 46287 11397
rect 46229 11009 46241 11385
rect 46275 11009 46287 11385
rect 46229 10997 46287 11009
rect 46343 11385 46401 11397
rect 46343 11009 46355 11385
rect 46389 11009 46401 11385
rect 46343 10997 46401 11009
rect 46601 11385 46659 11397
rect 46601 11009 46613 11385
rect 46647 11009 46659 11385
rect 46601 10997 46659 11009
rect 46715 11385 46773 11397
rect 46715 11009 46727 11385
rect 46761 11009 46773 11385
rect 46715 10997 46773 11009
rect 46973 11385 47031 11397
rect 46973 11009 46985 11385
rect 47019 11009 47031 11385
rect 46973 10997 47031 11009
rect 47087 11385 47145 11397
rect 47087 11009 47099 11385
rect 47133 11009 47145 11385
rect 47087 10997 47145 11009
rect 47345 11385 47403 11397
rect 47345 11009 47357 11385
rect 47391 11009 47403 11385
rect 47345 10997 47403 11009
rect 47459 11385 47517 11397
rect 47459 11009 47471 11385
rect 47505 11009 47517 11385
rect 47459 10997 47517 11009
rect 47717 11385 47775 11397
rect 47717 11009 47729 11385
rect 47763 11009 47775 11385
rect 47717 10997 47775 11009
rect 47831 11385 47889 11397
rect 47831 11009 47843 11385
rect 47877 11009 47889 11385
rect 47831 10997 47889 11009
rect 48089 11385 48147 11397
rect 48089 11009 48101 11385
rect 48135 11009 48147 11385
rect 48089 10997 48147 11009
rect 48203 11385 48261 11397
rect 48203 11009 48215 11385
rect 48249 11009 48261 11385
rect 48203 10997 48261 11009
rect 48461 11385 48519 11397
rect 48461 11009 48473 11385
rect 48507 11009 48519 11385
rect 48461 10997 48519 11009
rect 48575 11385 48633 11397
rect 48575 11009 48587 11385
rect 48621 11009 48633 11385
rect 48575 10997 48633 11009
rect 48833 11385 48891 11397
rect 48833 11009 48845 11385
rect 48879 11009 48891 11385
rect 48833 10997 48891 11009
rect 48947 11385 49005 11397
rect 48947 11009 48959 11385
rect 48993 11009 49005 11385
rect 48947 10997 49005 11009
rect 49205 11385 49263 11397
rect 49205 11009 49217 11385
rect 49251 11009 49263 11385
rect 49205 10997 49263 11009
rect 49319 11385 49377 11397
rect 49319 11009 49331 11385
rect 49365 11009 49377 11385
rect 49319 10997 49377 11009
rect 49577 11385 49635 11397
rect 49577 11009 49589 11385
rect 49623 11009 49635 11385
rect 49577 10997 49635 11009
rect 49691 11385 49749 11397
rect 49691 11009 49703 11385
rect 49737 11009 49749 11385
rect 49691 10997 49749 11009
rect 49949 11385 50007 11397
rect 49949 11009 49961 11385
rect 49995 11009 50007 11385
rect 49949 10997 50007 11009
rect 50063 11385 50121 11397
rect 50063 11009 50075 11385
rect 50109 11009 50121 11385
rect 50063 10997 50121 11009
rect 50321 11385 50379 11397
rect 50321 11009 50333 11385
rect 50367 11009 50379 11385
rect 50321 10997 50379 11009
rect 50435 11385 50493 11397
rect 50435 11009 50447 11385
rect 50481 11009 50493 11385
rect 50435 10997 50493 11009
rect 50693 11385 50751 11397
rect 50693 11009 50705 11385
rect 50739 11009 50751 11385
rect 50693 10997 50751 11009
rect 50807 11385 50865 11397
rect 50807 11009 50819 11385
rect 50853 11009 50865 11385
rect 50807 10997 50865 11009
rect 51065 11385 51123 11397
rect 51065 11009 51077 11385
rect 51111 11009 51123 11385
rect 51065 10997 51123 11009
rect 39275 8856 39333 8868
rect 39275 8480 39287 8856
rect 39321 8480 39333 8856
rect 39275 8468 39333 8480
rect 39533 8856 39591 8868
rect 39533 8480 39545 8856
rect 39579 8480 39591 8856
rect 39533 8468 39591 8480
rect 39647 8856 39705 8868
rect 39647 8480 39659 8856
rect 39693 8480 39705 8856
rect 39647 8468 39705 8480
rect 39905 8856 39963 8868
rect 39905 8480 39917 8856
rect 39951 8480 39963 8856
rect 39905 8468 39963 8480
rect 40019 8856 40077 8868
rect 40019 8480 40031 8856
rect 40065 8480 40077 8856
rect 40019 8468 40077 8480
rect 40277 8856 40335 8868
rect 40277 8480 40289 8856
rect 40323 8480 40335 8856
rect 40277 8468 40335 8480
rect 40391 8856 40449 8868
rect 40391 8480 40403 8856
rect 40437 8480 40449 8856
rect 40391 8468 40449 8480
rect 40649 8856 40707 8868
rect 40649 8480 40661 8856
rect 40695 8480 40707 8856
rect 40649 8468 40707 8480
rect 40763 8856 40821 8868
rect 40763 8480 40775 8856
rect 40809 8480 40821 8856
rect 40763 8468 40821 8480
rect 41021 8856 41079 8868
rect 41021 8480 41033 8856
rect 41067 8480 41079 8856
rect 41021 8468 41079 8480
rect 41135 8856 41193 8868
rect 41135 8480 41147 8856
rect 41181 8480 41193 8856
rect 41135 8468 41193 8480
rect 41393 8856 41451 8868
rect 41393 8480 41405 8856
rect 41439 8480 41451 8856
rect 41393 8468 41451 8480
rect 41507 8856 41565 8868
rect 41507 8480 41519 8856
rect 41553 8480 41565 8856
rect 41507 8468 41565 8480
rect 41765 8856 41823 8868
rect 41765 8480 41777 8856
rect 41811 8480 41823 8856
rect 41765 8468 41823 8480
rect 41879 8856 41937 8868
rect 41879 8480 41891 8856
rect 41925 8480 41937 8856
rect 41879 8468 41937 8480
rect 42137 8856 42195 8868
rect 42137 8480 42149 8856
rect 42183 8480 42195 8856
rect 42137 8468 42195 8480
rect 42251 8856 42309 8868
rect 42251 8480 42263 8856
rect 42297 8480 42309 8856
rect 42251 8468 42309 8480
rect 42509 8856 42567 8868
rect 42509 8480 42521 8856
rect 42555 8480 42567 8856
rect 42509 8468 42567 8480
rect 42623 8856 42681 8868
rect 42623 8480 42635 8856
rect 42669 8480 42681 8856
rect 42623 8468 42681 8480
rect 42881 8856 42939 8868
rect 42881 8480 42893 8856
rect 42927 8480 42939 8856
rect 42881 8468 42939 8480
rect 42995 8856 43053 8868
rect 42995 8480 43007 8856
rect 43041 8480 43053 8856
rect 42995 8468 43053 8480
rect 43253 8856 43311 8868
rect 43253 8480 43265 8856
rect 43299 8480 43311 8856
rect 43253 8468 43311 8480
rect 43367 8856 43425 8868
rect 43367 8480 43379 8856
rect 43413 8480 43425 8856
rect 43367 8468 43425 8480
rect 43625 8856 43683 8868
rect 43625 8480 43637 8856
rect 43671 8480 43683 8856
rect 43625 8468 43683 8480
rect 43739 8856 43797 8868
rect 43739 8480 43751 8856
rect 43785 8480 43797 8856
rect 43739 8468 43797 8480
rect 43997 8856 44055 8868
rect 43997 8480 44009 8856
rect 44043 8480 44055 8856
rect 43997 8468 44055 8480
rect 44111 8856 44169 8868
rect 44111 8480 44123 8856
rect 44157 8480 44169 8856
rect 44111 8468 44169 8480
rect 44369 8856 44427 8868
rect 44369 8480 44381 8856
rect 44415 8480 44427 8856
rect 44369 8468 44427 8480
rect 44483 8856 44541 8868
rect 44483 8480 44495 8856
rect 44529 8480 44541 8856
rect 44483 8468 44541 8480
rect 44741 8856 44799 8868
rect 44741 8480 44753 8856
rect 44787 8480 44799 8856
rect 44741 8468 44799 8480
rect 44855 8856 44913 8868
rect 44855 8480 44867 8856
rect 44901 8480 44913 8856
rect 44855 8468 44913 8480
rect 45113 8856 45171 8868
rect 45113 8480 45125 8856
rect 45159 8480 45171 8856
rect 45113 8468 45171 8480
rect 45227 8856 45285 8868
rect 45227 8480 45239 8856
rect 45273 8480 45285 8856
rect 45227 8468 45285 8480
rect 45485 8856 45543 8868
rect 45485 8480 45497 8856
rect 45531 8480 45543 8856
rect 45485 8468 45543 8480
rect 45599 8856 45657 8868
rect 45599 8480 45611 8856
rect 45645 8480 45657 8856
rect 45599 8468 45657 8480
rect 45857 8856 45915 8868
rect 45857 8480 45869 8856
rect 45903 8480 45915 8856
rect 45857 8468 45915 8480
rect 45971 8856 46029 8868
rect 45971 8480 45983 8856
rect 46017 8480 46029 8856
rect 45971 8468 46029 8480
rect 46229 8856 46287 8868
rect 46229 8480 46241 8856
rect 46275 8480 46287 8856
rect 46229 8468 46287 8480
rect 46343 8856 46401 8868
rect 46343 8480 46355 8856
rect 46389 8480 46401 8856
rect 46343 8468 46401 8480
rect 46601 8856 46659 8868
rect 46601 8480 46613 8856
rect 46647 8480 46659 8856
rect 46601 8468 46659 8480
rect 46715 8856 46773 8868
rect 46715 8480 46727 8856
rect 46761 8480 46773 8856
rect 46715 8468 46773 8480
rect 46973 8856 47031 8868
rect 46973 8480 46985 8856
rect 47019 8480 47031 8856
rect 46973 8468 47031 8480
rect 47087 8856 47145 8868
rect 47087 8480 47099 8856
rect 47133 8480 47145 8856
rect 47087 8468 47145 8480
rect 47345 8856 47403 8868
rect 47345 8480 47357 8856
rect 47391 8480 47403 8856
rect 47345 8468 47403 8480
rect 47459 8856 47517 8868
rect 47459 8480 47471 8856
rect 47505 8480 47517 8856
rect 47459 8468 47517 8480
rect 47717 8856 47775 8868
rect 47717 8480 47729 8856
rect 47763 8480 47775 8856
rect 47717 8468 47775 8480
rect 47831 8856 47889 8868
rect 47831 8480 47843 8856
rect 47877 8480 47889 8856
rect 47831 8468 47889 8480
rect 48089 8856 48147 8868
rect 48089 8480 48101 8856
rect 48135 8480 48147 8856
rect 48089 8468 48147 8480
rect 48203 8856 48261 8868
rect 48203 8480 48215 8856
rect 48249 8480 48261 8856
rect 48203 8468 48261 8480
rect 48461 8856 48519 8868
rect 48461 8480 48473 8856
rect 48507 8480 48519 8856
rect 48461 8468 48519 8480
rect 48575 8856 48633 8868
rect 48575 8480 48587 8856
rect 48621 8480 48633 8856
rect 48575 8468 48633 8480
rect 48833 8856 48891 8868
rect 48833 8480 48845 8856
rect 48879 8480 48891 8856
rect 48833 8468 48891 8480
rect 48947 8856 49005 8868
rect 48947 8480 48959 8856
rect 48993 8480 49005 8856
rect 48947 8468 49005 8480
rect 49205 8856 49263 8868
rect 49205 8480 49217 8856
rect 49251 8480 49263 8856
rect 49205 8468 49263 8480
rect 49319 8856 49377 8868
rect 49319 8480 49331 8856
rect 49365 8480 49377 8856
rect 49319 8468 49377 8480
rect 49577 8856 49635 8868
rect 49577 8480 49589 8856
rect 49623 8480 49635 8856
rect 49577 8468 49635 8480
rect 49691 8856 49749 8868
rect 49691 8480 49703 8856
rect 49737 8480 49749 8856
rect 49691 8468 49749 8480
rect 49949 8856 50007 8868
rect 49949 8480 49961 8856
rect 49995 8480 50007 8856
rect 49949 8468 50007 8480
rect 50063 8856 50121 8868
rect 50063 8480 50075 8856
rect 50109 8480 50121 8856
rect 50063 8468 50121 8480
rect 50321 8856 50379 8868
rect 50321 8480 50333 8856
rect 50367 8480 50379 8856
rect 50321 8468 50379 8480
rect 50435 8856 50493 8868
rect 50435 8480 50447 8856
rect 50481 8480 50493 8856
rect 50435 8468 50493 8480
rect 50693 8856 50751 8868
rect 50693 8480 50705 8856
rect 50739 8480 50751 8856
rect 50693 8468 50751 8480
rect 50807 8856 50865 8868
rect 50807 8480 50819 8856
rect 50853 8480 50865 8856
rect 50807 8468 50865 8480
rect 51065 8856 51123 8868
rect 51065 8480 51077 8856
rect 51111 8480 51123 8856
rect 51065 8468 51123 8480
rect 39275 8220 39333 8232
rect 39275 7844 39287 8220
rect 39321 7844 39333 8220
rect 39275 7832 39333 7844
rect 39533 8220 39591 8232
rect 39533 7844 39545 8220
rect 39579 7844 39591 8220
rect 39533 7832 39591 7844
rect 39647 8220 39705 8232
rect 39647 7844 39659 8220
rect 39693 7844 39705 8220
rect 39647 7832 39705 7844
rect 39905 8220 39963 8232
rect 39905 7844 39917 8220
rect 39951 7844 39963 8220
rect 39905 7832 39963 7844
rect 40019 8220 40077 8232
rect 40019 7844 40031 8220
rect 40065 7844 40077 8220
rect 40019 7832 40077 7844
rect 40277 8220 40335 8232
rect 40277 7844 40289 8220
rect 40323 7844 40335 8220
rect 40277 7832 40335 7844
rect 40391 8220 40449 8232
rect 40391 7844 40403 8220
rect 40437 7844 40449 8220
rect 40391 7832 40449 7844
rect 40649 8220 40707 8232
rect 40649 7844 40661 8220
rect 40695 7844 40707 8220
rect 40649 7832 40707 7844
rect 40763 8220 40821 8232
rect 40763 7844 40775 8220
rect 40809 7844 40821 8220
rect 40763 7832 40821 7844
rect 41021 8220 41079 8232
rect 41021 7844 41033 8220
rect 41067 7844 41079 8220
rect 41021 7832 41079 7844
rect 41135 8220 41193 8232
rect 41135 7844 41147 8220
rect 41181 7844 41193 8220
rect 41135 7832 41193 7844
rect 41393 8220 41451 8232
rect 41393 7844 41405 8220
rect 41439 7844 41451 8220
rect 41393 7832 41451 7844
rect 41507 8220 41565 8232
rect 41507 7844 41519 8220
rect 41553 7844 41565 8220
rect 41507 7832 41565 7844
rect 41765 8220 41823 8232
rect 41765 7844 41777 8220
rect 41811 7844 41823 8220
rect 41765 7832 41823 7844
rect 41879 8220 41937 8232
rect 41879 7844 41891 8220
rect 41925 7844 41937 8220
rect 41879 7832 41937 7844
rect 42137 8220 42195 8232
rect 42137 7844 42149 8220
rect 42183 7844 42195 8220
rect 42137 7832 42195 7844
rect 42251 8220 42309 8232
rect 42251 7844 42263 8220
rect 42297 7844 42309 8220
rect 42251 7832 42309 7844
rect 42509 8220 42567 8232
rect 42509 7844 42521 8220
rect 42555 7844 42567 8220
rect 42509 7832 42567 7844
rect 42623 8220 42681 8232
rect 42623 7844 42635 8220
rect 42669 7844 42681 8220
rect 42623 7832 42681 7844
rect 42881 8220 42939 8232
rect 42881 7844 42893 8220
rect 42927 7844 42939 8220
rect 42881 7832 42939 7844
rect 42995 8220 43053 8232
rect 42995 7844 43007 8220
rect 43041 7844 43053 8220
rect 42995 7832 43053 7844
rect 43253 8220 43311 8232
rect 43253 7844 43265 8220
rect 43299 7844 43311 8220
rect 43253 7832 43311 7844
rect 43367 8220 43425 8232
rect 43367 7844 43379 8220
rect 43413 7844 43425 8220
rect 43367 7832 43425 7844
rect 43625 8220 43683 8232
rect 43625 7844 43637 8220
rect 43671 7844 43683 8220
rect 43625 7832 43683 7844
rect 43739 8220 43797 8232
rect 43739 7844 43751 8220
rect 43785 7844 43797 8220
rect 43739 7832 43797 7844
rect 43997 8220 44055 8232
rect 43997 7844 44009 8220
rect 44043 7844 44055 8220
rect 43997 7832 44055 7844
rect 44111 8220 44169 8232
rect 44111 7844 44123 8220
rect 44157 7844 44169 8220
rect 44111 7832 44169 7844
rect 44369 8220 44427 8232
rect 44369 7844 44381 8220
rect 44415 7844 44427 8220
rect 44369 7832 44427 7844
rect 44483 8220 44541 8232
rect 44483 7844 44495 8220
rect 44529 7844 44541 8220
rect 44483 7832 44541 7844
rect 44741 8220 44799 8232
rect 44741 7844 44753 8220
rect 44787 7844 44799 8220
rect 44741 7832 44799 7844
rect 44855 8220 44913 8232
rect 44855 7844 44867 8220
rect 44901 7844 44913 8220
rect 44855 7832 44913 7844
rect 45113 8220 45171 8232
rect 45113 7844 45125 8220
rect 45159 7844 45171 8220
rect 45113 7832 45171 7844
rect 45227 8220 45285 8232
rect 45227 7844 45239 8220
rect 45273 7844 45285 8220
rect 45227 7832 45285 7844
rect 45485 8220 45543 8232
rect 45485 7844 45497 8220
rect 45531 7844 45543 8220
rect 45485 7832 45543 7844
rect 45599 8220 45657 8232
rect 45599 7844 45611 8220
rect 45645 7844 45657 8220
rect 45599 7832 45657 7844
rect 45857 8220 45915 8232
rect 45857 7844 45869 8220
rect 45903 7844 45915 8220
rect 45857 7832 45915 7844
rect 45971 8220 46029 8232
rect 45971 7844 45983 8220
rect 46017 7844 46029 8220
rect 45971 7832 46029 7844
rect 46229 8220 46287 8232
rect 46229 7844 46241 8220
rect 46275 7844 46287 8220
rect 46229 7832 46287 7844
rect 46343 8220 46401 8232
rect 46343 7844 46355 8220
rect 46389 7844 46401 8220
rect 46343 7832 46401 7844
rect 46601 8220 46659 8232
rect 46601 7844 46613 8220
rect 46647 7844 46659 8220
rect 46601 7832 46659 7844
rect 46715 8220 46773 8232
rect 46715 7844 46727 8220
rect 46761 7844 46773 8220
rect 46715 7832 46773 7844
rect 46973 8220 47031 8232
rect 46973 7844 46985 8220
rect 47019 7844 47031 8220
rect 46973 7832 47031 7844
rect 47087 8220 47145 8232
rect 47087 7844 47099 8220
rect 47133 7844 47145 8220
rect 47087 7832 47145 7844
rect 47345 8220 47403 8232
rect 47345 7844 47357 8220
rect 47391 7844 47403 8220
rect 47345 7832 47403 7844
rect 47459 8220 47517 8232
rect 47459 7844 47471 8220
rect 47505 7844 47517 8220
rect 47459 7832 47517 7844
rect 47717 8220 47775 8232
rect 47717 7844 47729 8220
rect 47763 7844 47775 8220
rect 47717 7832 47775 7844
rect 47831 8220 47889 8232
rect 47831 7844 47843 8220
rect 47877 7844 47889 8220
rect 47831 7832 47889 7844
rect 48089 8220 48147 8232
rect 48089 7844 48101 8220
rect 48135 7844 48147 8220
rect 48089 7832 48147 7844
rect 48203 8220 48261 8232
rect 48203 7844 48215 8220
rect 48249 7844 48261 8220
rect 48203 7832 48261 7844
rect 48461 8220 48519 8232
rect 48461 7844 48473 8220
rect 48507 7844 48519 8220
rect 48461 7832 48519 7844
rect 48575 8220 48633 8232
rect 48575 7844 48587 8220
rect 48621 7844 48633 8220
rect 48575 7832 48633 7844
rect 48833 8220 48891 8232
rect 48833 7844 48845 8220
rect 48879 7844 48891 8220
rect 48833 7832 48891 7844
rect 48947 8220 49005 8232
rect 48947 7844 48959 8220
rect 48993 7844 49005 8220
rect 48947 7832 49005 7844
rect 49205 8220 49263 8232
rect 49205 7844 49217 8220
rect 49251 7844 49263 8220
rect 49205 7832 49263 7844
rect 49319 8220 49377 8232
rect 49319 7844 49331 8220
rect 49365 7844 49377 8220
rect 49319 7832 49377 7844
rect 49577 8220 49635 8232
rect 49577 7844 49589 8220
rect 49623 7844 49635 8220
rect 49577 7832 49635 7844
rect 49691 8220 49749 8232
rect 49691 7844 49703 8220
rect 49737 7844 49749 8220
rect 49691 7832 49749 7844
rect 49949 8220 50007 8232
rect 49949 7844 49961 8220
rect 49995 7844 50007 8220
rect 49949 7832 50007 7844
rect 50063 8220 50121 8232
rect 50063 7844 50075 8220
rect 50109 7844 50121 8220
rect 50063 7832 50121 7844
rect 50321 8220 50379 8232
rect 50321 7844 50333 8220
rect 50367 7844 50379 8220
rect 50321 7832 50379 7844
rect 50435 8220 50493 8232
rect 50435 7844 50447 8220
rect 50481 7844 50493 8220
rect 50435 7832 50493 7844
rect 50693 8220 50751 8232
rect 50693 7844 50705 8220
rect 50739 7844 50751 8220
rect 50693 7832 50751 7844
rect 50807 8220 50865 8232
rect 50807 7844 50819 8220
rect 50853 7844 50865 8220
rect 50807 7832 50865 7844
rect 51065 8220 51123 8232
rect 51065 7844 51077 8220
rect 51111 7844 51123 8220
rect 51065 7832 51123 7844
rect 39275 7584 39333 7596
rect 39275 7208 39287 7584
rect 39321 7208 39333 7584
rect 39275 7196 39333 7208
rect 39533 7584 39591 7596
rect 39533 7208 39545 7584
rect 39579 7208 39591 7584
rect 39533 7196 39591 7208
rect 39647 7584 39705 7596
rect 39647 7208 39659 7584
rect 39693 7208 39705 7584
rect 39647 7196 39705 7208
rect 39905 7584 39963 7596
rect 39905 7208 39917 7584
rect 39951 7208 39963 7584
rect 39905 7196 39963 7208
rect 40019 7584 40077 7596
rect 40019 7208 40031 7584
rect 40065 7208 40077 7584
rect 40019 7196 40077 7208
rect 40277 7584 40335 7596
rect 40277 7208 40289 7584
rect 40323 7208 40335 7584
rect 40277 7196 40335 7208
rect 40391 7584 40449 7596
rect 40391 7208 40403 7584
rect 40437 7208 40449 7584
rect 40391 7196 40449 7208
rect 40649 7584 40707 7596
rect 40649 7208 40661 7584
rect 40695 7208 40707 7584
rect 40649 7196 40707 7208
rect 40763 7584 40821 7596
rect 40763 7208 40775 7584
rect 40809 7208 40821 7584
rect 40763 7196 40821 7208
rect 41021 7584 41079 7596
rect 41021 7208 41033 7584
rect 41067 7208 41079 7584
rect 41021 7196 41079 7208
rect 41135 7584 41193 7596
rect 41135 7208 41147 7584
rect 41181 7208 41193 7584
rect 41135 7196 41193 7208
rect 41393 7584 41451 7596
rect 41393 7208 41405 7584
rect 41439 7208 41451 7584
rect 41393 7196 41451 7208
rect 41507 7584 41565 7596
rect 41507 7208 41519 7584
rect 41553 7208 41565 7584
rect 41507 7196 41565 7208
rect 41765 7584 41823 7596
rect 41765 7208 41777 7584
rect 41811 7208 41823 7584
rect 41765 7196 41823 7208
rect 41879 7584 41937 7596
rect 41879 7208 41891 7584
rect 41925 7208 41937 7584
rect 41879 7196 41937 7208
rect 42137 7584 42195 7596
rect 42137 7208 42149 7584
rect 42183 7208 42195 7584
rect 42137 7196 42195 7208
rect 42251 7584 42309 7596
rect 42251 7208 42263 7584
rect 42297 7208 42309 7584
rect 42251 7196 42309 7208
rect 42509 7584 42567 7596
rect 42509 7208 42521 7584
rect 42555 7208 42567 7584
rect 42509 7196 42567 7208
rect 42623 7584 42681 7596
rect 42623 7208 42635 7584
rect 42669 7208 42681 7584
rect 42623 7196 42681 7208
rect 42881 7584 42939 7596
rect 42881 7208 42893 7584
rect 42927 7208 42939 7584
rect 42881 7196 42939 7208
rect 42995 7584 43053 7596
rect 42995 7208 43007 7584
rect 43041 7208 43053 7584
rect 42995 7196 43053 7208
rect 43253 7584 43311 7596
rect 43253 7208 43265 7584
rect 43299 7208 43311 7584
rect 43253 7196 43311 7208
rect 43367 7584 43425 7596
rect 43367 7208 43379 7584
rect 43413 7208 43425 7584
rect 43367 7196 43425 7208
rect 43625 7584 43683 7596
rect 43625 7208 43637 7584
rect 43671 7208 43683 7584
rect 43625 7196 43683 7208
rect 43739 7584 43797 7596
rect 43739 7208 43751 7584
rect 43785 7208 43797 7584
rect 43739 7196 43797 7208
rect 43997 7584 44055 7596
rect 43997 7208 44009 7584
rect 44043 7208 44055 7584
rect 43997 7196 44055 7208
rect 44111 7584 44169 7596
rect 44111 7208 44123 7584
rect 44157 7208 44169 7584
rect 44111 7196 44169 7208
rect 44369 7584 44427 7596
rect 44369 7208 44381 7584
rect 44415 7208 44427 7584
rect 44369 7196 44427 7208
rect 44483 7584 44541 7596
rect 44483 7208 44495 7584
rect 44529 7208 44541 7584
rect 44483 7196 44541 7208
rect 44741 7584 44799 7596
rect 44741 7208 44753 7584
rect 44787 7208 44799 7584
rect 44741 7196 44799 7208
rect 44855 7584 44913 7596
rect 44855 7208 44867 7584
rect 44901 7208 44913 7584
rect 44855 7196 44913 7208
rect 45113 7584 45171 7596
rect 45113 7208 45125 7584
rect 45159 7208 45171 7584
rect 45113 7196 45171 7208
rect 45227 7584 45285 7596
rect 45227 7208 45239 7584
rect 45273 7208 45285 7584
rect 45227 7196 45285 7208
rect 45485 7584 45543 7596
rect 45485 7208 45497 7584
rect 45531 7208 45543 7584
rect 45485 7196 45543 7208
rect 45599 7584 45657 7596
rect 45599 7208 45611 7584
rect 45645 7208 45657 7584
rect 45599 7196 45657 7208
rect 45857 7584 45915 7596
rect 45857 7208 45869 7584
rect 45903 7208 45915 7584
rect 45857 7196 45915 7208
rect 45971 7584 46029 7596
rect 45971 7208 45983 7584
rect 46017 7208 46029 7584
rect 45971 7196 46029 7208
rect 46229 7584 46287 7596
rect 46229 7208 46241 7584
rect 46275 7208 46287 7584
rect 46229 7196 46287 7208
rect 46343 7584 46401 7596
rect 46343 7208 46355 7584
rect 46389 7208 46401 7584
rect 46343 7196 46401 7208
rect 46601 7584 46659 7596
rect 46601 7208 46613 7584
rect 46647 7208 46659 7584
rect 46601 7196 46659 7208
rect 46715 7584 46773 7596
rect 46715 7208 46727 7584
rect 46761 7208 46773 7584
rect 46715 7196 46773 7208
rect 46973 7584 47031 7596
rect 46973 7208 46985 7584
rect 47019 7208 47031 7584
rect 46973 7196 47031 7208
rect 47087 7584 47145 7596
rect 47087 7208 47099 7584
rect 47133 7208 47145 7584
rect 47087 7196 47145 7208
rect 47345 7584 47403 7596
rect 47345 7208 47357 7584
rect 47391 7208 47403 7584
rect 47345 7196 47403 7208
rect 47459 7584 47517 7596
rect 47459 7208 47471 7584
rect 47505 7208 47517 7584
rect 47459 7196 47517 7208
rect 47717 7584 47775 7596
rect 47717 7208 47729 7584
rect 47763 7208 47775 7584
rect 47717 7196 47775 7208
rect 47831 7584 47889 7596
rect 47831 7208 47843 7584
rect 47877 7208 47889 7584
rect 47831 7196 47889 7208
rect 48089 7584 48147 7596
rect 48089 7208 48101 7584
rect 48135 7208 48147 7584
rect 48089 7196 48147 7208
rect 48203 7584 48261 7596
rect 48203 7208 48215 7584
rect 48249 7208 48261 7584
rect 48203 7196 48261 7208
rect 48461 7584 48519 7596
rect 48461 7208 48473 7584
rect 48507 7208 48519 7584
rect 48461 7196 48519 7208
rect 48575 7584 48633 7596
rect 48575 7208 48587 7584
rect 48621 7208 48633 7584
rect 48575 7196 48633 7208
rect 48833 7584 48891 7596
rect 48833 7208 48845 7584
rect 48879 7208 48891 7584
rect 48833 7196 48891 7208
rect 48947 7584 49005 7596
rect 48947 7208 48959 7584
rect 48993 7208 49005 7584
rect 48947 7196 49005 7208
rect 49205 7584 49263 7596
rect 49205 7208 49217 7584
rect 49251 7208 49263 7584
rect 49205 7196 49263 7208
rect 49319 7584 49377 7596
rect 49319 7208 49331 7584
rect 49365 7208 49377 7584
rect 49319 7196 49377 7208
rect 49577 7584 49635 7596
rect 49577 7208 49589 7584
rect 49623 7208 49635 7584
rect 49577 7196 49635 7208
rect 49691 7584 49749 7596
rect 49691 7208 49703 7584
rect 49737 7208 49749 7584
rect 49691 7196 49749 7208
rect 49949 7584 50007 7596
rect 49949 7208 49961 7584
rect 49995 7208 50007 7584
rect 49949 7196 50007 7208
rect 50063 7584 50121 7596
rect 50063 7208 50075 7584
rect 50109 7208 50121 7584
rect 50063 7196 50121 7208
rect 50321 7584 50379 7596
rect 50321 7208 50333 7584
rect 50367 7208 50379 7584
rect 50321 7196 50379 7208
rect 50435 7584 50493 7596
rect 50435 7208 50447 7584
rect 50481 7208 50493 7584
rect 50435 7196 50493 7208
rect 50693 7584 50751 7596
rect 50693 7208 50705 7584
rect 50739 7208 50751 7584
rect 50693 7196 50751 7208
rect 50807 7584 50865 7596
rect 50807 7208 50819 7584
rect 50853 7208 50865 7584
rect 50807 7196 50865 7208
rect 51065 7584 51123 7596
rect 51065 7208 51077 7584
rect 51111 7208 51123 7584
rect 51065 7196 51123 7208
rect 40763 6468 40821 6480
rect 40763 5692 40775 6468
rect 40809 5692 40821 6468
rect 40763 5680 40821 5692
rect 41021 6468 41079 6480
rect 41021 5692 41033 6468
rect 41067 5692 41079 6468
rect 41021 5680 41079 5692
rect 41135 6468 41193 6480
rect 41135 5692 41147 6468
rect 41181 5692 41193 6468
rect 41135 5680 41193 5692
rect 41393 6468 41451 6480
rect 41393 5692 41405 6468
rect 41439 5692 41451 6468
rect 41393 5680 41451 5692
rect 41507 6468 41565 6480
rect 41507 5692 41519 6468
rect 41553 5692 41565 6468
rect 41507 5680 41565 5692
rect 41765 6468 41823 6480
rect 41765 5692 41777 6468
rect 41811 5692 41823 6468
rect 41765 5680 41823 5692
rect 41879 6468 41937 6480
rect 41879 5692 41891 6468
rect 41925 5692 41937 6468
rect 41879 5680 41937 5692
rect 42137 6468 42195 6480
rect 42137 5692 42149 6468
rect 42183 5692 42195 6468
rect 42137 5680 42195 5692
rect 42251 6468 42309 6480
rect 42251 5692 42263 6468
rect 42297 5692 42309 6468
rect 42251 5680 42309 5692
rect 42509 6468 42567 6480
rect 42509 5692 42521 6468
rect 42555 5692 42567 6468
rect 42509 5680 42567 5692
rect 42623 6468 42681 6480
rect 42623 5692 42635 6468
rect 42669 5692 42681 6468
rect 42623 5680 42681 5692
rect 42881 6468 42939 6480
rect 42881 5692 42893 6468
rect 42927 5692 42939 6468
rect 42881 5680 42939 5692
rect 42995 6468 43053 6480
rect 42995 5692 43007 6468
rect 43041 5692 43053 6468
rect 42995 5680 43053 5692
rect 43253 6468 43311 6480
rect 43253 5692 43265 6468
rect 43299 5692 43311 6468
rect 43253 5680 43311 5692
rect 43367 6468 43425 6480
rect 43367 5692 43379 6468
rect 43413 5692 43425 6468
rect 43367 5680 43425 5692
rect 43625 6468 43683 6480
rect 43625 5692 43637 6468
rect 43671 5692 43683 6468
rect 43625 5680 43683 5692
rect 40763 5432 40821 5444
rect 40763 4656 40775 5432
rect 40809 4656 40821 5432
rect 40763 4644 40821 4656
rect 41021 5432 41079 5444
rect 41021 4656 41033 5432
rect 41067 4656 41079 5432
rect 41021 4644 41079 4656
rect 41135 5432 41193 5444
rect 41135 4656 41147 5432
rect 41181 4656 41193 5432
rect 41135 4644 41193 4656
rect 41393 5432 41451 5444
rect 41393 4656 41405 5432
rect 41439 4656 41451 5432
rect 41393 4644 41451 4656
rect 41507 5432 41565 5444
rect 41507 4656 41519 5432
rect 41553 4656 41565 5432
rect 41507 4644 41565 4656
rect 41765 5432 41823 5444
rect 41765 4656 41777 5432
rect 41811 4656 41823 5432
rect 41765 4644 41823 4656
rect 41879 5432 41937 5444
rect 41879 4656 41891 5432
rect 41925 4656 41937 5432
rect 41879 4644 41937 4656
rect 42137 5432 42195 5444
rect 42137 4656 42149 5432
rect 42183 4656 42195 5432
rect 42137 4644 42195 4656
rect 42251 5432 42309 5444
rect 42251 4656 42263 5432
rect 42297 4656 42309 5432
rect 42251 4644 42309 4656
rect 42509 5432 42567 5444
rect 42509 4656 42521 5432
rect 42555 4656 42567 5432
rect 42509 4644 42567 4656
rect 42623 5432 42681 5444
rect 42623 4656 42635 5432
rect 42669 4656 42681 5432
rect 42623 4644 42681 4656
rect 42881 5432 42939 5444
rect 42881 4656 42893 5432
rect 42927 4656 42939 5432
rect 42881 4644 42939 4656
rect 42995 5432 43053 5444
rect 42995 4656 43007 5432
rect 43041 4656 43053 5432
rect 42995 4644 43053 4656
rect 43253 5432 43311 5444
rect 43253 4656 43265 5432
rect 43299 4656 43311 5432
rect 43253 4644 43311 4656
rect 43367 5432 43425 5444
rect 43367 4656 43379 5432
rect 43413 4656 43425 5432
rect 43367 4644 43425 4656
rect 43625 5432 43683 5444
rect 43625 4656 43637 5432
rect 43671 4656 43683 5432
rect 43625 4644 43683 4656
rect 40763 4396 40821 4408
rect 40763 3620 40775 4396
rect 40809 3620 40821 4396
rect 40763 3608 40821 3620
rect 41021 4396 41079 4408
rect 41021 3620 41033 4396
rect 41067 3620 41079 4396
rect 41021 3608 41079 3620
rect 41135 4396 41193 4408
rect 41135 3620 41147 4396
rect 41181 3620 41193 4396
rect 41135 3608 41193 3620
rect 41393 4396 41451 4408
rect 41393 3620 41405 4396
rect 41439 3620 41451 4396
rect 41393 3608 41451 3620
rect 41507 4396 41565 4408
rect 41507 3620 41519 4396
rect 41553 3620 41565 4396
rect 41507 3608 41565 3620
rect 41765 4396 41823 4408
rect 41765 3620 41777 4396
rect 41811 3620 41823 4396
rect 41765 3608 41823 3620
rect 41879 4396 41937 4408
rect 41879 3620 41891 4396
rect 41925 3620 41937 4396
rect 41879 3608 41937 3620
rect 42137 4396 42195 4408
rect 42137 3620 42149 4396
rect 42183 3620 42195 4396
rect 42137 3608 42195 3620
rect 42251 4396 42309 4408
rect 42251 3620 42263 4396
rect 42297 3620 42309 4396
rect 42251 3608 42309 3620
rect 42509 4396 42567 4408
rect 42509 3620 42521 4396
rect 42555 3620 42567 4396
rect 42509 3608 42567 3620
rect 42623 4396 42681 4408
rect 42623 3620 42635 4396
rect 42669 3620 42681 4396
rect 42623 3608 42681 3620
rect 42881 4396 42939 4408
rect 42881 3620 42893 4396
rect 42927 3620 42939 4396
rect 42881 3608 42939 3620
rect 42995 4396 43053 4408
rect 42995 3620 43007 4396
rect 43041 3620 43053 4396
rect 42995 3608 43053 3620
rect 43253 4396 43311 4408
rect 43253 3620 43265 4396
rect 43299 3620 43311 4396
rect 43253 3608 43311 3620
rect 43367 4396 43425 4408
rect 43367 3620 43379 4396
rect 43413 3620 43425 4396
rect 43367 3608 43425 3620
rect 43625 4396 43683 4408
rect 43625 3620 43637 4396
rect 43671 3620 43683 4396
rect 43625 3608 43683 3620
rect 40763 3360 40821 3372
rect 40763 2584 40775 3360
rect 40809 2584 40821 3360
rect 40763 2572 40821 2584
rect 41021 3360 41079 3372
rect 41021 2584 41033 3360
rect 41067 2584 41079 3360
rect 41021 2572 41079 2584
rect 41135 3360 41193 3372
rect 41135 2584 41147 3360
rect 41181 2584 41193 3360
rect 41135 2572 41193 2584
rect 41393 3360 41451 3372
rect 41393 2584 41405 3360
rect 41439 2584 41451 3360
rect 41393 2572 41451 2584
rect 41507 3360 41565 3372
rect 41507 2584 41519 3360
rect 41553 2584 41565 3360
rect 41507 2572 41565 2584
rect 41765 3360 41823 3372
rect 41765 2584 41777 3360
rect 41811 2584 41823 3360
rect 41765 2572 41823 2584
rect 41879 3360 41937 3372
rect 41879 2584 41891 3360
rect 41925 2584 41937 3360
rect 41879 2572 41937 2584
rect 42137 3360 42195 3372
rect 42137 2584 42149 3360
rect 42183 2584 42195 3360
rect 42137 2572 42195 2584
rect 42251 3360 42309 3372
rect 42251 2584 42263 3360
rect 42297 2584 42309 3360
rect 42251 2572 42309 2584
rect 42509 3360 42567 3372
rect 42509 2584 42521 3360
rect 42555 2584 42567 3360
rect 42509 2572 42567 2584
rect 42623 3360 42681 3372
rect 42623 2584 42635 3360
rect 42669 2584 42681 3360
rect 42623 2572 42681 2584
rect 42881 3360 42939 3372
rect 42881 2584 42893 3360
rect 42927 2584 42939 3360
rect 42881 2572 42939 2584
rect 42995 3360 43053 3372
rect 42995 2584 43007 3360
rect 43041 2584 43053 3360
rect 42995 2572 43053 2584
rect 43253 3360 43311 3372
rect 43253 2584 43265 3360
rect 43299 2584 43311 3360
rect 43253 2572 43311 2584
rect 43367 3360 43425 3372
rect 43367 2584 43379 3360
rect 43413 2584 43425 3360
rect 43367 2572 43425 2584
rect 43625 3360 43683 3372
rect 43625 2584 43637 3360
rect 43671 2584 43683 3360
rect 43625 2572 43683 2584
<< ndiffc >>
rect 40775 19336 40809 19512
rect 41033 19336 41067 19512
rect 41147 19336 41181 19512
rect 41405 19336 41439 19512
rect 41519 19336 41553 19512
rect 41777 19336 41811 19512
rect 41891 19336 41925 19512
rect 42149 19336 42183 19512
rect 42263 19336 42297 19512
rect 42521 19336 42555 19512
rect 42635 19336 42669 19512
rect 42893 19336 42927 19512
rect 43007 19336 43041 19512
rect 43265 19336 43299 19512
rect 43379 19336 43413 19512
rect 43637 19336 43671 19512
rect 43751 19336 43785 19512
rect 44009 19336 44043 19512
rect 44123 19336 44157 19512
rect 44381 19336 44415 19512
rect 44495 19336 44529 19512
rect 44753 19336 44787 19512
rect 44867 19336 44901 19512
rect 45125 19336 45159 19512
rect 45239 19336 45273 19512
rect 45497 19336 45531 19512
rect 45611 19336 45645 19512
rect 45869 19336 45903 19512
rect 45983 19336 46017 19512
rect 46241 19336 46275 19512
rect 46355 19336 46389 19512
rect 46613 19336 46647 19512
rect 46727 19336 46761 19512
rect 46985 19336 47019 19512
rect 47099 19336 47133 19512
rect 47357 19336 47391 19512
rect 47471 19336 47505 19512
rect 47729 19336 47763 19512
rect 47843 19336 47877 19512
rect 48101 19336 48135 19512
rect 48215 19336 48249 19512
rect 48473 19336 48507 19512
rect 48587 19336 48621 19512
rect 48845 19336 48879 19512
rect 48959 19336 48993 19512
rect 49217 19336 49251 19512
rect 49331 19336 49365 19512
rect 49589 19336 49623 19512
rect 40775 18918 40809 19094
rect 41033 18918 41067 19094
rect 41147 18918 41181 19094
rect 41405 18918 41439 19094
rect 41519 18918 41553 19094
rect 41777 18918 41811 19094
rect 41891 18918 41925 19094
rect 42149 18918 42183 19094
rect 42263 18918 42297 19094
rect 42521 18918 42555 19094
rect 42635 18918 42669 19094
rect 42893 18918 42927 19094
rect 43007 18918 43041 19094
rect 43265 18918 43299 19094
rect 43379 18918 43413 19094
rect 43637 18918 43671 19094
rect 43751 18918 43785 19094
rect 44009 18918 44043 19094
rect 44123 18918 44157 19094
rect 44381 18918 44415 19094
rect 44495 18918 44529 19094
rect 44753 18918 44787 19094
rect 44867 18918 44901 19094
rect 45125 18918 45159 19094
rect 45239 18918 45273 19094
rect 45497 18918 45531 19094
rect 45611 18918 45645 19094
rect 45869 18918 45903 19094
rect 45983 18918 46017 19094
rect 46241 18918 46275 19094
rect 46355 18918 46389 19094
rect 46613 18918 46647 19094
rect 46727 18918 46761 19094
rect 46985 18918 47019 19094
rect 47099 18918 47133 19094
rect 47357 18918 47391 19094
rect 47471 18918 47505 19094
rect 47729 18918 47763 19094
rect 47843 18918 47877 19094
rect 48101 18918 48135 19094
rect 48215 18918 48249 19094
rect 48473 18918 48507 19094
rect 48587 18918 48621 19094
rect 48845 18918 48879 19094
rect 48959 18918 48993 19094
rect 49217 18918 49251 19094
rect 49331 18918 49365 19094
rect 49589 18918 49623 19094
rect 40775 18500 40809 18676
rect 41033 18500 41067 18676
rect 41147 18500 41181 18676
rect 41405 18500 41439 18676
rect 41519 18500 41553 18676
rect 41777 18500 41811 18676
rect 41891 18500 41925 18676
rect 42149 18500 42183 18676
rect 42263 18500 42297 18676
rect 42521 18500 42555 18676
rect 42635 18500 42669 18676
rect 42893 18500 42927 18676
rect 43007 18500 43041 18676
rect 43265 18500 43299 18676
rect 43379 18500 43413 18676
rect 43637 18500 43671 18676
rect 43751 18500 43785 18676
rect 44009 18500 44043 18676
rect 44123 18500 44157 18676
rect 44381 18500 44415 18676
rect 44495 18500 44529 18676
rect 44753 18500 44787 18676
rect 44867 18500 44901 18676
rect 45125 18500 45159 18676
rect 45239 18500 45273 18676
rect 45497 18500 45531 18676
rect 45611 18500 45645 18676
rect 45869 18500 45903 18676
rect 45983 18500 46017 18676
rect 46241 18500 46275 18676
rect 46355 18500 46389 18676
rect 46613 18500 46647 18676
rect 46727 18500 46761 18676
rect 46985 18500 47019 18676
rect 47099 18500 47133 18676
rect 47357 18500 47391 18676
rect 47471 18500 47505 18676
rect 47729 18500 47763 18676
rect 47843 18500 47877 18676
rect 48101 18500 48135 18676
rect 48215 18500 48249 18676
rect 48473 18500 48507 18676
rect 48587 18500 48621 18676
rect 48845 18500 48879 18676
rect 48959 18500 48993 18676
rect 49217 18500 49251 18676
rect 49331 18500 49365 18676
rect 49589 18500 49623 18676
rect 40775 18082 40809 18258
rect 41033 18082 41067 18258
rect 41147 18082 41181 18258
rect 41405 18082 41439 18258
rect 41519 18082 41553 18258
rect 41777 18082 41811 18258
rect 41891 18082 41925 18258
rect 42149 18082 42183 18258
rect 42263 18082 42297 18258
rect 42521 18082 42555 18258
rect 42635 18082 42669 18258
rect 42893 18082 42927 18258
rect 43007 18082 43041 18258
rect 43265 18082 43299 18258
rect 43379 18082 43413 18258
rect 43637 18082 43671 18258
rect 43751 18082 43785 18258
rect 44009 18082 44043 18258
rect 44123 18082 44157 18258
rect 44381 18082 44415 18258
rect 44495 18082 44529 18258
rect 44753 18082 44787 18258
rect 44867 18082 44901 18258
rect 45125 18082 45159 18258
rect 45239 18082 45273 18258
rect 45497 18082 45531 18258
rect 45611 18082 45645 18258
rect 45869 18082 45903 18258
rect 45983 18082 46017 18258
rect 46241 18082 46275 18258
rect 46355 18082 46389 18258
rect 46613 18082 46647 18258
rect 46727 18082 46761 18258
rect 46985 18082 47019 18258
rect 47099 18082 47133 18258
rect 47357 18082 47391 18258
rect 47471 18082 47505 18258
rect 47729 18082 47763 18258
rect 47843 18082 47877 18258
rect 48101 18082 48135 18258
rect 48215 18082 48249 18258
rect 48473 18082 48507 18258
rect 48587 18082 48621 18258
rect 48845 18082 48879 18258
rect 48959 18082 48993 18258
rect 49217 18082 49251 18258
rect 49331 18082 49365 18258
rect 49589 18082 49623 18258
rect 40775 1607 40809 1783
rect 41033 1607 41067 1783
rect 41147 1607 41181 1783
rect 41405 1607 41439 1783
rect 41519 1607 41553 1783
rect 41777 1607 41811 1783
rect 41891 1607 41925 1783
rect 42149 1607 42183 1783
rect 42263 1607 42297 1783
rect 42521 1607 42555 1783
rect 42635 1607 42669 1783
rect 42893 1607 42927 1783
rect 43007 1607 43041 1783
rect 43265 1607 43299 1783
rect 43379 1607 43413 1783
rect 43637 1607 43671 1783
rect 43751 1607 43785 1783
rect 44009 1607 44043 1783
rect 44123 1607 44157 1783
rect 44381 1607 44415 1783
rect 44495 1607 44529 1783
rect 44753 1607 44787 1783
rect 44867 1607 44901 1783
rect 45125 1607 45159 1783
rect 45239 1607 45273 1783
rect 45497 1607 45531 1783
rect 45611 1607 45645 1783
rect 45869 1607 45903 1783
rect 45983 1607 46017 1783
rect 46241 1607 46275 1783
rect 46355 1607 46389 1783
rect 46613 1607 46647 1783
rect 46727 1607 46761 1783
rect 46985 1607 47019 1783
rect 47099 1607 47133 1783
rect 47357 1607 47391 1783
rect 47471 1607 47505 1783
rect 47729 1607 47763 1783
rect 47843 1607 47877 1783
rect 48101 1607 48135 1783
rect 48215 1607 48249 1783
rect 48473 1607 48507 1783
rect 48587 1607 48621 1783
rect 48845 1607 48879 1783
rect 48959 1607 48993 1783
rect 49217 1607 49251 1783
rect 49331 1607 49365 1783
rect 49589 1607 49623 1783
rect 40775 1189 40809 1365
rect 41033 1189 41067 1365
rect 41147 1189 41181 1365
rect 41405 1189 41439 1365
rect 41519 1189 41553 1365
rect 41777 1189 41811 1365
rect 41891 1189 41925 1365
rect 42149 1189 42183 1365
rect 42263 1189 42297 1365
rect 42521 1189 42555 1365
rect 42635 1189 42669 1365
rect 42893 1189 42927 1365
rect 43007 1189 43041 1365
rect 43265 1189 43299 1365
rect 43379 1189 43413 1365
rect 43637 1189 43671 1365
rect 43751 1189 43785 1365
rect 44009 1189 44043 1365
rect 44123 1189 44157 1365
rect 44381 1189 44415 1365
rect 44495 1189 44529 1365
rect 44753 1189 44787 1365
rect 44867 1189 44901 1365
rect 45125 1189 45159 1365
rect 45239 1189 45273 1365
rect 45497 1189 45531 1365
rect 45611 1189 45645 1365
rect 45869 1189 45903 1365
rect 45983 1189 46017 1365
rect 46241 1189 46275 1365
rect 46355 1189 46389 1365
rect 46613 1189 46647 1365
rect 46727 1189 46761 1365
rect 46985 1189 47019 1365
rect 47099 1189 47133 1365
rect 47357 1189 47391 1365
rect 47471 1189 47505 1365
rect 47729 1189 47763 1365
rect 47843 1189 47877 1365
rect 48101 1189 48135 1365
rect 48215 1189 48249 1365
rect 48473 1189 48507 1365
rect 48587 1189 48621 1365
rect 48845 1189 48879 1365
rect 48959 1189 48993 1365
rect 49217 1189 49251 1365
rect 49331 1189 49365 1365
rect 49589 1189 49623 1365
rect 40775 771 40809 947
rect 41033 771 41067 947
rect 41147 771 41181 947
rect 41405 771 41439 947
rect 41519 771 41553 947
rect 41777 771 41811 947
rect 41891 771 41925 947
rect 42149 771 42183 947
rect 42263 771 42297 947
rect 42521 771 42555 947
rect 42635 771 42669 947
rect 42893 771 42927 947
rect 43007 771 43041 947
rect 43265 771 43299 947
rect 43379 771 43413 947
rect 43637 771 43671 947
rect 43751 771 43785 947
rect 44009 771 44043 947
rect 44123 771 44157 947
rect 44381 771 44415 947
rect 44495 771 44529 947
rect 44753 771 44787 947
rect 44867 771 44901 947
rect 45125 771 45159 947
rect 45239 771 45273 947
rect 45497 771 45531 947
rect 45611 771 45645 947
rect 45869 771 45903 947
rect 45983 771 46017 947
rect 46241 771 46275 947
rect 46355 771 46389 947
rect 46613 771 46647 947
rect 46727 771 46761 947
rect 46985 771 47019 947
rect 47099 771 47133 947
rect 47357 771 47391 947
rect 47471 771 47505 947
rect 47729 771 47763 947
rect 47843 771 47877 947
rect 48101 771 48135 947
rect 48215 771 48249 947
rect 48473 771 48507 947
rect 48587 771 48621 947
rect 48845 771 48879 947
rect 48959 771 48993 947
rect 49217 771 49251 947
rect 49331 771 49365 947
rect 49589 771 49623 947
rect 40775 353 40809 529
rect 41033 353 41067 529
rect 41147 353 41181 529
rect 41405 353 41439 529
rect 41519 353 41553 529
rect 41777 353 41811 529
rect 41891 353 41925 529
rect 42149 353 42183 529
rect 42263 353 42297 529
rect 42521 353 42555 529
rect 42635 353 42669 529
rect 42893 353 42927 529
rect 43007 353 43041 529
rect 43265 353 43299 529
rect 43379 353 43413 529
rect 43637 353 43671 529
rect 43751 353 43785 529
rect 44009 353 44043 529
rect 44123 353 44157 529
rect 44381 353 44415 529
rect 44495 353 44529 529
rect 44753 353 44787 529
rect 44867 353 44901 529
rect 45125 353 45159 529
rect 45239 353 45273 529
rect 45497 353 45531 529
rect 45611 353 45645 529
rect 45869 353 45903 529
rect 45983 353 46017 529
rect 46241 353 46275 529
rect 46355 353 46389 529
rect 46613 353 46647 529
rect 46727 353 46761 529
rect 46985 353 47019 529
rect 47099 353 47133 529
rect 47357 353 47391 529
rect 47471 353 47505 529
rect 47729 353 47763 529
rect 47843 353 47877 529
rect 48101 353 48135 529
rect 48215 353 48249 529
rect 48473 353 48507 529
rect 48587 353 48621 529
rect 48845 353 48879 529
rect 48959 353 48993 529
rect 49217 353 49251 529
rect 49331 353 49365 529
rect 49589 353 49623 529
<< pdiffc >>
rect 40775 16505 40809 17281
rect 41033 16505 41067 17281
rect 41147 16505 41181 17281
rect 41405 16505 41439 17281
rect 41519 16505 41553 17281
rect 41777 16505 41811 17281
rect 41891 16505 41925 17281
rect 42149 16505 42183 17281
rect 42263 16505 42297 17281
rect 42521 16505 42555 17281
rect 42635 16505 42669 17281
rect 42893 16505 42927 17281
rect 43007 16505 43041 17281
rect 43265 16505 43299 17281
rect 43379 16505 43413 17281
rect 43637 16505 43671 17281
rect 40775 15469 40809 16245
rect 41033 15469 41067 16245
rect 41147 15469 41181 16245
rect 41405 15469 41439 16245
rect 41519 15469 41553 16245
rect 41777 15469 41811 16245
rect 41891 15469 41925 16245
rect 42149 15469 42183 16245
rect 42263 15469 42297 16245
rect 42521 15469 42555 16245
rect 42635 15469 42669 16245
rect 42893 15469 42927 16245
rect 43007 15469 43041 16245
rect 43265 15469 43299 16245
rect 43379 15469 43413 16245
rect 43637 15469 43671 16245
rect 40775 14433 40809 15209
rect 41033 14433 41067 15209
rect 41147 14433 41181 15209
rect 41405 14433 41439 15209
rect 41519 14433 41553 15209
rect 41777 14433 41811 15209
rect 41891 14433 41925 15209
rect 42149 14433 42183 15209
rect 42263 14433 42297 15209
rect 42521 14433 42555 15209
rect 42635 14433 42669 15209
rect 42893 14433 42927 15209
rect 43007 14433 43041 15209
rect 43265 14433 43299 15209
rect 43379 14433 43413 15209
rect 43637 14433 43671 15209
rect 40775 13397 40809 14173
rect 41033 13397 41067 14173
rect 41147 13397 41181 14173
rect 41405 13397 41439 14173
rect 41519 13397 41553 14173
rect 41777 13397 41811 14173
rect 41891 13397 41925 14173
rect 42149 13397 42183 14173
rect 42263 13397 42297 14173
rect 42521 13397 42555 14173
rect 42635 13397 42669 14173
rect 42893 13397 42927 14173
rect 43007 13397 43041 14173
rect 43265 13397 43299 14173
rect 43379 13397 43413 14173
rect 43637 13397 43671 14173
rect 39287 12281 39321 12657
rect 39545 12281 39579 12657
rect 39659 12281 39693 12657
rect 39917 12281 39951 12657
rect 40031 12281 40065 12657
rect 40289 12281 40323 12657
rect 40403 12281 40437 12657
rect 40661 12281 40695 12657
rect 40775 12281 40809 12657
rect 41033 12281 41067 12657
rect 41147 12281 41181 12657
rect 41405 12281 41439 12657
rect 41519 12281 41553 12657
rect 41777 12281 41811 12657
rect 41891 12281 41925 12657
rect 42149 12281 42183 12657
rect 42263 12281 42297 12657
rect 42521 12281 42555 12657
rect 42635 12281 42669 12657
rect 42893 12281 42927 12657
rect 43007 12281 43041 12657
rect 43265 12281 43299 12657
rect 43379 12281 43413 12657
rect 43637 12281 43671 12657
rect 43751 12281 43785 12657
rect 44009 12281 44043 12657
rect 44123 12281 44157 12657
rect 44381 12281 44415 12657
rect 44495 12281 44529 12657
rect 44753 12281 44787 12657
rect 44867 12281 44901 12657
rect 45125 12281 45159 12657
rect 45239 12281 45273 12657
rect 45497 12281 45531 12657
rect 45611 12281 45645 12657
rect 45869 12281 45903 12657
rect 45983 12281 46017 12657
rect 46241 12281 46275 12657
rect 46355 12281 46389 12657
rect 46613 12281 46647 12657
rect 46727 12281 46761 12657
rect 46985 12281 47019 12657
rect 47099 12281 47133 12657
rect 47357 12281 47391 12657
rect 47471 12281 47505 12657
rect 47729 12281 47763 12657
rect 47843 12281 47877 12657
rect 48101 12281 48135 12657
rect 48215 12281 48249 12657
rect 48473 12281 48507 12657
rect 48587 12281 48621 12657
rect 48845 12281 48879 12657
rect 48959 12281 48993 12657
rect 49217 12281 49251 12657
rect 49331 12281 49365 12657
rect 49589 12281 49623 12657
rect 49703 12281 49737 12657
rect 49961 12281 49995 12657
rect 50075 12281 50109 12657
rect 50333 12281 50367 12657
rect 50447 12281 50481 12657
rect 50705 12281 50739 12657
rect 50819 12281 50853 12657
rect 51077 12281 51111 12657
rect 39287 11645 39321 12021
rect 39545 11645 39579 12021
rect 39659 11645 39693 12021
rect 39917 11645 39951 12021
rect 40031 11645 40065 12021
rect 40289 11645 40323 12021
rect 40403 11645 40437 12021
rect 40661 11645 40695 12021
rect 40775 11645 40809 12021
rect 41033 11645 41067 12021
rect 41147 11645 41181 12021
rect 41405 11645 41439 12021
rect 41519 11645 41553 12021
rect 41777 11645 41811 12021
rect 41891 11645 41925 12021
rect 42149 11645 42183 12021
rect 42263 11645 42297 12021
rect 42521 11645 42555 12021
rect 42635 11645 42669 12021
rect 42893 11645 42927 12021
rect 43007 11645 43041 12021
rect 43265 11645 43299 12021
rect 43379 11645 43413 12021
rect 43637 11645 43671 12021
rect 43751 11645 43785 12021
rect 44009 11645 44043 12021
rect 44123 11645 44157 12021
rect 44381 11645 44415 12021
rect 44495 11645 44529 12021
rect 44753 11645 44787 12021
rect 44867 11645 44901 12021
rect 45125 11645 45159 12021
rect 45239 11645 45273 12021
rect 45497 11645 45531 12021
rect 45611 11645 45645 12021
rect 45869 11645 45903 12021
rect 45983 11645 46017 12021
rect 46241 11645 46275 12021
rect 46355 11645 46389 12021
rect 46613 11645 46647 12021
rect 46727 11645 46761 12021
rect 46985 11645 47019 12021
rect 47099 11645 47133 12021
rect 47357 11645 47391 12021
rect 47471 11645 47505 12021
rect 47729 11645 47763 12021
rect 47843 11645 47877 12021
rect 48101 11645 48135 12021
rect 48215 11645 48249 12021
rect 48473 11645 48507 12021
rect 48587 11645 48621 12021
rect 48845 11645 48879 12021
rect 48959 11645 48993 12021
rect 49217 11645 49251 12021
rect 49331 11645 49365 12021
rect 49589 11645 49623 12021
rect 49703 11645 49737 12021
rect 49961 11645 49995 12021
rect 50075 11645 50109 12021
rect 50333 11645 50367 12021
rect 50447 11645 50481 12021
rect 50705 11645 50739 12021
rect 50819 11645 50853 12021
rect 51077 11645 51111 12021
rect 39287 11009 39321 11385
rect 39545 11009 39579 11385
rect 39659 11009 39693 11385
rect 39917 11009 39951 11385
rect 40031 11009 40065 11385
rect 40289 11009 40323 11385
rect 40403 11009 40437 11385
rect 40661 11009 40695 11385
rect 40775 11009 40809 11385
rect 41033 11009 41067 11385
rect 41147 11009 41181 11385
rect 41405 11009 41439 11385
rect 41519 11009 41553 11385
rect 41777 11009 41811 11385
rect 41891 11009 41925 11385
rect 42149 11009 42183 11385
rect 42263 11009 42297 11385
rect 42521 11009 42555 11385
rect 42635 11009 42669 11385
rect 42893 11009 42927 11385
rect 43007 11009 43041 11385
rect 43265 11009 43299 11385
rect 43379 11009 43413 11385
rect 43637 11009 43671 11385
rect 43751 11009 43785 11385
rect 44009 11009 44043 11385
rect 44123 11009 44157 11385
rect 44381 11009 44415 11385
rect 44495 11009 44529 11385
rect 44753 11009 44787 11385
rect 44867 11009 44901 11385
rect 45125 11009 45159 11385
rect 45239 11009 45273 11385
rect 45497 11009 45531 11385
rect 45611 11009 45645 11385
rect 45869 11009 45903 11385
rect 45983 11009 46017 11385
rect 46241 11009 46275 11385
rect 46355 11009 46389 11385
rect 46613 11009 46647 11385
rect 46727 11009 46761 11385
rect 46985 11009 47019 11385
rect 47099 11009 47133 11385
rect 47357 11009 47391 11385
rect 47471 11009 47505 11385
rect 47729 11009 47763 11385
rect 47843 11009 47877 11385
rect 48101 11009 48135 11385
rect 48215 11009 48249 11385
rect 48473 11009 48507 11385
rect 48587 11009 48621 11385
rect 48845 11009 48879 11385
rect 48959 11009 48993 11385
rect 49217 11009 49251 11385
rect 49331 11009 49365 11385
rect 49589 11009 49623 11385
rect 49703 11009 49737 11385
rect 49961 11009 49995 11385
rect 50075 11009 50109 11385
rect 50333 11009 50367 11385
rect 50447 11009 50481 11385
rect 50705 11009 50739 11385
rect 50819 11009 50853 11385
rect 51077 11009 51111 11385
rect 39287 8480 39321 8856
rect 39545 8480 39579 8856
rect 39659 8480 39693 8856
rect 39917 8480 39951 8856
rect 40031 8480 40065 8856
rect 40289 8480 40323 8856
rect 40403 8480 40437 8856
rect 40661 8480 40695 8856
rect 40775 8480 40809 8856
rect 41033 8480 41067 8856
rect 41147 8480 41181 8856
rect 41405 8480 41439 8856
rect 41519 8480 41553 8856
rect 41777 8480 41811 8856
rect 41891 8480 41925 8856
rect 42149 8480 42183 8856
rect 42263 8480 42297 8856
rect 42521 8480 42555 8856
rect 42635 8480 42669 8856
rect 42893 8480 42927 8856
rect 43007 8480 43041 8856
rect 43265 8480 43299 8856
rect 43379 8480 43413 8856
rect 43637 8480 43671 8856
rect 43751 8480 43785 8856
rect 44009 8480 44043 8856
rect 44123 8480 44157 8856
rect 44381 8480 44415 8856
rect 44495 8480 44529 8856
rect 44753 8480 44787 8856
rect 44867 8480 44901 8856
rect 45125 8480 45159 8856
rect 45239 8480 45273 8856
rect 45497 8480 45531 8856
rect 45611 8480 45645 8856
rect 45869 8480 45903 8856
rect 45983 8480 46017 8856
rect 46241 8480 46275 8856
rect 46355 8480 46389 8856
rect 46613 8480 46647 8856
rect 46727 8480 46761 8856
rect 46985 8480 47019 8856
rect 47099 8480 47133 8856
rect 47357 8480 47391 8856
rect 47471 8480 47505 8856
rect 47729 8480 47763 8856
rect 47843 8480 47877 8856
rect 48101 8480 48135 8856
rect 48215 8480 48249 8856
rect 48473 8480 48507 8856
rect 48587 8480 48621 8856
rect 48845 8480 48879 8856
rect 48959 8480 48993 8856
rect 49217 8480 49251 8856
rect 49331 8480 49365 8856
rect 49589 8480 49623 8856
rect 49703 8480 49737 8856
rect 49961 8480 49995 8856
rect 50075 8480 50109 8856
rect 50333 8480 50367 8856
rect 50447 8480 50481 8856
rect 50705 8480 50739 8856
rect 50819 8480 50853 8856
rect 51077 8480 51111 8856
rect 39287 7844 39321 8220
rect 39545 7844 39579 8220
rect 39659 7844 39693 8220
rect 39917 7844 39951 8220
rect 40031 7844 40065 8220
rect 40289 7844 40323 8220
rect 40403 7844 40437 8220
rect 40661 7844 40695 8220
rect 40775 7844 40809 8220
rect 41033 7844 41067 8220
rect 41147 7844 41181 8220
rect 41405 7844 41439 8220
rect 41519 7844 41553 8220
rect 41777 7844 41811 8220
rect 41891 7844 41925 8220
rect 42149 7844 42183 8220
rect 42263 7844 42297 8220
rect 42521 7844 42555 8220
rect 42635 7844 42669 8220
rect 42893 7844 42927 8220
rect 43007 7844 43041 8220
rect 43265 7844 43299 8220
rect 43379 7844 43413 8220
rect 43637 7844 43671 8220
rect 43751 7844 43785 8220
rect 44009 7844 44043 8220
rect 44123 7844 44157 8220
rect 44381 7844 44415 8220
rect 44495 7844 44529 8220
rect 44753 7844 44787 8220
rect 44867 7844 44901 8220
rect 45125 7844 45159 8220
rect 45239 7844 45273 8220
rect 45497 7844 45531 8220
rect 45611 7844 45645 8220
rect 45869 7844 45903 8220
rect 45983 7844 46017 8220
rect 46241 7844 46275 8220
rect 46355 7844 46389 8220
rect 46613 7844 46647 8220
rect 46727 7844 46761 8220
rect 46985 7844 47019 8220
rect 47099 7844 47133 8220
rect 47357 7844 47391 8220
rect 47471 7844 47505 8220
rect 47729 7844 47763 8220
rect 47843 7844 47877 8220
rect 48101 7844 48135 8220
rect 48215 7844 48249 8220
rect 48473 7844 48507 8220
rect 48587 7844 48621 8220
rect 48845 7844 48879 8220
rect 48959 7844 48993 8220
rect 49217 7844 49251 8220
rect 49331 7844 49365 8220
rect 49589 7844 49623 8220
rect 49703 7844 49737 8220
rect 49961 7844 49995 8220
rect 50075 7844 50109 8220
rect 50333 7844 50367 8220
rect 50447 7844 50481 8220
rect 50705 7844 50739 8220
rect 50819 7844 50853 8220
rect 51077 7844 51111 8220
rect 39287 7208 39321 7584
rect 39545 7208 39579 7584
rect 39659 7208 39693 7584
rect 39917 7208 39951 7584
rect 40031 7208 40065 7584
rect 40289 7208 40323 7584
rect 40403 7208 40437 7584
rect 40661 7208 40695 7584
rect 40775 7208 40809 7584
rect 41033 7208 41067 7584
rect 41147 7208 41181 7584
rect 41405 7208 41439 7584
rect 41519 7208 41553 7584
rect 41777 7208 41811 7584
rect 41891 7208 41925 7584
rect 42149 7208 42183 7584
rect 42263 7208 42297 7584
rect 42521 7208 42555 7584
rect 42635 7208 42669 7584
rect 42893 7208 42927 7584
rect 43007 7208 43041 7584
rect 43265 7208 43299 7584
rect 43379 7208 43413 7584
rect 43637 7208 43671 7584
rect 43751 7208 43785 7584
rect 44009 7208 44043 7584
rect 44123 7208 44157 7584
rect 44381 7208 44415 7584
rect 44495 7208 44529 7584
rect 44753 7208 44787 7584
rect 44867 7208 44901 7584
rect 45125 7208 45159 7584
rect 45239 7208 45273 7584
rect 45497 7208 45531 7584
rect 45611 7208 45645 7584
rect 45869 7208 45903 7584
rect 45983 7208 46017 7584
rect 46241 7208 46275 7584
rect 46355 7208 46389 7584
rect 46613 7208 46647 7584
rect 46727 7208 46761 7584
rect 46985 7208 47019 7584
rect 47099 7208 47133 7584
rect 47357 7208 47391 7584
rect 47471 7208 47505 7584
rect 47729 7208 47763 7584
rect 47843 7208 47877 7584
rect 48101 7208 48135 7584
rect 48215 7208 48249 7584
rect 48473 7208 48507 7584
rect 48587 7208 48621 7584
rect 48845 7208 48879 7584
rect 48959 7208 48993 7584
rect 49217 7208 49251 7584
rect 49331 7208 49365 7584
rect 49589 7208 49623 7584
rect 49703 7208 49737 7584
rect 49961 7208 49995 7584
rect 50075 7208 50109 7584
rect 50333 7208 50367 7584
rect 50447 7208 50481 7584
rect 50705 7208 50739 7584
rect 50819 7208 50853 7584
rect 51077 7208 51111 7584
rect 40775 5692 40809 6468
rect 41033 5692 41067 6468
rect 41147 5692 41181 6468
rect 41405 5692 41439 6468
rect 41519 5692 41553 6468
rect 41777 5692 41811 6468
rect 41891 5692 41925 6468
rect 42149 5692 42183 6468
rect 42263 5692 42297 6468
rect 42521 5692 42555 6468
rect 42635 5692 42669 6468
rect 42893 5692 42927 6468
rect 43007 5692 43041 6468
rect 43265 5692 43299 6468
rect 43379 5692 43413 6468
rect 43637 5692 43671 6468
rect 40775 4656 40809 5432
rect 41033 4656 41067 5432
rect 41147 4656 41181 5432
rect 41405 4656 41439 5432
rect 41519 4656 41553 5432
rect 41777 4656 41811 5432
rect 41891 4656 41925 5432
rect 42149 4656 42183 5432
rect 42263 4656 42297 5432
rect 42521 4656 42555 5432
rect 42635 4656 42669 5432
rect 42893 4656 42927 5432
rect 43007 4656 43041 5432
rect 43265 4656 43299 5432
rect 43379 4656 43413 5432
rect 43637 4656 43671 5432
rect 40775 3620 40809 4396
rect 41033 3620 41067 4396
rect 41147 3620 41181 4396
rect 41405 3620 41439 4396
rect 41519 3620 41553 4396
rect 41777 3620 41811 4396
rect 41891 3620 41925 4396
rect 42149 3620 42183 4396
rect 42263 3620 42297 4396
rect 42521 3620 42555 4396
rect 42635 3620 42669 4396
rect 42893 3620 42927 4396
rect 43007 3620 43041 4396
rect 43265 3620 43299 4396
rect 43379 3620 43413 4396
rect 43637 3620 43671 4396
rect 40775 2584 40809 3360
rect 41033 2584 41067 3360
rect 41147 2584 41181 3360
rect 41405 2584 41439 3360
rect 41519 2584 41553 3360
rect 41777 2584 41811 3360
rect 41891 2584 41925 3360
rect 42149 2584 42183 3360
rect 42263 2584 42297 3360
rect 42521 2584 42555 3360
rect 42635 2584 42669 3360
rect 42893 2584 42927 3360
rect 43007 2584 43041 3360
rect 43265 2584 43299 3360
rect 43379 2584 43413 3360
rect 43637 2584 43671 3360
<< psubdiff >>
rect 40661 19664 40757 19698
rect 49641 19664 49737 19698
rect 40661 19602 40695 19664
rect 49703 19602 49737 19664
rect 40661 17930 40695 17992
rect 49703 17930 49737 17992
rect 40661 17896 40757 17930
rect 49641 17896 49737 17930
rect 45825 16548 45921 16582
rect 46059 16548 46155 16582
rect 45825 16486 45859 16548
rect 46121 16486 46155 16548
rect 45825 15392 45859 15454
rect 46121 15392 46155 15454
rect 45825 15358 45921 15392
rect 46059 15358 46155 15392
rect 39375 6836 39471 6870
rect 39927 6836 40023 6870
rect 39375 6774 39409 6836
rect 39989 6774 40023 6836
rect 39375 4780 39409 4842
rect 39989 4780 40023 4842
rect 39375 4746 39471 4780
rect 39927 4746 40023 4780
rect 44531 6196 44627 6230
rect 45083 6196 45179 6230
rect 44531 6134 44565 6196
rect 45145 6134 45179 6196
rect 44531 4140 44565 4202
rect 45145 4140 45179 4202
rect 44531 4106 44627 4140
rect 45083 4106 45179 4140
rect 45825 4473 45921 4507
rect 46059 4473 46155 4507
rect 45825 4411 45859 4473
rect 46121 4411 46155 4473
rect 45825 3317 45859 3379
rect 46121 3317 46155 3379
rect 45825 3283 45921 3317
rect 46059 3283 46155 3317
rect 40661 1935 40757 1969
rect 49641 1935 49737 1969
rect 40661 1873 40695 1935
rect 49703 1873 49737 1935
rect 40661 201 40695 263
rect 49703 201 49737 263
rect 40661 167 40757 201
rect 49641 167 49737 201
<< nsubdiff >>
rect 40661 17442 40757 17476
rect 43689 17442 43785 17476
rect 40661 17380 40695 17442
rect 43751 17380 43785 17442
rect 40661 13236 40695 13298
rect 43751 13236 43785 13298
rect 40661 13202 40757 13236
rect 43689 13202 43785 13236
rect 39173 12818 39269 12852
rect 51129 12818 51225 12852
rect 39173 12756 39207 12818
rect 51191 12756 51225 12818
rect 39173 10848 39207 10910
rect 51191 10848 51225 10910
rect 39173 10814 39269 10848
rect 51129 10814 51225 10848
rect 39173 9017 39269 9051
rect 51129 9017 51225 9051
rect 39173 8955 39207 9017
rect 51191 8955 51225 9017
rect 39173 7047 39207 7109
rect 51191 7047 51225 7109
rect 39173 7013 39269 7047
rect 51129 7013 51225 7047
rect 40661 6629 40757 6663
rect 43689 6629 43785 6663
rect 40661 6567 40695 6629
rect 43751 6567 43785 6629
rect 40661 2423 40695 2485
rect 43751 2423 43785 2485
rect 40661 2389 40757 2423
rect 43689 2389 43785 2423
<< psubdiffcont >>
rect 40757 19664 49641 19698
rect 40661 17992 40695 19602
rect 49703 17992 49737 19602
rect 40757 17896 49641 17930
rect 45921 16548 46059 16582
rect 45825 15454 45859 16486
rect 46121 15454 46155 16486
rect 45921 15358 46059 15392
rect 39471 6836 39927 6870
rect 39375 4842 39409 6774
rect 39989 4842 40023 6774
rect 39471 4746 39927 4780
rect 44627 6196 45083 6230
rect 44531 4202 44565 6134
rect 45145 4202 45179 6134
rect 44627 4106 45083 4140
rect 45921 4473 46059 4507
rect 45825 3379 45859 4411
rect 46121 3379 46155 4411
rect 45921 3283 46059 3317
rect 40757 1935 49641 1969
rect 40661 263 40695 1873
rect 49703 263 49737 1873
rect 40757 167 49641 201
<< nsubdiffcont >>
rect 40757 17442 43689 17476
rect 40661 13298 40695 17380
rect 43751 13298 43785 17380
rect 40757 13202 43689 13236
rect 39269 12818 51129 12852
rect 39173 10910 39207 12756
rect 51191 10910 51225 12756
rect 39269 10814 51129 10848
rect 39269 9017 51129 9051
rect 39173 7109 39207 8955
rect 51191 7109 51225 8955
rect 39269 7013 51129 7047
rect 40757 6629 43689 6663
rect 40661 2485 40695 6567
rect 43751 2485 43785 6567
rect 40757 2389 43689 2423
<< poly >>
rect 40821 19596 41021 19612
rect 40821 19562 40837 19596
rect 41005 19562 41021 19596
rect 40821 19524 41021 19562
rect 41193 19596 41393 19612
rect 41193 19562 41209 19596
rect 41377 19562 41393 19596
rect 41193 19524 41393 19562
rect 41565 19596 41765 19612
rect 41565 19562 41581 19596
rect 41749 19562 41765 19596
rect 41565 19524 41765 19562
rect 41937 19596 42137 19612
rect 41937 19562 41953 19596
rect 42121 19562 42137 19596
rect 41937 19524 42137 19562
rect 42309 19596 42509 19612
rect 42309 19562 42325 19596
rect 42493 19562 42509 19596
rect 42309 19524 42509 19562
rect 42681 19596 42881 19612
rect 42681 19562 42697 19596
rect 42865 19562 42881 19596
rect 42681 19524 42881 19562
rect 43053 19596 43253 19612
rect 43053 19562 43069 19596
rect 43237 19562 43253 19596
rect 43053 19524 43253 19562
rect 43425 19596 43625 19612
rect 43425 19562 43441 19596
rect 43609 19562 43625 19596
rect 43425 19524 43625 19562
rect 43797 19596 43997 19612
rect 43797 19562 43813 19596
rect 43981 19562 43997 19596
rect 43797 19524 43997 19562
rect 44169 19596 44369 19612
rect 44169 19562 44185 19596
rect 44353 19562 44369 19596
rect 44169 19524 44369 19562
rect 44541 19596 44741 19612
rect 44541 19562 44557 19596
rect 44725 19562 44741 19596
rect 44541 19524 44741 19562
rect 44913 19596 45113 19612
rect 44913 19562 44929 19596
rect 45097 19562 45113 19596
rect 44913 19524 45113 19562
rect 45285 19596 45485 19612
rect 45285 19562 45301 19596
rect 45469 19562 45485 19596
rect 45285 19524 45485 19562
rect 45657 19596 45857 19612
rect 45657 19562 45673 19596
rect 45841 19562 45857 19596
rect 45657 19524 45857 19562
rect 46029 19596 46229 19612
rect 46029 19562 46045 19596
rect 46213 19562 46229 19596
rect 46029 19524 46229 19562
rect 46401 19596 46601 19612
rect 46401 19562 46417 19596
rect 46585 19562 46601 19596
rect 46401 19524 46601 19562
rect 46773 19596 46973 19612
rect 46773 19562 46789 19596
rect 46957 19562 46973 19596
rect 46773 19524 46973 19562
rect 47145 19596 47345 19612
rect 47145 19562 47161 19596
rect 47329 19562 47345 19596
rect 47145 19524 47345 19562
rect 47517 19596 47717 19612
rect 47517 19562 47533 19596
rect 47701 19562 47717 19596
rect 47517 19524 47717 19562
rect 47889 19596 48089 19612
rect 47889 19562 47905 19596
rect 48073 19562 48089 19596
rect 47889 19524 48089 19562
rect 48261 19596 48461 19612
rect 48261 19562 48277 19596
rect 48445 19562 48461 19596
rect 48261 19524 48461 19562
rect 48633 19596 48833 19612
rect 48633 19562 48649 19596
rect 48817 19562 48833 19596
rect 48633 19524 48833 19562
rect 49005 19596 49205 19612
rect 49005 19562 49021 19596
rect 49189 19562 49205 19596
rect 49005 19524 49205 19562
rect 49377 19596 49577 19612
rect 49377 19562 49393 19596
rect 49561 19562 49577 19596
rect 49377 19524 49577 19562
rect 40821 19286 41021 19324
rect 40821 19252 40837 19286
rect 41005 19252 41021 19286
rect 40821 19236 41021 19252
rect 41193 19286 41393 19324
rect 41193 19252 41209 19286
rect 41377 19252 41393 19286
rect 41193 19236 41393 19252
rect 41565 19286 41765 19324
rect 41565 19252 41581 19286
rect 41749 19252 41765 19286
rect 41565 19236 41765 19252
rect 41937 19286 42137 19324
rect 41937 19252 41953 19286
rect 42121 19252 42137 19286
rect 41937 19236 42137 19252
rect 42309 19286 42509 19324
rect 42309 19252 42325 19286
rect 42493 19252 42509 19286
rect 42309 19236 42509 19252
rect 42681 19286 42881 19324
rect 42681 19252 42697 19286
rect 42865 19252 42881 19286
rect 42681 19236 42881 19252
rect 43053 19286 43253 19324
rect 43053 19252 43069 19286
rect 43237 19252 43253 19286
rect 43053 19236 43253 19252
rect 43425 19286 43625 19324
rect 43425 19252 43441 19286
rect 43609 19252 43625 19286
rect 43425 19236 43625 19252
rect 43797 19286 43997 19324
rect 43797 19252 43813 19286
rect 43981 19252 43997 19286
rect 43797 19236 43997 19252
rect 44169 19286 44369 19324
rect 44169 19252 44185 19286
rect 44353 19252 44369 19286
rect 44169 19236 44369 19252
rect 44541 19286 44741 19324
rect 44541 19252 44557 19286
rect 44725 19252 44741 19286
rect 44541 19236 44741 19252
rect 44913 19286 45113 19324
rect 44913 19252 44929 19286
rect 45097 19252 45113 19286
rect 44913 19236 45113 19252
rect 45285 19286 45485 19324
rect 45285 19252 45301 19286
rect 45469 19252 45485 19286
rect 45285 19236 45485 19252
rect 45657 19286 45857 19324
rect 45657 19252 45673 19286
rect 45841 19252 45857 19286
rect 45657 19236 45857 19252
rect 46029 19286 46229 19324
rect 46029 19252 46045 19286
rect 46213 19252 46229 19286
rect 46029 19236 46229 19252
rect 46401 19286 46601 19324
rect 46401 19252 46417 19286
rect 46585 19252 46601 19286
rect 46401 19236 46601 19252
rect 46773 19286 46973 19324
rect 46773 19252 46789 19286
rect 46957 19252 46973 19286
rect 46773 19236 46973 19252
rect 47145 19286 47345 19324
rect 47145 19252 47161 19286
rect 47329 19252 47345 19286
rect 47145 19236 47345 19252
rect 47517 19286 47717 19324
rect 47517 19252 47533 19286
rect 47701 19252 47717 19286
rect 47517 19236 47717 19252
rect 47889 19286 48089 19324
rect 47889 19252 47905 19286
rect 48073 19252 48089 19286
rect 47889 19236 48089 19252
rect 48261 19286 48461 19324
rect 48261 19252 48277 19286
rect 48445 19252 48461 19286
rect 48261 19236 48461 19252
rect 48633 19286 48833 19324
rect 48633 19252 48649 19286
rect 48817 19252 48833 19286
rect 48633 19236 48833 19252
rect 49005 19286 49205 19324
rect 49005 19252 49021 19286
rect 49189 19252 49205 19286
rect 49005 19236 49205 19252
rect 49377 19286 49577 19324
rect 49377 19252 49393 19286
rect 49561 19252 49577 19286
rect 49377 19236 49577 19252
rect 40821 19178 41021 19194
rect 40821 19144 40837 19178
rect 41005 19144 41021 19178
rect 40821 19106 41021 19144
rect 41193 19178 41393 19194
rect 41193 19144 41209 19178
rect 41377 19144 41393 19178
rect 41193 19106 41393 19144
rect 41565 19178 41765 19194
rect 41565 19144 41581 19178
rect 41749 19144 41765 19178
rect 41565 19106 41765 19144
rect 41937 19178 42137 19194
rect 41937 19144 41953 19178
rect 42121 19144 42137 19178
rect 41937 19106 42137 19144
rect 42309 19178 42509 19194
rect 42309 19144 42325 19178
rect 42493 19144 42509 19178
rect 42309 19106 42509 19144
rect 42681 19178 42881 19194
rect 42681 19144 42697 19178
rect 42865 19144 42881 19178
rect 42681 19106 42881 19144
rect 43053 19178 43253 19194
rect 43053 19144 43069 19178
rect 43237 19144 43253 19178
rect 43053 19106 43253 19144
rect 43425 19178 43625 19194
rect 43425 19144 43441 19178
rect 43609 19144 43625 19178
rect 43425 19106 43625 19144
rect 43797 19178 43997 19194
rect 43797 19144 43813 19178
rect 43981 19144 43997 19178
rect 43797 19106 43997 19144
rect 44169 19178 44369 19194
rect 44169 19144 44185 19178
rect 44353 19144 44369 19178
rect 44169 19106 44369 19144
rect 44541 19178 44741 19194
rect 44541 19144 44557 19178
rect 44725 19144 44741 19178
rect 44541 19106 44741 19144
rect 44913 19178 45113 19194
rect 44913 19144 44929 19178
rect 45097 19144 45113 19178
rect 44913 19106 45113 19144
rect 45285 19178 45485 19194
rect 45285 19144 45301 19178
rect 45469 19144 45485 19178
rect 45285 19106 45485 19144
rect 45657 19178 45857 19194
rect 45657 19144 45673 19178
rect 45841 19144 45857 19178
rect 45657 19106 45857 19144
rect 46029 19178 46229 19194
rect 46029 19144 46045 19178
rect 46213 19144 46229 19178
rect 46029 19106 46229 19144
rect 46401 19178 46601 19194
rect 46401 19144 46417 19178
rect 46585 19144 46601 19178
rect 46401 19106 46601 19144
rect 46773 19178 46973 19194
rect 46773 19144 46789 19178
rect 46957 19144 46973 19178
rect 46773 19106 46973 19144
rect 47145 19178 47345 19194
rect 47145 19144 47161 19178
rect 47329 19144 47345 19178
rect 47145 19106 47345 19144
rect 47517 19178 47717 19194
rect 47517 19144 47533 19178
rect 47701 19144 47717 19178
rect 47517 19106 47717 19144
rect 47889 19178 48089 19194
rect 47889 19144 47905 19178
rect 48073 19144 48089 19178
rect 47889 19106 48089 19144
rect 48261 19178 48461 19194
rect 48261 19144 48277 19178
rect 48445 19144 48461 19178
rect 48261 19106 48461 19144
rect 48633 19178 48833 19194
rect 48633 19144 48649 19178
rect 48817 19144 48833 19178
rect 48633 19106 48833 19144
rect 49005 19178 49205 19194
rect 49005 19144 49021 19178
rect 49189 19144 49205 19178
rect 49005 19106 49205 19144
rect 49377 19178 49577 19194
rect 49377 19144 49393 19178
rect 49561 19144 49577 19178
rect 49377 19106 49577 19144
rect 40821 18868 41021 18906
rect 40821 18834 40837 18868
rect 41005 18834 41021 18868
rect 40821 18818 41021 18834
rect 41193 18868 41393 18906
rect 41193 18834 41209 18868
rect 41377 18834 41393 18868
rect 41193 18818 41393 18834
rect 41565 18868 41765 18906
rect 41565 18834 41581 18868
rect 41749 18834 41765 18868
rect 41565 18818 41765 18834
rect 41937 18868 42137 18906
rect 41937 18834 41953 18868
rect 42121 18834 42137 18868
rect 41937 18818 42137 18834
rect 42309 18868 42509 18906
rect 42309 18834 42325 18868
rect 42493 18834 42509 18868
rect 42309 18818 42509 18834
rect 42681 18868 42881 18906
rect 42681 18834 42697 18868
rect 42865 18834 42881 18868
rect 42681 18818 42881 18834
rect 43053 18868 43253 18906
rect 43053 18834 43069 18868
rect 43237 18834 43253 18868
rect 43053 18818 43253 18834
rect 43425 18868 43625 18906
rect 43425 18834 43441 18868
rect 43609 18834 43625 18868
rect 43425 18818 43625 18834
rect 43797 18868 43997 18906
rect 43797 18834 43813 18868
rect 43981 18834 43997 18868
rect 43797 18818 43997 18834
rect 44169 18868 44369 18906
rect 44169 18834 44185 18868
rect 44353 18834 44369 18868
rect 44169 18818 44369 18834
rect 44541 18868 44741 18906
rect 44541 18834 44557 18868
rect 44725 18834 44741 18868
rect 44541 18818 44741 18834
rect 44913 18868 45113 18906
rect 44913 18834 44929 18868
rect 45097 18834 45113 18868
rect 44913 18818 45113 18834
rect 45285 18868 45485 18906
rect 45285 18834 45301 18868
rect 45469 18834 45485 18868
rect 45285 18818 45485 18834
rect 45657 18868 45857 18906
rect 45657 18834 45673 18868
rect 45841 18834 45857 18868
rect 45657 18818 45857 18834
rect 46029 18868 46229 18906
rect 46029 18834 46045 18868
rect 46213 18834 46229 18868
rect 46029 18818 46229 18834
rect 46401 18868 46601 18906
rect 46401 18834 46417 18868
rect 46585 18834 46601 18868
rect 46401 18818 46601 18834
rect 46773 18868 46973 18906
rect 46773 18834 46789 18868
rect 46957 18834 46973 18868
rect 46773 18818 46973 18834
rect 47145 18868 47345 18906
rect 47145 18834 47161 18868
rect 47329 18834 47345 18868
rect 47145 18818 47345 18834
rect 47517 18868 47717 18906
rect 47517 18834 47533 18868
rect 47701 18834 47717 18868
rect 47517 18818 47717 18834
rect 47889 18868 48089 18906
rect 47889 18834 47905 18868
rect 48073 18834 48089 18868
rect 47889 18818 48089 18834
rect 48261 18868 48461 18906
rect 48261 18834 48277 18868
rect 48445 18834 48461 18868
rect 48261 18818 48461 18834
rect 48633 18868 48833 18906
rect 48633 18834 48649 18868
rect 48817 18834 48833 18868
rect 48633 18818 48833 18834
rect 49005 18868 49205 18906
rect 49005 18834 49021 18868
rect 49189 18834 49205 18868
rect 49005 18818 49205 18834
rect 49377 18868 49577 18906
rect 49377 18834 49393 18868
rect 49561 18834 49577 18868
rect 49377 18818 49577 18834
rect 40821 18760 41021 18776
rect 40821 18726 40837 18760
rect 41005 18726 41021 18760
rect 40821 18688 41021 18726
rect 41193 18760 41393 18776
rect 41193 18726 41209 18760
rect 41377 18726 41393 18760
rect 41193 18688 41393 18726
rect 41565 18760 41765 18776
rect 41565 18726 41581 18760
rect 41749 18726 41765 18760
rect 41565 18688 41765 18726
rect 41937 18760 42137 18776
rect 41937 18726 41953 18760
rect 42121 18726 42137 18760
rect 41937 18688 42137 18726
rect 42309 18760 42509 18776
rect 42309 18726 42325 18760
rect 42493 18726 42509 18760
rect 42309 18688 42509 18726
rect 42681 18760 42881 18776
rect 42681 18726 42697 18760
rect 42865 18726 42881 18760
rect 42681 18688 42881 18726
rect 43053 18760 43253 18776
rect 43053 18726 43069 18760
rect 43237 18726 43253 18760
rect 43053 18688 43253 18726
rect 43425 18760 43625 18776
rect 43425 18726 43441 18760
rect 43609 18726 43625 18760
rect 43425 18688 43625 18726
rect 43797 18760 43997 18776
rect 43797 18726 43813 18760
rect 43981 18726 43997 18760
rect 43797 18688 43997 18726
rect 44169 18760 44369 18776
rect 44169 18726 44185 18760
rect 44353 18726 44369 18760
rect 44169 18688 44369 18726
rect 44541 18760 44741 18776
rect 44541 18726 44557 18760
rect 44725 18726 44741 18760
rect 44541 18688 44741 18726
rect 44913 18760 45113 18776
rect 44913 18726 44929 18760
rect 45097 18726 45113 18760
rect 44913 18688 45113 18726
rect 45285 18760 45485 18776
rect 45285 18726 45301 18760
rect 45469 18726 45485 18760
rect 45285 18688 45485 18726
rect 45657 18760 45857 18776
rect 45657 18726 45673 18760
rect 45841 18726 45857 18760
rect 45657 18688 45857 18726
rect 46029 18760 46229 18776
rect 46029 18726 46045 18760
rect 46213 18726 46229 18760
rect 46029 18688 46229 18726
rect 46401 18760 46601 18776
rect 46401 18726 46417 18760
rect 46585 18726 46601 18760
rect 46401 18688 46601 18726
rect 46773 18760 46973 18776
rect 46773 18726 46789 18760
rect 46957 18726 46973 18760
rect 46773 18688 46973 18726
rect 47145 18760 47345 18776
rect 47145 18726 47161 18760
rect 47329 18726 47345 18760
rect 47145 18688 47345 18726
rect 47517 18760 47717 18776
rect 47517 18726 47533 18760
rect 47701 18726 47717 18760
rect 47517 18688 47717 18726
rect 47889 18760 48089 18776
rect 47889 18726 47905 18760
rect 48073 18726 48089 18760
rect 47889 18688 48089 18726
rect 48261 18760 48461 18776
rect 48261 18726 48277 18760
rect 48445 18726 48461 18760
rect 48261 18688 48461 18726
rect 48633 18760 48833 18776
rect 48633 18726 48649 18760
rect 48817 18726 48833 18760
rect 48633 18688 48833 18726
rect 49005 18760 49205 18776
rect 49005 18726 49021 18760
rect 49189 18726 49205 18760
rect 49005 18688 49205 18726
rect 49377 18760 49577 18776
rect 49377 18726 49393 18760
rect 49561 18726 49577 18760
rect 49377 18688 49577 18726
rect 40821 18450 41021 18488
rect 40821 18416 40837 18450
rect 41005 18416 41021 18450
rect 40821 18400 41021 18416
rect 41193 18450 41393 18488
rect 41193 18416 41209 18450
rect 41377 18416 41393 18450
rect 41193 18400 41393 18416
rect 41565 18450 41765 18488
rect 41565 18416 41581 18450
rect 41749 18416 41765 18450
rect 41565 18400 41765 18416
rect 41937 18450 42137 18488
rect 41937 18416 41953 18450
rect 42121 18416 42137 18450
rect 41937 18400 42137 18416
rect 42309 18450 42509 18488
rect 42309 18416 42325 18450
rect 42493 18416 42509 18450
rect 42309 18400 42509 18416
rect 42681 18450 42881 18488
rect 42681 18416 42697 18450
rect 42865 18416 42881 18450
rect 42681 18400 42881 18416
rect 43053 18450 43253 18488
rect 43053 18416 43069 18450
rect 43237 18416 43253 18450
rect 43053 18400 43253 18416
rect 43425 18450 43625 18488
rect 43425 18416 43441 18450
rect 43609 18416 43625 18450
rect 43425 18400 43625 18416
rect 43797 18450 43997 18488
rect 43797 18416 43813 18450
rect 43981 18416 43997 18450
rect 43797 18400 43997 18416
rect 44169 18450 44369 18488
rect 44169 18416 44185 18450
rect 44353 18416 44369 18450
rect 44169 18400 44369 18416
rect 44541 18450 44741 18488
rect 44541 18416 44557 18450
rect 44725 18416 44741 18450
rect 44541 18400 44741 18416
rect 44913 18450 45113 18488
rect 44913 18416 44929 18450
rect 45097 18416 45113 18450
rect 44913 18400 45113 18416
rect 45285 18450 45485 18488
rect 45285 18416 45301 18450
rect 45469 18416 45485 18450
rect 45285 18400 45485 18416
rect 45657 18450 45857 18488
rect 45657 18416 45673 18450
rect 45841 18416 45857 18450
rect 45657 18400 45857 18416
rect 46029 18450 46229 18488
rect 46029 18416 46045 18450
rect 46213 18416 46229 18450
rect 46029 18400 46229 18416
rect 46401 18450 46601 18488
rect 46401 18416 46417 18450
rect 46585 18416 46601 18450
rect 46401 18400 46601 18416
rect 46773 18450 46973 18488
rect 46773 18416 46789 18450
rect 46957 18416 46973 18450
rect 46773 18400 46973 18416
rect 47145 18450 47345 18488
rect 47145 18416 47161 18450
rect 47329 18416 47345 18450
rect 47145 18400 47345 18416
rect 47517 18450 47717 18488
rect 47517 18416 47533 18450
rect 47701 18416 47717 18450
rect 47517 18400 47717 18416
rect 47889 18450 48089 18488
rect 47889 18416 47905 18450
rect 48073 18416 48089 18450
rect 47889 18400 48089 18416
rect 48261 18450 48461 18488
rect 48261 18416 48277 18450
rect 48445 18416 48461 18450
rect 48261 18400 48461 18416
rect 48633 18450 48833 18488
rect 48633 18416 48649 18450
rect 48817 18416 48833 18450
rect 48633 18400 48833 18416
rect 49005 18450 49205 18488
rect 49005 18416 49021 18450
rect 49189 18416 49205 18450
rect 49005 18400 49205 18416
rect 49377 18450 49577 18488
rect 49377 18416 49393 18450
rect 49561 18416 49577 18450
rect 49377 18400 49577 18416
rect 40821 18342 41021 18358
rect 40821 18308 40837 18342
rect 41005 18308 41021 18342
rect 40821 18270 41021 18308
rect 41193 18342 41393 18358
rect 41193 18308 41209 18342
rect 41377 18308 41393 18342
rect 41193 18270 41393 18308
rect 41565 18342 41765 18358
rect 41565 18308 41581 18342
rect 41749 18308 41765 18342
rect 41565 18270 41765 18308
rect 41937 18342 42137 18358
rect 41937 18308 41953 18342
rect 42121 18308 42137 18342
rect 41937 18270 42137 18308
rect 42309 18342 42509 18358
rect 42309 18308 42325 18342
rect 42493 18308 42509 18342
rect 42309 18270 42509 18308
rect 42681 18342 42881 18358
rect 42681 18308 42697 18342
rect 42865 18308 42881 18342
rect 42681 18270 42881 18308
rect 43053 18342 43253 18358
rect 43053 18308 43069 18342
rect 43237 18308 43253 18342
rect 43053 18270 43253 18308
rect 43425 18342 43625 18358
rect 43425 18308 43441 18342
rect 43609 18308 43625 18342
rect 43425 18270 43625 18308
rect 43797 18342 43997 18358
rect 43797 18308 43813 18342
rect 43981 18308 43997 18342
rect 43797 18270 43997 18308
rect 44169 18342 44369 18358
rect 44169 18308 44185 18342
rect 44353 18308 44369 18342
rect 44169 18270 44369 18308
rect 44541 18342 44741 18358
rect 44541 18308 44557 18342
rect 44725 18308 44741 18342
rect 44541 18270 44741 18308
rect 44913 18342 45113 18358
rect 44913 18308 44929 18342
rect 45097 18308 45113 18342
rect 44913 18270 45113 18308
rect 45285 18342 45485 18358
rect 45285 18308 45301 18342
rect 45469 18308 45485 18342
rect 45285 18270 45485 18308
rect 45657 18342 45857 18358
rect 45657 18308 45673 18342
rect 45841 18308 45857 18342
rect 45657 18270 45857 18308
rect 46029 18342 46229 18358
rect 46029 18308 46045 18342
rect 46213 18308 46229 18342
rect 46029 18270 46229 18308
rect 46401 18342 46601 18358
rect 46401 18308 46417 18342
rect 46585 18308 46601 18342
rect 46401 18270 46601 18308
rect 46773 18342 46973 18358
rect 46773 18308 46789 18342
rect 46957 18308 46973 18342
rect 46773 18270 46973 18308
rect 47145 18342 47345 18358
rect 47145 18308 47161 18342
rect 47329 18308 47345 18342
rect 47145 18270 47345 18308
rect 47517 18342 47717 18358
rect 47517 18308 47533 18342
rect 47701 18308 47717 18342
rect 47517 18270 47717 18308
rect 47889 18342 48089 18358
rect 47889 18308 47905 18342
rect 48073 18308 48089 18342
rect 47889 18270 48089 18308
rect 48261 18342 48461 18358
rect 48261 18308 48277 18342
rect 48445 18308 48461 18342
rect 48261 18270 48461 18308
rect 48633 18342 48833 18358
rect 48633 18308 48649 18342
rect 48817 18308 48833 18342
rect 48633 18270 48833 18308
rect 49005 18342 49205 18358
rect 49005 18308 49021 18342
rect 49189 18308 49205 18342
rect 49005 18270 49205 18308
rect 49377 18342 49577 18358
rect 49377 18308 49393 18342
rect 49561 18308 49577 18342
rect 49377 18270 49577 18308
rect 40821 18032 41021 18070
rect 40821 17998 40837 18032
rect 41005 17998 41021 18032
rect 40821 17982 41021 17998
rect 41193 18032 41393 18070
rect 41193 17998 41209 18032
rect 41377 17998 41393 18032
rect 41193 17982 41393 17998
rect 41565 18032 41765 18070
rect 41565 17998 41581 18032
rect 41749 17998 41765 18032
rect 41565 17982 41765 17998
rect 41937 18032 42137 18070
rect 41937 17998 41953 18032
rect 42121 17998 42137 18032
rect 41937 17982 42137 17998
rect 42309 18032 42509 18070
rect 42309 17998 42325 18032
rect 42493 17998 42509 18032
rect 42309 17982 42509 17998
rect 42681 18032 42881 18070
rect 42681 17998 42697 18032
rect 42865 17998 42881 18032
rect 42681 17982 42881 17998
rect 43053 18032 43253 18070
rect 43053 17998 43069 18032
rect 43237 17998 43253 18032
rect 43053 17982 43253 17998
rect 43425 18032 43625 18070
rect 43425 17998 43441 18032
rect 43609 17998 43625 18032
rect 43425 17982 43625 17998
rect 43797 18032 43997 18070
rect 43797 17998 43813 18032
rect 43981 17998 43997 18032
rect 43797 17982 43997 17998
rect 44169 18032 44369 18070
rect 44169 17998 44185 18032
rect 44353 17998 44369 18032
rect 44169 17982 44369 17998
rect 44541 18032 44741 18070
rect 44541 17998 44557 18032
rect 44725 17998 44741 18032
rect 44541 17982 44741 17998
rect 44913 18032 45113 18070
rect 44913 17998 44929 18032
rect 45097 17998 45113 18032
rect 44913 17982 45113 17998
rect 45285 18032 45485 18070
rect 45285 17998 45301 18032
rect 45469 17998 45485 18032
rect 45285 17982 45485 17998
rect 45657 18032 45857 18070
rect 45657 17998 45673 18032
rect 45841 17998 45857 18032
rect 45657 17982 45857 17998
rect 46029 18032 46229 18070
rect 46029 17998 46045 18032
rect 46213 17998 46229 18032
rect 46029 17982 46229 17998
rect 46401 18032 46601 18070
rect 46401 17998 46417 18032
rect 46585 17998 46601 18032
rect 46401 17982 46601 17998
rect 46773 18032 46973 18070
rect 46773 17998 46789 18032
rect 46957 17998 46973 18032
rect 46773 17982 46973 17998
rect 47145 18032 47345 18070
rect 47145 17998 47161 18032
rect 47329 17998 47345 18032
rect 47145 17982 47345 17998
rect 47517 18032 47717 18070
rect 47517 17998 47533 18032
rect 47701 17998 47717 18032
rect 47517 17982 47717 17998
rect 47889 18032 48089 18070
rect 47889 17998 47905 18032
rect 48073 17998 48089 18032
rect 47889 17982 48089 17998
rect 48261 18032 48461 18070
rect 48261 17998 48277 18032
rect 48445 17998 48461 18032
rect 48261 17982 48461 17998
rect 48633 18032 48833 18070
rect 48633 17998 48649 18032
rect 48817 17998 48833 18032
rect 48633 17982 48833 17998
rect 49005 18032 49205 18070
rect 49005 17998 49021 18032
rect 49189 17998 49205 18032
rect 49005 17982 49205 17998
rect 49377 18032 49577 18070
rect 49377 17998 49393 18032
rect 49561 17998 49577 18032
rect 49377 17982 49577 17998
rect 40821 17374 41021 17390
rect 40821 17340 40837 17374
rect 41005 17340 41021 17374
rect 40821 17293 41021 17340
rect 41193 17374 41393 17390
rect 41193 17340 41209 17374
rect 41377 17340 41393 17374
rect 41193 17293 41393 17340
rect 41565 17374 41765 17390
rect 41565 17340 41581 17374
rect 41749 17340 41765 17374
rect 41565 17293 41765 17340
rect 41937 17374 42137 17390
rect 41937 17340 41953 17374
rect 42121 17340 42137 17374
rect 41937 17293 42137 17340
rect 42309 17374 42509 17390
rect 42309 17340 42325 17374
rect 42493 17340 42509 17374
rect 42309 17293 42509 17340
rect 42681 17374 42881 17390
rect 42681 17340 42697 17374
rect 42865 17340 42881 17374
rect 42681 17293 42881 17340
rect 43053 17374 43253 17390
rect 43053 17340 43069 17374
rect 43237 17340 43253 17374
rect 43053 17293 43253 17340
rect 43425 17374 43625 17390
rect 43425 17340 43441 17374
rect 43609 17340 43625 17374
rect 43425 17293 43625 17340
rect 40821 16446 41021 16493
rect 40821 16412 40837 16446
rect 41005 16412 41021 16446
rect 40821 16396 41021 16412
rect 41193 16446 41393 16493
rect 41193 16412 41209 16446
rect 41377 16412 41393 16446
rect 41193 16396 41393 16412
rect 41565 16446 41765 16493
rect 41565 16412 41581 16446
rect 41749 16412 41765 16446
rect 41565 16396 41765 16412
rect 41937 16446 42137 16493
rect 41937 16412 41953 16446
rect 42121 16412 42137 16446
rect 41937 16396 42137 16412
rect 42309 16446 42509 16493
rect 42309 16412 42325 16446
rect 42493 16412 42509 16446
rect 42309 16396 42509 16412
rect 42681 16446 42881 16493
rect 42681 16412 42697 16446
rect 42865 16412 42881 16446
rect 42681 16396 42881 16412
rect 43053 16446 43253 16493
rect 43053 16412 43069 16446
rect 43237 16412 43253 16446
rect 43053 16396 43253 16412
rect 43425 16446 43625 16493
rect 43425 16412 43441 16446
rect 43609 16412 43625 16446
rect 43425 16396 43625 16412
rect 40821 16338 41021 16354
rect 40821 16304 40837 16338
rect 41005 16304 41021 16338
rect 40821 16257 41021 16304
rect 41193 16338 41393 16354
rect 41193 16304 41209 16338
rect 41377 16304 41393 16338
rect 41193 16257 41393 16304
rect 41565 16338 41765 16354
rect 41565 16304 41581 16338
rect 41749 16304 41765 16338
rect 41565 16257 41765 16304
rect 41937 16338 42137 16354
rect 41937 16304 41953 16338
rect 42121 16304 42137 16338
rect 41937 16257 42137 16304
rect 42309 16338 42509 16354
rect 42309 16304 42325 16338
rect 42493 16304 42509 16338
rect 42309 16257 42509 16304
rect 42681 16338 42881 16354
rect 42681 16304 42697 16338
rect 42865 16304 42881 16338
rect 42681 16257 42881 16304
rect 43053 16338 43253 16354
rect 43053 16304 43069 16338
rect 43237 16304 43253 16338
rect 43053 16257 43253 16304
rect 43425 16338 43625 16354
rect 43425 16304 43441 16338
rect 43609 16304 43625 16338
rect 43425 16257 43625 16304
rect 40821 15410 41021 15457
rect 40821 15376 40837 15410
rect 41005 15376 41021 15410
rect 40821 15360 41021 15376
rect 41193 15410 41393 15457
rect 41193 15376 41209 15410
rect 41377 15376 41393 15410
rect 41193 15360 41393 15376
rect 41565 15410 41765 15457
rect 41565 15376 41581 15410
rect 41749 15376 41765 15410
rect 41565 15360 41765 15376
rect 41937 15410 42137 15457
rect 41937 15376 41953 15410
rect 42121 15376 42137 15410
rect 41937 15360 42137 15376
rect 42309 15410 42509 15457
rect 42309 15376 42325 15410
rect 42493 15376 42509 15410
rect 42309 15360 42509 15376
rect 42681 15410 42881 15457
rect 42681 15376 42697 15410
rect 42865 15376 42881 15410
rect 42681 15360 42881 15376
rect 43053 15410 43253 15457
rect 43053 15376 43069 15410
rect 43237 15376 43253 15410
rect 43053 15360 43253 15376
rect 43425 15410 43625 15457
rect 43425 15376 43441 15410
rect 43609 15376 43625 15410
rect 43425 15360 43625 15376
rect 40821 15302 41021 15318
rect 40821 15268 40837 15302
rect 41005 15268 41021 15302
rect 40821 15221 41021 15268
rect 41193 15302 41393 15318
rect 41193 15268 41209 15302
rect 41377 15268 41393 15302
rect 41193 15221 41393 15268
rect 41565 15302 41765 15318
rect 41565 15268 41581 15302
rect 41749 15268 41765 15302
rect 41565 15221 41765 15268
rect 41937 15302 42137 15318
rect 41937 15268 41953 15302
rect 42121 15268 42137 15302
rect 41937 15221 42137 15268
rect 42309 15302 42509 15318
rect 42309 15268 42325 15302
rect 42493 15268 42509 15302
rect 42309 15221 42509 15268
rect 42681 15302 42881 15318
rect 42681 15268 42697 15302
rect 42865 15268 42881 15302
rect 42681 15221 42881 15268
rect 43053 15302 43253 15318
rect 43053 15268 43069 15302
rect 43237 15268 43253 15302
rect 43053 15221 43253 15268
rect 43425 15302 43625 15318
rect 43425 15268 43441 15302
rect 43609 15268 43625 15302
rect 43425 15221 43625 15268
rect 40821 14374 41021 14421
rect 40821 14340 40837 14374
rect 41005 14340 41021 14374
rect 40821 14324 41021 14340
rect 41193 14374 41393 14421
rect 41193 14340 41209 14374
rect 41377 14340 41393 14374
rect 41193 14324 41393 14340
rect 41565 14374 41765 14421
rect 41565 14340 41581 14374
rect 41749 14340 41765 14374
rect 41565 14324 41765 14340
rect 41937 14374 42137 14421
rect 41937 14340 41953 14374
rect 42121 14340 42137 14374
rect 41937 14324 42137 14340
rect 42309 14374 42509 14421
rect 42309 14340 42325 14374
rect 42493 14340 42509 14374
rect 42309 14324 42509 14340
rect 42681 14374 42881 14421
rect 42681 14340 42697 14374
rect 42865 14340 42881 14374
rect 42681 14324 42881 14340
rect 43053 14374 43253 14421
rect 43053 14340 43069 14374
rect 43237 14340 43253 14374
rect 43053 14324 43253 14340
rect 43425 14374 43625 14421
rect 43425 14340 43441 14374
rect 43609 14340 43625 14374
rect 43425 14324 43625 14340
rect 40821 14266 41021 14282
rect 40821 14232 40837 14266
rect 41005 14232 41021 14266
rect 40821 14185 41021 14232
rect 41193 14266 41393 14282
rect 41193 14232 41209 14266
rect 41377 14232 41393 14266
rect 41193 14185 41393 14232
rect 41565 14266 41765 14282
rect 41565 14232 41581 14266
rect 41749 14232 41765 14266
rect 41565 14185 41765 14232
rect 41937 14266 42137 14282
rect 41937 14232 41953 14266
rect 42121 14232 42137 14266
rect 41937 14185 42137 14232
rect 42309 14266 42509 14282
rect 42309 14232 42325 14266
rect 42493 14232 42509 14266
rect 42309 14185 42509 14232
rect 42681 14266 42881 14282
rect 42681 14232 42697 14266
rect 42865 14232 42881 14266
rect 42681 14185 42881 14232
rect 43053 14266 43253 14282
rect 43053 14232 43069 14266
rect 43237 14232 43253 14266
rect 43053 14185 43253 14232
rect 43425 14266 43625 14282
rect 43425 14232 43441 14266
rect 43609 14232 43625 14266
rect 43425 14185 43625 14232
rect 40821 13338 41021 13385
rect 40821 13304 40837 13338
rect 41005 13304 41021 13338
rect 40821 13288 41021 13304
rect 41193 13338 41393 13385
rect 41193 13304 41209 13338
rect 41377 13304 41393 13338
rect 41193 13288 41393 13304
rect 41565 13338 41765 13385
rect 41565 13304 41581 13338
rect 41749 13304 41765 13338
rect 41565 13288 41765 13304
rect 41937 13338 42137 13385
rect 41937 13304 41953 13338
rect 42121 13304 42137 13338
rect 41937 13288 42137 13304
rect 42309 13338 42509 13385
rect 42309 13304 42325 13338
rect 42493 13304 42509 13338
rect 42309 13288 42509 13304
rect 42681 13338 42881 13385
rect 42681 13304 42697 13338
rect 42865 13304 42881 13338
rect 42681 13288 42881 13304
rect 43053 13338 43253 13385
rect 43053 13304 43069 13338
rect 43237 13304 43253 13338
rect 43053 13288 43253 13304
rect 43425 13338 43625 13385
rect 43425 13304 43441 13338
rect 43609 13304 43625 13338
rect 43425 13288 43625 13304
rect 39333 12750 39533 12766
rect 39333 12716 39349 12750
rect 39517 12716 39533 12750
rect 39333 12669 39533 12716
rect 39705 12750 39905 12766
rect 39705 12716 39721 12750
rect 39889 12716 39905 12750
rect 39705 12669 39905 12716
rect 40077 12750 40277 12766
rect 40077 12716 40093 12750
rect 40261 12716 40277 12750
rect 40077 12669 40277 12716
rect 40449 12750 40649 12766
rect 40449 12716 40465 12750
rect 40633 12716 40649 12750
rect 40449 12669 40649 12716
rect 40821 12750 41021 12766
rect 40821 12716 40837 12750
rect 41005 12716 41021 12750
rect 40821 12669 41021 12716
rect 41193 12750 41393 12766
rect 41193 12716 41209 12750
rect 41377 12716 41393 12750
rect 41193 12669 41393 12716
rect 41565 12750 41765 12766
rect 41565 12716 41581 12750
rect 41749 12716 41765 12750
rect 41565 12669 41765 12716
rect 41937 12750 42137 12766
rect 41937 12716 41953 12750
rect 42121 12716 42137 12750
rect 41937 12669 42137 12716
rect 42309 12750 42509 12766
rect 42309 12716 42325 12750
rect 42493 12716 42509 12750
rect 42309 12669 42509 12716
rect 42681 12750 42881 12766
rect 42681 12716 42697 12750
rect 42865 12716 42881 12750
rect 42681 12669 42881 12716
rect 43053 12750 43253 12766
rect 43053 12716 43069 12750
rect 43237 12716 43253 12750
rect 43053 12669 43253 12716
rect 43425 12750 43625 12766
rect 43425 12716 43441 12750
rect 43609 12716 43625 12750
rect 43425 12669 43625 12716
rect 43797 12750 43997 12766
rect 43797 12716 43813 12750
rect 43981 12716 43997 12750
rect 43797 12669 43997 12716
rect 44169 12750 44369 12766
rect 44169 12716 44185 12750
rect 44353 12716 44369 12750
rect 44169 12669 44369 12716
rect 44541 12750 44741 12766
rect 44541 12716 44557 12750
rect 44725 12716 44741 12750
rect 44541 12669 44741 12716
rect 44913 12750 45113 12766
rect 44913 12716 44929 12750
rect 45097 12716 45113 12750
rect 44913 12669 45113 12716
rect 45285 12750 45485 12766
rect 45285 12716 45301 12750
rect 45469 12716 45485 12750
rect 45285 12669 45485 12716
rect 45657 12750 45857 12766
rect 45657 12716 45673 12750
rect 45841 12716 45857 12750
rect 45657 12669 45857 12716
rect 46029 12750 46229 12766
rect 46029 12716 46045 12750
rect 46213 12716 46229 12750
rect 46029 12669 46229 12716
rect 46401 12750 46601 12766
rect 46401 12716 46417 12750
rect 46585 12716 46601 12750
rect 46401 12669 46601 12716
rect 46773 12750 46973 12766
rect 46773 12716 46789 12750
rect 46957 12716 46973 12750
rect 46773 12669 46973 12716
rect 47145 12750 47345 12766
rect 47145 12716 47161 12750
rect 47329 12716 47345 12750
rect 47145 12669 47345 12716
rect 47517 12750 47717 12766
rect 47517 12716 47533 12750
rect 47701 12716 47717 12750
rect 47517 12669 47717 12716
rect 47889 12750 48089 12766
rect 47889 12716 47905 12750
rect 48073 12716 48089 12750
rect 47889 12669 48089 12716
rect 48261 12750 48461 12766
rect 48261 12716 48277 12750
rect 48445 12716 48461 12750
rect 48261 12669 48461 12716
rect 48633 12750 48833 12766
rect 48633 12716 48649 12750
rect 48817 12716 48833 12750
rect 48633 12669 48833 12716
rect 49005 12750 49205 12766
rect 49005 12716 49021 12750
rect 49189 12716 49205 12750
rect 49005 12669 49205 12716
rect 49377 12750 49577 12766
rect 49377 12716 49393 12750
rect 49561 12716 49577 12750
rect 49377 12669 49577 12716
rect 49749 12750 49949 12766
rect 49749 12716 49765 12750
rect 49933 12716 49949 12750
rect 49749 12669 49949 12716
rect 50121 12750 50321 12766
rect 50121 12716 50137 12750
rect 50305 12716 50321 12750
rect 50121 12669 50321 12716
rect 50493 12750 50693 12766
rect 50493 12716 50509 12750
rect 50677 12716 50693 12750
rect 50493 12669 50693 12716
rect 50865 12750 51065 12766
rect 50865 12716 50881 12750
rect 51049 12716 51065 12750
rect 50865 12669 51065 12716
rect 39333 12222 39533 12269
rect 39333 12188 39349 12222
rect 39517 12188 39533 12222
rect 39333 12172 39533 12188
rect 39705 12222 39905 12269
rect 39705 12188 39721 12222
rect 39889 12188 39905 12222
rect 39705 12172 39905 12188
rect 40077 12222 40277 12269
rect 40077 12188 40093 12222
rect 40261 12188 40277 12222
rect 40077 12172 40277 12188
rect 40449 12222 40649 12269
rect 40449 12188 40465 12222
rect 40633 12188 40649 12222
rect 40449 12172 40649 12188
rect 40821 12222 41021 12269
rect 40821 12188 40837 12222
rect 41005 12188 41021 12222
rect 40821 12172 41021 12188
rect 41193 12222 41393 12269
rect 41193 12188 41209 12222
rect 41377 12188 41393 12222
rect 41193 12172 41393 12188
rect 41565 12222 41765 12269
rect 41565 12188 41581 12222
rect 41749 12188 41765 12222
rect 41565 12172 41765 12188
rect 41937 12222 42137 12269
rect 41937 12188 41953 12222
rect 42121 12188 42137 12222
rect 41937 12172 42137 12188
rect 42309 12222 42509 12269
rect 42309 12188 42325 12222
rect 42493 12188 42509 12222
rect 42309 12172 42509 12188
rect 42681 12222 42881 12269
rect 42681 12188 42697 12222
rect 42865 12188 42881 12222
rect 42681 12172 42881 12188
rect 43053 12222 43253 12269
rect 43053 12188 43069 12222
rect 43237 12188 43253 12222
rect 43053 12172 43253 12188
rect 43425 12222 43625 12269
rect 43425 12188 43441 12222
rect 43609 12188 43625 12222
rect 43425 12172 43625 12188
rect 43797 12222 43997 12269
rect 43797 12188 43813 12222
rect 43981 12188 43997 12222
rect 43797 12172 43997 12188
rect 44169 12222 44369 12269
rect 44169 12188 44185 12222
rect 44353 12188 44369 12222
rect 44169 12172 44369 12188
rect 44541 12222 44741 12269
rect 44541 12188 44557 12222
rect 44725 12188 44741 12222
rect 44541 12172 44741 12188
rect 44913 12222 45113 12269
rect 44913 12188 44929 12222
rect 45097 12188 45113 12222
rect 44913 12172 45113 12188
rect 45285 12222 45485 12269
rect 45285 12188 45301 12222
rect 45469 12188 45485 12222
rect 45285 12172 45485 12188
rect 45657 12222 45857 12269
rect 45657 12188 45673 12222
rect 45841 12188 45857 12222
rect 45657 12172 45857 12188
rect 46029 12222 46229 12269
rect 46029 12188 46045 12222
rect 46213 12188 46229 12222
rect 46029 12172 46229 12188
rect 46401 12222 46601 12269
rect 46401 12188 46417 12222
rect 46585 12188 46601 12222
rect 46401 12172 46601 12188
rect 46773 12222 46973 12269
rect 46773 12188 46789 12222
rect 46957 12188 46973 12222
rect 46773 12172 46973 12188
rect 47145 12222 47345 12269
rect 47145 12188 47161 12222
rect 47329 12188 47345 12222
rect 47145 12172 47345 12188
rect 47517 12222 47717 12269
rect 47517 12188 47533 12222
rect 47701 12188 47717 12222
rect 47517 12172 47717 12188
rect 47889 12222 48089 12269
rect 47889 12188 47905 12222
rect 48073 12188 48089 12222
rect 47889 12172 48089 12188
rect 48261 12222 48461 12269
rect 48261 12188 48277 12222
rect 48445 12188 48461 12222
rect 48261 12172 48461 12188
rect 48633 12222 48833 12269
rect 48633 12188 48649 12222
rect 48817 12188 48833 12222
rect 48633 12172 48833 12188
rect 49005 12222 49205 12269
rect 49005 12188 49021 12222
rect 49189 12188 49205 12222
rect 49005 12172 49205 12188
rect 49377 12222 49577 12269
rect 49377 12188 49393 12222
rect 49561 12188 49577 12222
rect 49377 12172 49577 12188
rect 49749 12222 49949 12269
rect 49749 12188 49765 12222
rect 49933 12188 49949 12222
rect 49749 12172 49949 12188
rect 50121 12222 50321 12269
rect 50121 12188 50137 12222
rect 50305 12188 50321 12222
rect 50121 12172 50321 12188
rect 50493 12222 50693 12269
rect 50493 12188 50509 12222
rect 50677 12188 50693 12222
rect 50493 12172 50693 12188
rect 50865 12222 51065 12269
rect 50865 12188 50881 12222
rect 51049 12188 51065 12222
rect 50865 12172 51065 12188
rect 39333 12114 39533 12130
rect 39333 12080 39349 12114
rect 39517 12080 39533 12114
rect 39333 12033 39533 12080
rect 39705 12114 39905 12130
rect 39705 12080 39721 12114
rect 39889 12080 39905 12114
rect 39705 12033 39905 12080
rect 40077 12114 40277 12130
rect 40077 12080 40093 12114
rect 40261 12080 40277 12114
rect 40077 12033 40277 12080
rect 40449 12114 40649 12130
rect 40449 12080 40465 12114
rect 40633 12080 40649 12114
rect 40449 12033 40649 12080
rect 40821 12114 41021 12130
rect 40821 12080 40837 12114
rect 41005 12080 41021 12114
rect 40821 12033 41021 12080
rect 41193 12114 41393 12130
rect 41193 12080 41209 12114
rect 41377 12080 41393 12114
rect 41193 12033 41393 12080
rect 41565 12114 41765 12130
rect 41565 12080 41581 12114
rect 41749 12080 41765 12114
rect 41565 12033 41765 12080
rect 41937 12114 42137 12130
rect 41937 12080 41953 12114
rect 42121 12080 42137 12114
rect 41937 12033 42137 12080
rect 42309 12114 42509 12130
rect 42309 12080 42325 12114
rect 42493 12080 42509 12114
rect 42309 12033 42509 12080
rect 42681 12114 42881 12130
rect 42681 12080 42697 12114
rect 42865 12080 42881 12114
rect 42681 12033 42881 12080
rect 43053 12114 43253 12130
rect 43053 12080 43069 12114
rect 43237 12080 43253 12114
rect 43053 12033 43253 12080
rect 43425 12114 43625 12130
rect 43425 12080 43441 12114
rect 43609 12080 43625 12114
rect 43425 12033 43625 12080
rect 43797 12114 43997 12130
rect 43797 12080 43813 12114
rect 43981 12080 43997 12114
rect 43797 12033 43997 12080
rect 44169 12114 44369 12130
rect 44169 12080 44185 12114
rect 44353 12080 44369 12114
rect 44169 12033 44369 12080
rect 44541 12114 44741 12130
rect 44541 12080 44557 12114
rect 44725 12080 44741 12114
rect 44541 12033 44741 12080
rect 44913 12114 45113 12130
rect 44913 12080 44929 12114
rect 45097 12080 45113 12114
rect 44913 12033 45113 12080
rect 45285 12114 45485 12130
rect 45285 12080 45301 12114
rect 45469 12080 45485 12114
rect 45285 12033 45485 12080
rect 45657 12114 45857 12130
rect 45657 12080 45673 12114
rect 45841 12080 45857 12114
rect 45657 12033 45857 12080
rect 46029 12114 46229 12130
rect 46029 12080 46045 12114
rect 46213 12080 46229 12114
rect 46029 12033 46229 12080
rect 46401 12114 46601 12130
rect 46401 12080 46417 12114
rect 46585 12080 46601 12114
rect 46401 12033 46601 12080
rect 46773 12114 46973 12130
rect 46773 12080 46789 12114
rect 46957 12080 46973 12114
rect 46773 12033 46973 12080
rect 47145 12114 47345 12130
rect 47145 12080 47161 12114
rect 47329 12080 47345 12114
rect 47145 12033 47345 12080
rect 47517 12114 47717 12130
rect 47517 12080 47533 12114
rect 47701 12080 47717 12114
rect 47517 12033 47717 12080
rect 47889 12114 48089 12130
rect 47889 12080 47905 12114
rect 48073 12080 48089 12114
rect 47889 12033 48089 12080
rect 48261 12114 48461 12130
rect 48261 12080 48277 12114
rect 48445 12080 48461 12114
rect 48261 12033 48461 12080
rect 48633 12114 48833 12130
rect 48633 12080 48649 12114
rect 48817 12080 48833 12114
rect 48633 12033 48833 12080
rect 49005 12114 49205 12130
rect 49005 12080 49021 12114
rect 49189 12080 49205 12114
rect 49005 12033 49205 12080
rect 49377 12114 49577 12130
rect 49377 12080 49393 12114
rect 49561 12080 49577 12114
rect 49377 12033 49577 12080
rect 49749 12114 49949 12130
rect 49749 12080 49765 12114
rect 49933 12080 49949 12114
rect 49749 12033 49949 12080
rect 50121 12114 50321 12130
rect 50121 12080 50137 12114
rect 50305 12080 50321 12114
rect 50121 12033 50321 12080
rect 50493 12114 50693 12130
rect 50493 12080 50509 12114
rect 50677 12080 50693 12114
rect 50493 12033 50693 12080
rect 50865 12114 51065 12130
rect 50865 12080 50881 12114
rect 51049 12080 51065 12114
rect 50865 12033 51065 12080
rect 39333 11586 39533 11633
rect 39333 11552 39349 11586
rect 39517 11552 39533 11586
rect 39333 11536 39533 11552
rect 39705 11586 39905 11633
rect 39705 11552 39721 11586
rect 39889 11552 39905 11586
rect 39705 11536 39905 11552
rect 40077 11586 40277 11633
rect 40077 11552 40093 11586
rect 40261 11552 40277 11586
rect 40077 11536 40277 11552
rect 40449 11586 40649 11633
rect 40449 11552 40465 11586
rect 40633 11552 40649 11586
rect 40449 11536 40649 11552
rect 40821 11586 41021 11633
rect 40821 11552 40837 11586
rect 41005 11552 41021 11586
rect 40821 11536 41021 11552
rect 41193 11586 41393 11633
rect 41193 11552 41209 11586
rect 41377 11552 41393 11586
rect 41193 11536 41393 11552
rect 41565 11586 41765 11633
rect 41565 11552 41581 11586
rect 41749 11552 41765 11586
rect 41565 11536 41765 11552
rect 41937 11586 42137 11633
rect 41937 11552 41953 11586
rect 42121 11552 42137 11586
rect 41937 11536 42137 11552
rect 42309 11586 42509 11633
rect 42309 11552 42325 11586
rect 42493 11552 42509 11586
rect 42309 11536 42509 11552
rect 42681 11586 42881 11633
rect 42681 11552 42697 11586
rect 42865 11552 42881 11586
rect 42681 11536 42881 11552
rect 43053 11586 43253 11633
rect 43053 11552 43069 11586
rect 43237 11552 43253 11586
rect 43053 11536 43253 11552
rect 43425 11586 43625 11633
rect 43425 11552 43441 11586
rect 43609 11552 43625 11586
rect 43425 11536 43625 11552
rect 43797 11586 43997 11633
rect 43797 11552 43813 11586
rect 43981 11552 43997 11586
rect 43797 11536 43997 11552
rect 44169 11586 44369 11633
rect 44169 11552 44185 11586
rect 44353 11552 44369 11586
rect 44169 11536 44369 11552
rect 44541 11586 44741 11633
rect 44541 11552 44557 11586
rect 44725 11552 44741 11586
rect 44541 11536 44741 11552
rect 44913 11586 45113 11633
rect 44913 11552 44929 11586
rect 45097 11552 45113 11586
rect 44913 11536 45113 11552
rect 45285 11586 45485 11633
rect 45285 11552 45301 11586
rect 45469 11552 45485 11586
rect 45285 11536 45485 11552
rect 45657 11586 45857 11633
rect 45657 11552 45673 11586
rect 45841 11552 45857 11586
rect 45657 11536 45857 11552
rect 46029 11586 46229 11633
rect 46029 11552 46045 11586
rect 46213 11552 46229 11586
rect 46029 11536 46229 11552
rect 46401 11586 46601 11633
rect 46401 11552 46417 11586
rect 46585 11552 46601 11586
rect 46401 11536 46601 11552
rect 46773 11586 46973 11633
rect 46773 11552 46789 11586
rect 46957 11552 46973 11586
rect 46773 11536 46973 11552
rect 47145 11586 47345 11633
rect 47145 11552 47161 11586
rect 47329 11552 47345 11586
rect 47145 11536 47345 11552
rect 47517 11586 47717 11633
rect 47517 11552 47533 11586
rect 47701 11552 47717 11586
rect 47517 11536 47717 11552
rect 47889 11586 48089 11633
rect 47889 11552 47905 11586
rect 48073 11552 48089 11586
rect 47889 11536 48089 11552
rect 48261 11586 48461 11633
rect 48261 11552 48277 11586
rect 48445 11552 48461 11586
rect 48261 11536 48461 11552
rect 48633 11586 48833 11633
rect 48633 11552 48649 11586
rect 48817 11552 48833 11586
rect 48633 11536 48833 11552
rect 49005 11586 49205 11633
rect 49005 11552 49021 11586
rect 49189 11552 49205 11586
rect 49005 11536 49205 11552
rect 49377 11586 49577 11633
rect 49377 11552 49393 11586
rect 49561 11552 49577 11586
rect 49377 11536 49577 11552
rect 49749 11586 49949 11633
rect 49749 11552 49765 11586
rect 49933 11552 49949 11586
rect 49749 11536 49949 11552
rect 50121 11586 50321 11633
rect 50121 11552 50137 11586
rect 50305 11552 50321 11586
rect 50121 11536 50321 11552
rect 50493 11586 50693 11633
rect 50493 11552 50509 11586
rect 50677 11552 50693 11586
rect 50493 11536 50693 11552
rect 50865 11586 51065 11633
rect 50865 11552 50881 11586
rect 51049 11552 51065 11586
rect 50865 11536 51065 11552
rect 39333 11478 39533 11494
rect 39333 11444 39349 11478
rect 39517 11444 39533 11478
rect 39333 11397 39533 11444
rect 39705 11478 39905 11494
rect 39705 11444 39721 11478
rect 39889 11444 39905 11478
rect 39705 11397 39905 11444
rect 40077 11478 40277 11494
rect 40077 11444 40093 11478
rect 40261 11444 40277 11478
rect 40077 11397 40277 11444
rect 40449 11478 40649 11494
rect 40449 11444 40465 11478
rect 40633 11444 40649 11478
rect 40449 11397 40649 11444
rect 40821 11478 41021 11494
rect 40821 11444 40837 11478
rect 41005 11444 41021 11478
rect 40821 11397 41021 11444
rect 41193 11478 41393 11494
rect 41193 11444 41209 11478
rect 41377 11444 41393 11478
rect 41193 11397 41393 11444
rect 41565 11478 41765 11494
rect 41565 11444 41581 11478
rect 41749 11444 41765 11478
rect 41565 11397 41765 11444
rect 41937 11478 42137 11494
rect 41937 11444 41953 11478
rect 42121 11444 42137 11478
rect 41937 11397 42137 11444
rect 42309 11478 42509 11494
rect 42309 11444 42325 11478
rect 42493 11444 42509 11478
rect 42309 11397 42509 11444
rect 42681 11478 42881 11494
rect 42681 11444 42697 11478
rect 42865 11444 42881 11478
rect 42681 11397 42881 11444
rect 43053 11478 43253 11494
rect 43053 11444 43069 11478
rect 43237 11444 43253 11478
rect 43053 11397 43253 11444
rect 43425 11478 43625 11494
rect 43425 11444 43441 11478
rect 43609 11444 43625 11478
rect 43425 11397 43625 11444
rect 43797 11478 43997 11494
rect 43797 11444 43813 11478
rect 43981 11444 43997 11478
rect 43797 11397 43997 11444
rect 44169 11478 44369 11494
rect 44169 11444 44185 11478
rect 44353 11444 44369 11478
rect 44169 11397 44369 11444
rect 44541 11478 44741 11494
rect 44541 11444 44557 11478
rect 44725 11444 44741 11478
rect 44541 11397 44741 11444
rect 44913 11478 45113 11494
rect 44913 11444 44929 11478
rect 45097 11444 45113 11478
rect 44913 11397 45113 11444
rect 45285 11478 45485 11494
rect 45285 11444 45301 11478
rect 45469 11444 45485 11478
rect 45285 11397 45485 11444
rect 45657 11478 45857 11494
rect 45657 11444 45673 11478
rect 45841 11444 45857 11478
rect 45657 11397 45857 11444
rect 46029 11478 46229 11494
rect 46029 11444 46045 11478
rect 46213 11444 46229 11478
rect 46029 11397 46229 11444
rect 46401 11478 46601 11494
rect 46401 11444 46417 11478
rect 46585 11444 46601 11478
rect 46401 11397 46601 11444
rect 46773 11478 46973 11494
rect 46773 11444 46789 11478
rect 46957 11444 46973 11478
rect 46773 11397 46973 11444
rect 47145 11478 47345 11494
rect 47145 11444 47161 11478
rect 47329 11444 47345 11478
rect 47145 11397 47345 11444
rect 47517 11478 47717 11494
rect 47517 11444 47533 11478
rect 47701 11444 47717 11478
rect 47517 11397 47717 11444
rect 47889 11478 48089 11494
rect 47889 11444 47905 11478
rect 48073 11444 48089 11478
rect 47889 11397 48089 11444
rect 48261 11478 48461 11494
rect 48261 11444 48277 11478
rect 48445 11444 48461 11478
rect 48261 11397 48461 11444
rect 48633 11478 48833 11494
rect 48633 11444 48649 11478
rect 48817 11444 48833 11478
rect 48633 11397 48833 11444
rect 49005 11478 49205 11494
rect 49005 11444 49021 11478
rect 49189 11444 49205 11478
rect 49005 11397 49205 11444
rect 49377 11478 49577 11494
rect 49377 11444 49393 11478
rect 49561 11444 49577 11478
rect 49377 11397 49577 11444
rect 49749 11478 49949 11494
rect 49749 11444 49765 11478
rect 49933 11444 49949 11478
rect 49749 11397 49949 11444
rect 50121 11478 50321 11494
rect 50121 11444 50137 11478
rect 50305 11444 50321 11478
rect 50121 11397 50321 11444
rect 50493 11478 50693 11494
rect 50493 11444 50509 11478
rect 50677 11444 50693 11478
rect 50493 11397 50693 11444
rect 50865 11478 51065 11494
rect 50865 11444 50881 11478
rect 51049 11444 51065 11478
rect 50865 11397 51065 11444
rect 39333 10950 39533 10997
rect 39333 10916 39349 10950
rect 39517 10916 39533 10950
rect 39333 10900 39533 10916
rect 39705 10950 39905 10997
rect 39705 10916 39721 10950
rect 39889 10916 39905 10950
rect 39705 10900 39905 10916
rect 40077 10950 40277 10997
rect 40077 10916 40093 10950
rect 40261 10916 40277 10950
rect 40077 10900 40277 10916
rect 40449 10950 40649 10997
rect 40449 10916 40465 10950
rect 40633 10916 40649 10950
rect 40449 10900 40649 10916
rect 40821 10950 41021 10997
rect 40821 10916 40837 10950
rect 41005 10916 41021 10950
rect 40821 10900 41021 10916
rect 41193 10950 41393 10997
rect 41193 10916 41209 10950
rect 41377 10916 41393 10950
rect 41193 10900 41393 10916
rect 41565 10950 41765 10997
rect 41565 10916 41581 10950
rect 41749 10916 41765 10950
rect 41565 10900 41765 10916
rect 41937 10950 42137 10997
rect 41937 10916 41953 10950
rect 42121 10916 42137 10950
rect 41937 10900 42137 10916
rect 42309 10950 42509 10997
rect 42309 10916 42325 10950
rect 42493 10916 42509 10950
rect 42309 10900 42509 10916
rect 42681 10950 42881 10997
rect 42681 10916 42697 10950
rect 42865 10916 42881 10950
rect 42681 10900 42881 10916
rect 43053 10950 43253 10997
rect 43053 10916 43069 10950
rect 43237 10916 43253 10950
rect 43053 10900 43253 10916
rect 43425 10950 43625 10997
rect 43425 10916 43441 10950
rect 43609 10916 43625 10950
rect 43425 10900 43625 10916
rect 43797 10950 43997 10997
rect 43797 10916 43813 10950
rect 43981 10916 43997 10950
rect 43797 10900 43997 10916
rect 44169 10950 44369 10997
rect 44169 10916 44185 10950
rect 44353 10916 44369 10950
rect 44169 10900 44369 10916
rect 44541 10950 44741 10997
rect 44541 10916 44557 10950
rect 44725 10916 44741 10950
rect 44541 10900 44741 10916
rect 44913 10950 45113 10997
rect 44913 10916 44929 10950
rect 45097 10916 45113 10950
rect 44913 10900 45113 10916
rect 45285 10950 45485 10997
rect 45285 10916 45301 10950
rect 45469 10916 45485 10950
rect 45285 10900 45485 10916
rect 45657 10950 45857 10997
rect 45657 10916 45673 10950
rect 45841 10916 45857 10950
rect 45657 10900 45857 10916
rect 46029 10950 46229 10997
rect 46029 10916 46045 10950
rect 46213 10916 46229 10950
rect 46029 10900 46229 10916
rect 46401 10950 46601 10997
rect 46401 10916 46417 10950
rect 46585 10916 46601 10950
rect 46401 10900 46601 10916
rect 46773 10950 46973 10997
rect 46773 10916 46789 10950
rect 46957 10916 46973 10950
rect 46773 10900 46973 10916
rect 47145 10950 47345 10997
rect 47145 10916 47161 10950
rect 47329 10916 47345 10950
rect 47145 10900 47345 10916
rect 47517 10950 47717 10997
rect 47517 10916 47533 10950
rect 47701 10916 47717 10950
rect 47517 10900 47717 10916
rect 47889 10950 48089 10997
rect 47889 10916 47905 10950
rect 48073 10916 48089 10950
rect 47889 10900 48089 10916
rect 48261 10950 48461 10997
rect 48261 10916 48277 10950
rect 48445 10916 48461 10950
rect 48261 10900 48461 10916
rect 48633 10950 48833 10997
rect 48633 10916 48649 10950
rect 48817 10916 48833 10950
rect 48633 10900 48833 10916
rect 49005 10950 49205 10997
rect 49005 10916 49021 10950
rect 49189 10916 49205 10950
rect 49005 10900 49205 10916
rect 49377 10950 49577 10997
rect 49377 10916 49393 10950
rect 49561 10916 49577 10950
rect 49377 10900 49577 10916
rect 49749 10950 49949 10997
rect 49749 10916 49765 10950
rect 49933 10916 49949 10950
rect 49749 10900 49949 10916
rect 50121 10950 50321 10997
rect 50121 10916 50137 10950
rect 50305 10916 50321 10950
rect 50121 10900 50321 10916
rect 50493 10950 50693 10997
rect 50493 10916 50509 10950
rect 50677 10916 50693 10950
rect 50493 10900 50693 10916
rect 50865 10950 51065 10997
rect 50865 10916 50881 10950
rect 51049 10916 51065 10950
rect 50865 10900 51065 10916
rect 39333 8949 39533 8965
rect 39333 8915 39349 8949
rect 39517 8915 39533 8949
rect 39333 8868 39533 8915
rect 39705 8949 39905 8965
rect 39705 8915 39721 8949
rect 39889 8915 39905 8949
rect 39705 8868 39905 8915
rect 40077 8949 40277 8965
rect 40077 8915 40093 8949
rect 40261 8915 40277 8949
rect 40077 8868 40277 8915
rect 40449 8949 40649 8965
rect 40449 8915 40465 8949
rect 40633 8915 40649 8949
rect 40449 8868 40649 8915
rect 40821 8949 41021 8965
rect 40821 8915 40837 8949
rect 41005 8915 41021 8949
rect 40821 8868 41021 8915
rect 41193 8949 41393 8965
rect 41193 8915 41209 8949
rect 41377 8915 41393 8949
rect 41193 8868 41393 8915
rect 41565 8949 41765 8965
rect 41565 8915 41581 8949
rect 41749 8915 41765 8949
rect 41565 8868 41765 8915
rect 41937 8949 42137 8965
rect 41937 8915 41953 8949
rect 42121 8915 42137 8949
rect 41937 8868 42137 8915
rect 42309 8949 42509 8965
rect 42309 8915 42325 8949
rect 42493 8915 42509 8949
rect 42309 8868 42509 8915
rect 42681 8949 42881 8965
rect 42681 8915 42697 8949
rect 42865 8915 42881 8949
rect 42681 8868 42881 8915
rect 43053 8949 43253 8965
rect 43053 8915 43069 8949
rect 43237 8915 43253 8949
rect 43053 8868 43253 8915
rect 43425 8949 43625 8965
rect 43425 8915 43441 8949
rect 43609 8915 43625 8949
rect 43425 8868 43625 8915
rect 43797 8949 43997 8965
rect 43797 8915 43813 8949
rect 43981 8915 43997 8949
rect 43797 8868 43997 8915
rect 44169 8949 44369 8965
rect 44169 8915 44185 8949
rect 44353 8915 44369 8949
rect 44169 8868 44369 8915
rect 44541 8949 44741 8965
rect 44541 8915 44557 8949
rect 44725 8915 44741 8949
rect 44541 8868 44741 8915
rect 44913 8949 45113 8965
rect 44913 8915 44929 8949
rect 45097 8915 45113 8949
rect 44913 8868 45113 8915
rect 45285 8949 45485 8965
rect 45285 8915 45301 8949
rect 45469 8915 45485 8949
rect 45285 8868 45485 8915
rect 45657 8949 45857 8965
rect 45657 8915 45673 8949
rect 45841 8915 45857 8949
rect 45657 8868 45857 8915
rect 46029 8949 46229 8965
rect 46029 8915 46045 8949
rect 46213 8915 46229 8949
rect 46029 8868 46229 8915
rect 46401 8949 46601 8965
rect 46401 8915 46417 8949
rect 46585 8915 46601 8949
rect 46401 8868 46601 8915
rect 46773 8949 46973 8965
rect 46773 8915 46789 8949
rect 46957 8915 46973 8949
rect 46773 8868 46973 8915
rect 47145 8949 47345 8965
rect 47145 8915 47161 8949
rect 47329 8915 47345 8949
rect 47145 8868 47345 8915
rect 47517 8949 47717 8965
rect 47517 8915 47533 8949
rect 47701 8915 47717 8949
rect 47517 8868 47717 8915
rect 47889 8949 48089 8965
rect 47889 8915 47905 8949
rect 48073 8915 48089 8949
rect 47889 8868 48089 8915
rect 48261 8949 48461 8965
rect 48261 8915 48277 8949
rect 48445 8915 48461 8949
rect 48261 8868 48461 8915
rect 48633 8949 48833 8965
rect 48633 8915 48649 8949
rect 48817 8915 48833 8949
rect 48633 8868 48833 8915
rect 49005 8949 49205 8965
rect 49005 8915 49021 8949
rect 49189 8915 49205 8949
rect 49005 8868 49205 8915
rect 49377 8949 49577 8965
rect 49377 8915 49393 8949
rect 49561 8915 49577 8949
rect 49377 8868 49577 8915
rect 49749 8949 49949 8965
rect 49749 8915 49765 8949
rect 49933 8915 49949 8949
rect 49749 8868 49949 8915
rect 50121 8949 50321 8965
rect 50121 8915 50137 8949
rect 50305 8915 50321 8949
rect 50121 8868 50321 8915
rect 50493 8949 50693 8965
rect 50493 8915 50509 8949
rect 50677 8915 50693 8949
rect 50493 8868 50693 8915
rect 50865 8949 51065 8965
rect 50865 8915 50881 8949
rect 51049 8915 51065 8949
rect 50865 8868 51065 8915
rect 39333 8421 39533 8468
rect 39333 8387 39349 8421
rect 39517 8387 39533 8421
rect 39333 8371 39533 8387
rect 39705 8421 39905 8468
rect 39705 8387 39721 8421
rect 39889 8387 39905 8421
rect 39705 8371 39905 8387
rect 40077 8421 40277 8468
rect 40077 8387 40093 8421
rect 40261 8387 40277 8421
rect 40077 8371 40277 8387
rect 40449 8421 40649 8468
rect 40449 8387 40465 8421
rect 40633 8387 40649 8421
rect 40449 8371 40649 8387
rect 40821 8421 41021 8468
rect 40821 8387 40837 8421
rect 41005 8387 41021 8421
rect 40821 8371 41021 8387
rect 41193 8421 41393 8468
rect 41193 8387 41209 8421
rect 41377 8387 41393 8421
rect 41193 8371 41393 8387
rect 41565 8421 41765 8468
rect 41565 8387 41581 8421
rect 41749 8387 41765 8421
rect 41565 8371 41765 8387
rect 41937 8421 42137 8468
rect 41937 8387 41953 8421
rect 42121 8387 42137 8421
rect 41937 8371 42137 8387
rect 42309 8421 42509 8468
rect 42309 8387 42325 8421
rect 42493 8387 42509 8421
rect 42309 8371 42509 8387
rect 42681 8421 42881 8468
rect 42681 8387 42697 8421
rect 42865 8387 42881 8421
rect 42681 8371 42881 8387
rect 43053 8421 43253 8468
rect 43053 8387 43069 8421
rect 43237 8387 43253 8421
rect 43053 8371 43253 8387
rect 43425 8421 43625 8468
rect 43425 8387 43441 8421
rect 43609 8387 43625 8421
rect 43425 8371 43625 8387
rect 43797 8421 43997 8468
rect 43797 8387 43813 8421
rect 43981 8387 43997 8421
rect 43797 8371 43997 8387
rect 44169 8421 44369 8468
rect 44169 8387 44185 8421
rect 44353 8387 44369 8421
rect 44169 8371 44369 8387
rect 44541 8421 44741 8468
rect 44541 8387 44557 8421
rect 44725 8387 44741 8421
rect 44541 8371 44741 8387
rect 44913 8421 45113 8468
rect 44913 8387 44929 8421
rect 45097 8387 45113 8421
rect 44913 8371 45113 8387
rect 45285 8421 45485 8468
rect 45285 8387 45301 8421
rect 45469 8387 45485 8421
rect 45285 8371 45485 8387
rect 45657 8421 45857 8468
rect 45657 8387 45673 8421
rect 45841 8387 45857 8421
rect 45657 8371 45857 8387
rect 46029 8421 46229 8468
rect 46029 8387 46045 8421
rect 46213 8387 46229 8421
rect 46029 8371 46229 8387
rect 46401 8421 46601 8468
rect 46401 8387 46417 8421
rect 46585 8387 46601 8421
rect 46401 8371 46601 8387
rect 46773 8421 46973 8468
rect 46773 8387 46789 8421
rect 46957 8387 46973 8421
rect 46773 8371 46973 8387
rect 47145 8421 47345 8468
rect 47145 8387 47161 8421
rect 47329 8387 47345 8421
rect 47145 8371 47345 8387
rect 47517 8421 47717 8468
rect 47517 8387 47533 8421
rect 47701 8387 47717 8421
rect 47517 8371 47717 8387
rect 47889 8421 48089 8468
rect 47889 8387 47905 8421
rect 48073 8387 48089 8421
rect 47889 8371 48089 8387
rect 48261 8421 48461 8468
rect 48261 8387 48277 8421
rect 48445 8387 48461 8421
rect 48261 8371 48461 8387
rect 48633 8421 48833 8468
rect 48633 8387 48649 8421
rect 48817 8387 48833 8421
rect 48633 8371 48833 8387
rect 49005 8421 49205 8468
rect 49005 8387 49021 8421
rect 49189 8387 49205 8421
rect 49005 8371 49205 8387
rect 49377 8421 49577 8468
rect 49377 8387 49393 8421
rect 49561 8387 49577 8421
rect 49377 8371 49577 8387
rect 49749 8421 49949 8468
rect 49749 8387 49765 8421
rect 49933 8387 49949 8421
rect 49749 8371 49949 8387
rect 50121 8421 50321 8468
rect 50121 8387 50137 8421
rect 50305 8387 50321 8421
rect 50121 8371 50321 8387
rect 50493 8421 50693 8468
rect 50493 8387 50509 8421
rect 50677 8387 50693 8421
rect 50493 8371 50693 8387
rect 50865 8421 51065 8468
rect 50865 8387 50881 8421
rect 51049 8387 51065 8421
rect 50865 8371 51065 8387
rect 39333 8313 39533 8329
rect 39333 8279 39349 8313
rect 39517 8279 39533 8313
rect 39333 8232 39533 8279
rect 39705 8313 39905 8329
rect 39705 8279 39721 8313
rect 39889 8279 39905 8313
rect 39705 8232 39905 8279
rect 40077 8313 40277 8329
rect 40077 8279 40093 8313
rect 40261 8279 40277 8313
rect 40077 8232 40277 8279
rect 40449 8313 40649 8329
rect 40449 8279 40465 8313
rect 40633 8279 40649 8313
rect 40449 8232 40649 8279
rect 40821 8313 41021 8329
rect 40821 8279 40837 8313
rect 41005 8279 41021 8313
rect 40821 8232 41021 8279
rect 41193 8313 41393 8329
rect 41193 8279 41209 8313
rect 41377 8279 41393 8313
rect 41193 8232 41393 8279
rect 41565 8313 41765 8329
rect 41565 8279 41581 8313
rect 41749 8279 41765 8313
rect 41565 8232 41765 8279
rect 41937 8313 42137 8329
rect 41937 8279 41953 8313
rect 42121 8279 42137 8313
rect 41937 8232 42137 8279
rect 42309 8313 42509 8329
rect 42309 8279 42325 8313
rect 42493 8279 42509 8313
rect 42309 8232 42509 8279
rect 42681 8313 42881 8329
rect 42681 8279 42697 8313
rect 42865 8279 42881 8313
rect 42681 8232 42881 8279
rect 43053 8313 43253 8329
rect 43053 8279 43069 8313
rect 43237 8279 43253 8313
rect 43053 8232 43253 8279
rect 43425 8313 43625 8329
rect 43425 8279 43441 8313
rect 43609 8279 43625 8313
rect 43425 8232 43625 8279
rect 43797 8313 43997 8329
rect 43797 8279 43813 8313
rect 43981 8279 43997 8313
rect 43797 8232 43997 8279
rect 44169 8313 44369 8329
rect 44169 8279 44185 8313
rect 44353 8279 44369 8313
rect 44169 8232 44369 8279
rect 44541 8313 44741 8329
rect 44541 8279 44557 8313
rect 44725 8279 44741 8313
rect 44541 8232 44741 8279
rect 44913 8313 45113 8329
rect 44913 8279 44929 8313
rect 45097 8279 45113 8313
rect 44913 8232 45113 8279
rect 45285 8313 45485 8329
rect 45285 8279 45301 8313
rect 45469 8279 45485 8313
rect 45285 8232 45485 8279
rect 45657 8313 45857 8329
rect 45657 8279 45673 8313
rect 45841 8279 45857 8313
rect 45657 8232 45857 8279
rect 46029 8313 46229 8329
rect 46029 8279 46045 8313
rect 46213 8279 46229 8313
rect 46029 8232 46229 8279
rect 46401 8313 46601 8329
rect 46401 8279 46417 8313
rect 46585 8279 46601 8313
rect 46401 8232 46601 8279
rect 46773 8313 46973 8329
rect 46773 8279 46789 8313
rect 46957 8279 46973 8313
rect 46773 8232 46973 8279
rect 47145 8313 47345 8329
rect 47145 8279 47161 8313
rect 47329 8279 47345 8313
rect 47145 8232 47345 8279
rect 47517 8313 47717 8329
rect 47517 8279 47533 8313
rect 47701 8279 47717 8313
rect 47517 8232 47717 8279
rect 47889 8313 48089 8329
rect 47889 8279 47905 8313
rect 48073 8279 48089 8313
rect 47889 8232 48089 8279
rect 48261 8313 48461 8329
rect 48261 8279 48277 8313
rect 48445 8279 48461 8313
rect 48261 8232 48461 8279
rect 48633 8313 48833 8329
rect 48633 8279 48649 8313
rect 48817 8279 48833 8313
rect 48633 8232 48833 8279
rect 49005 8313 49205 8329
rect 49005 8279 49021 8313
rect 49189 8279 49205 8313
rect 49005 8232 49205 8279
rect 49377 8313 49577 8329
rect 49377 8279 49393 8313
rect 49561 8279 49577 8313
rect 49377 8232 49577 8279
rect 49749 8313 49949 8329
rect 49749 8279 49765 8313
rect 49933 8279 49949 8313
rect 49749 8232 49949 8279
rect 50121 8313 50321 8329
rect 50121 8279 50137 8313
rect 50305 8279 50321 8313
rect 50121 8232 50321 8279
rect 50493 8313 50693 8329
rect 50493 8279 50509 8313
rect 50677 8279 50693 8313
rect 50493 8232 50693 8279
rect 50865 8313 51065 8329
rect 50865 8279 50881 8313
rect 51049 8279 51065 8313
rect 50865 8232 51065 8279
rect 39333 7785 39533 7832
rect 39333 7751 39349 7785
rect 39517 7751 39533 7785
rect 39333 7735 39533 7751
rect 39705 7785 39905 7832
rect 39705 7751 39721 7785
rect 39889 7751 39905 7785
rect 39705 7735 39905 7751
rect 40077 7785 40277 7832
rect 40077 7751 40093 7785
rect 40261 7751 40277 7785
rect 40077 7735 40277 7751
rect 40449 7785 40649 7832
rect 40449 7751 40465 7785
rect 40633 7751 40649 7785
rect 40449 7735 40649 7751
rect 40821 7785 41021 7832
rect 40821 7751 40837 7785
rect 41005 7751 41021 7785
rect 40821 7735 41021 7751
rect 41193 7785 41393 7832
rect 41193 7751 41209 7785
rect 41377 7751 41393 7785
rect 41193 7735 41393 7751
rect 41565 7785 41765 7832
rect 41565 7751 41581 7785
rect 41749 7751 41765 7785
rect 41565 7735 41765 7751
rect 41937 7785 42137 7832
rect 41937 7751 41953 7785
rect 42121 7751 42137 7785
rect 41937 7735 42137 7751
rect 42309 7785 42509 7832
rect 42309 7751 42325 7785
rect 42493 7751 42509 7785
rect 42309 7735 42509 7751
rect 42681 7785 42881 7832
rect 42681 7751 42697 7785
rect 42865 7751 42881 7785
rect 42681 7735 42881 7751
rect 43053 7785 43253 7832
rect 43053 7751 43069 7785
rect 43237 7751 43253 7785
rect 43053 7735 43253 7751
rect 43425 7785 43625 7832
rect 43425 7751 43441 7785
rect 43609 7751 43625 7785
rect 43425 7735 43625 7751
rect 43797 7785 43997 7832
rect 43797 7751 43813 7785
rect 43981 7751 43997 7785
rect 43797 7735 43997 7751
rect 44169 7785 44369 7832
rect 44169 7751 44185 7785
rect 44353 7751 44369 7785
rect 44169 7735 44369 7751
rect 44541 7785 44741 7832
rect 44541 7751 44557 7785
rect 44725 7751 44741 7785
rect 44541 7735 44741 7751
rect 44913 7785 45113 7832
rect 44913 7751 44929 7785
rect 45097 7751 45113 7785
rect 44913 7735 45113 7751
rect 45285 7785 45485 7832
rect 45285 7751 45301 7785
rect 45469 7751 45485 7785
rect 45285 7735 45485 7751
rect 45657 7785 45857 7832
rect 45657 7751 45673 7785
rect 45841 7751 45857 7785
rect 45657 7735 45857 7751
rect 46029 7785 46229 7832
rect 46029 7751 46045 7785
rect 46213 7751 46229 7785
rect 46029 7735 46229 7751
rect 46401 7785 46601 7832
rect 46401 7751 46417 7785
rect 46585 7751 46601 7785
rect 46401 7735 46601 7751
rect 46773 7785 46973 7832
rect 46773 7751 46789 7785
rect 46957 7751 46973 7785
rect 46773 7735 46973 7751
rect 47145 7785 47345 7832
rect 47145 7751 47161 7785
rect 47329 7751 47345 7785
rect 47145 7735 47345 7751
rect 47517 7785 47717 7832
rect 47517 7751 47533 7785
rect 47701 7751 47717 7785
rect 47517 7735 47717 7751
rect 47889 7785 48089 7832
rect 47889 7751 47905 7785
rect 48073 7751 48089 7785
rect 47889 7735 48089 7751
rect 48261 7785 48461 7832
rect 48261 7751 48277 7785
rect 48445 7751 48461 7785
rect 48261 7735 48461 7751
rect 48633 7785 48833 7832
rect 48633 7751 48649 7785
rect 48817 7751 48833 7785
rect 48633 7735 48833 7751
rect 49005 7785 49205 7832
rect 49005 7751 49021 7785
rect 49189 7751 49205 7785
rect 49005 7735 49205 7751
rect 49377 7785 49577 7832
rect 49377 7751 49393 7785
rect 49561 7751 49577 7785
rect 49377 7735 49577 7751
rect 49749 7785 49949 7832
rect 49749 7751 49765 7785
rect 49933 7751 49949 7785
rect 49749 7735 49949 7751
rect 50121 7785 50321 7832
rect 50121 7751 50137 7785
rect 50305 7751 50321 7785
rect 50121 7735 50321 7751
rect 50493 7785 50693 7832
rect 50493 7751 50509 7785
rect 50677 7751 50693 7785
rect 50493 7735 50693 7751
rect 50865 7785 51065 7832
rect 50865 7751 50881 7785
rect 51049 7751 51065 7785
rect 50865 7735 51065 7751
rect 39333 7677 39533 7693
rect 39333 7643 39349 7677
rect 39517 7643 39533 7677
rect 39333 7596 39533 7643
rect 39705 7677 39905 7693
rect 39705 7643 39721 7677
rect 39889 7643 39905 7677
rect 39705 7596 39905 7643
rect 40077 7677 40277 7693
rect 40077 7643 40093 7677
rect 40261 7643 40277 7677
rect 40077 7596 40277 7643
rect 40449 7677 40649 7693
rect 40449 7643 40465 7677
rect 40633 7643 40649 7677
rect 40449 7596 40649 7643
rect 40821 7677 41021 7693
rect 40821 7643 40837 7677
rect 41005 7643 41021 7677
rect 40821 7596 41021 7643
rect 41193 7677 41393 7693
rect 41193 7643 41209 7677
rect 41377 7643 41393 7677
rect 41193 7596 41393 7643
rect 41565 7677 41765 7693
rect 41565 7643 41581 7677
rect 41749 7643 41765 7677
rect 41565 7596 41765 7643
rect 41937 7677 42137 7693
rect 41937 7643 41953 7677
rect 42121 7643 42137 7677
rect 41937 7596 42137 7643
rect 42309 7677 42509 7693
rect 42309 7643 42325 7677
rect 42493 7643 42509 7677
rect 42309 7596 42509 7643
rect 42681 7677 42881 7693
rect 42681 7643 42697 7677
rect 42865 7643 42881 7677
rect 42681 7596 42881 7643
rect 43053 7677 43253 7693
rect 43053 7643 43069 7677
rect 43237 7643 43253 7677
rect 43053 7596 43253 7643
rect 43425 7677 43625 7693
rect 43425 7643 43441 7677
rect 43609 7643 43625 7677
rect 43425 7596 43625 7643
rect 43797 7677 43997 7693
rect 43797 7643 43813 7677
rect 43981 7643 43997 7677
rect 43797 7596 43997 7643
rect 44169 7677 44369 7693
rect 44169 7643 44185 7677
rect 44353 7643 44369 7677
rect 44169 7596 44369 7643
rect 44541 7677 44741 7693
rect 44541 7643 44557 7677
rect 44725 7643 44741 7677
rect 44541 7596 44741 7643
rect 44913 7677 45113 7693
rect 44913 7643 44929 7677
rect 45097 7643 45113 7677
rect 44913 7596 45113 7643
rect 45285 7677 45485 7693
rect 45285 7643 45301 7677
rect 45469 7643 45485 7677
rect 45285 7596 45485 7643
rect 45657 7677 45857 7693
rect 45657 7643 45673 7677
rect 45841 7643 45857 7677
rect 45657 7596 45857 7643
rect 46029 7677 46229 7693
rect 46029 7643 46045 7677
rect 46213 7643 46229 7677
rect 46029 7596 46229 7643
rect 46401 7677 46601 7693
rect 46401 7643 46417 7677
rect 46585 7643 46601 7677
rect 46401 7596 46601 7643
rect 46773 7677 46973 7693
rect 46773 7643 46789 7677
rect 46957 7643 46973 7677
rect 46773 7596 46973 7643
rect 47145 7677 47345 7693
rect 47145 7643 47161 7677
rect 47329 7643 47345 7677
rect 47145 7596 47345 7643
rect 47517 7677 47717 7693
rect 47517 7643 47533 7677
rect 47701 7643 47717 7677
rect 47517 7596 47717 7643
rect 47889 7677 48089 7693
rect 47889 7643 47905 7677
rect 48073 7643 48089 7677
rect 47889 7596 48089 7643
rect 48261 7677 48461 7693
rect 48261 7643 48277 7677
rect 48445 7643 48461 7677
rect 48261 7596 48461 7643
rect 48633 7677 48833 7693
rect 48633 7643 48649 7677
rect 48817 7643 48833 7677
rect 48633 7596 48833 7643
rect 49005 7677 49205 7693
rect 49005 7643 49021 7677
rect 49189 7643 49205 7677
rect 49005 7596 49205 7643
rect 49377 7677 49577 7693
rect 49377 7643 49393 7677
rect 49561 7643 49577 7677
rect 49377 7596 49577 7643
rect 49749 7677 49949 7693
rect 49749 7643 49765 7677
rect 49933 7643 49949 7677
rect 49749 7596 49949 7643
rect 50121 7677 50321 7693
rect 50121 7643 50137 7677
rect 50305 7643 50321 7677
rect 50121 7596 50321 7643
rect 50493 7677 50693 7693
rect 50493 7643 50509 7677
rect 50677 7643 50693 7677
rect 50493 7596 50693 7643
rect 50865 7677 51065 7693
rect 50865 7643 50881 7677
rect 51049 7643 51065 7677
rect 50865 7596 51065 7643
rect 39333 7149 39533 7196
rect 39333 7115 39349 7149
rect 39517 7115 39533 7149
rect 39333 7099 39533 7115
rect 39705 7149 39905 7196
rect 39705 7115 39721 7149
rect 39889 7115 39905 7149
rect 39705 7099 39905 7115
rect 40077 7149 40277 7196
rect 40077 7115 40093 7149
rect 40261 7115 40277 7149
rect 40077 7099 40277 7115
rect 40449 7149 40649 7196
rect 40449 7115 40465 7149
rect 40633 7115 40649 7149
rect 40449 7099 40649 7115
rect 40821 7149 41021 7196
rect 40821 7115 40837 7149
rect 41005 7115 41021 7149
rect 40821 7099 41021 7115
rect 41193 7149 41393 7196
rect 41193 7115 41209 7149
rect 41377 7115 41393 7149
rect 41193 7099 41393 7115
rect 41565 7149 41765 7196
rect 41565 7115 41581 7149
rect 41749 7115 41765 7149
rect 41565 7099 41765 7115
rect 41937 7149 42137 7196
rect 41937 7115 41953 7149
rect 42121 7115 42137 7149
rect 41937 7099 42137 7115
rect 42309 7149 42509 7196
rect 42309 7115 42325 7149
rect 42493 7115 42509 7149
rect 42309 7099 42509 7115
rect 42681 7149 42881 7196
rect 42681 7115 42697 7149
rect 42865 7115 42881 7149
rect 42681 7099 42881 7115
rect 43053 7149 43253 7196
rect 43053 7115 43069 7149
rect 43237 7115 43253 7149
rect 43053 7099 43253 7115
rect 43425 7149 43625 7196
rect 43425 7115 43441 7149
rect 43609 7115 43625 7149
rect 43425 7099 43625 7115
rect 43797 7149 43997 7196
rect 43797 7115 43813 7149
rect 43981 7115 43997 7149
rect 43797 7099 43997 7115
rect 44169 7149 44369 7196
rect 44169 7115 44185 7149
rect 44353 7115 44369 7149
rect 44169 7099 44369 7115
rect 44541 7149 44741 7196
rect 44541 7115 44557 7149
rect 44725 7115 44741 7149
rect 44541 7099 44741 7115
rect 44913 7149 45113 7196
rect 44913 7115 44929 7149
rect 45097 7115 45113 7149
rect 44913 7099 45113 7115
rect 45285 7149 45485 7196
rect 45285 7115 45301 7149
rect 45469 7115 45485 7149
rect 45285 7099 45485 7115
rect 45657 7149 45857 7196
rect 45657 7115 45673 7149
rect 45841 7115 45857 7149
rect 45657 7099 45857 7115
rect 46029 7149 46229 7196
rect 46029 7115 46045 7149
rect 46213 7115 46229 7149
rect 46029 7099 46229 7115
rect 46401 7149 46601 7196
rect 46401 7115 46417 7149
rect 46585 7115 46601 7149
rect 46401 7099 46601 7115
rect 46773 7149 46973 7196
rect 46773 7115 46789 7149
rect 46957 7115 46973 7149
rect 46773 7099 46973 7115
rect 47145 7149 47345 7196
rect 47145 7115 47161 7149
rect 47329 7115 47345 7149
rect 47145 7099 47345 7115
rect 47517 7149 47717 7196
rect 47517 7115 47533 7149
rect 47701 7115 47717 7149
rect 47517 7099 47717 7115
rect 47889 7149 48089 7196
rect 47889 7115 47905 7149
rect 48073 7115 48089 7149
rect 47889 7099 48089 7115
rect 48261 7149 48461 7196
rect 48261 7115 48277 7149
rect 48445 7115 48461 7149
rect 48261 7099 48461 7115
rect 48633 7149 48833 7196
rect 48633 7115 48649 7149
rect 48817 7115 48833 7149
rect 48633 7099 48833 7115
rect 49005 7149 49205 7196
rect 49005 7115 49021 7149
rect 49189 7115 49205 7149
rect 49005 7099 49205 7115
rect 49377 7149 49577 7196
rect 49377 7115 49393 7149
rect 49561 7115 49577 7149
rect 49377 7099 49577 7115
rect 49749 7149 49949 7196
rect 49749 7115 49765 7149
rect 49933 7115 49949 7149
rect 49749 7099 49949 7115
rect 50121 7149 50321 7196
rect 50121 7115 50137 7149
rect 50305 7115 50321 7149
rect 50121 7099 50321 7115
rect 50493 7149 50693 7196
rect 50493 7115 50509 7149
rect 50677 7115 50693 7149
rect 50493 7099 50693 7115
rect 50865 7149 51065 7196
rect 50865 7115 50881 7149
rect 51049 7115 51065 7149
rect 50865 7099 51065 7115
rect 40821 6561 41021 6577
rect 40821 6527 40837 6561
rect 41005 6527 41021 6561
rect 40821 6480 41021 6527
rect 41193 6561 41393 6577
rect 41193 6527 41209 6561
rect 41377 6527 41393 6561
rect 41193 6480 41393 6527
rect 41565 6561 41765 6577
rect 41565 6527 41581 6561
rect 41749 6527 41765 6561
rect 41565 6480 41765 6527
rect 41937 6561 42137 6577
rect 41937 6527 41953 6561
rect 42121 6527 42137 6561
rect 41937 6480 42137 6527
rect 42309 6561 42509 6577
rect 42309 6527 42325 6561
rect 42493 6527 42509 6561
rect 42309 6480 42509 6527
rect 42681 6561 42881 6577
rect 42681 6527 42697 6561
rect 42865 6527 42881 6561
rect 42681 6480 42881 6527
rect 43053 6561 43253 6577
rect 43053 6527 43069 6561
rect 43237 6527 43253 6561
rect 43053 6480 43253 6527
rect 43425 6561 43625 6577
rect 43425 6527 43441 6561
rect 43609 6527 43625 6561
rect 43425 6480 43625 6527
rect 40821 5633 41021 5680
rect 40821 5599 40837 5633
rect 41005 5599 41021 5633
rect 40821 5583 41021 5599
rect 41193 5633 41393 5680
rect 41193 5599 41209 5633
rect 41377 5599 41393 5633
rect 41193 5583 41393 5599
rect 41565 5633 41765 5680
rect 41565 5599 41581 5633
rect 41749 5599 41765 5633
rect 41565 5583 41765 5599
rect 41937 5633 42137 5680
rect 41937 5599 41953 5633
rect 42121 5599 42137 5633
rect 41937 5583 42137 5599
rect 42309 5633 42509 5680
rect 42309 5599 42325 5633
rect 42493 5599 42509 5633
rect 42309 5583 42509 5599
rect 42681 5633 42881 5680
rect 42681 5599 42697 5633
rect 42865 5599 42881 5633
rect 42681 5583 42881 5599
rect 43053 5633 43253 5680
rect 43053 5599 43069 5633
rect 43237 5599 43253 5633
rect 43053 5583 43253 5599
rect 43425 5633 43625 5680
rect 43425 5599 43441 5633
rect 43609 5599 43625 5633
rect 43425 5583 43625 5599
rect 40821 5525 41021 5541
rect 40821 5491 40837 5525
rect 41005 5491 41021 5525
rect 40821 5444 41021 5491
rect 41193 5525 41393 5541
rect 41193 5491 41209 5525
rect 41377 5491 41393 5525
rect 41193 5444 41393 5491
rect 41565 5525 41765 5541
rect 41565 5491 41581 5525
rect 41749 5491 41765 5525
rect 41565 5444 41765 5491
rect 41937 5525 42137 5541
rect 41937 5491 41953 5525
rect 42121 5491 42137 5525
rect 41937 5444 42137 5491
rect 42309 5525 42509 5541
rect 42309 5491 42325 5525
rect 42493 5491 42509 5525
rect 42309 5444 42509 5491
rect 42681 5525 42881 5541
rect 42681 5491 42697 5525
rect 42865 5491 42881 5525
rect 42681 5444 42881 5491
rect 43053 5525 43253 5541
rect 43053 5491 43069 5525
rect 43237 5491 43253 5525
rect 43053 5444 43253 5491
rect 43425 5525 43625 5541
rect 43425 5491 43441 5525
rect 43609 5491 43625 5525
rect 43425 5444 43625 5491
rect 40821 4597 41021 4644
rect 40821 4563 40837 4597
rect 41005 4563 41021 4597
rect 40821 4547 41021 4563
rect 41193 4597 41393 4644
rect 41193 4563 41209 4597
rect 41377 4563 41393 4597
rect 41193 4547 41393 4563
rect 41565 4597 41765 4644
rect 41565 4563 41581 4597
rect 41749 4563 41765 4597
rect 41565 4547 41765 4563
rect 41937 4597 42137 4644
rect 41937 4563 41953 4597
rect 42121 4563 42137 4597
rect 41937 4547 42137 4563
rect 42309 4597 42509 4644
rect 42309 4563 42325 4597
rect 42493 4563 42509 4597
rect 42309 4547 42509 4563
rect 42681 4597 42881 4644
rect 42681 4563 42697 4597
rect 42865 4563 42881 4597
rect 42681 4547 42881 4563
rect 43053 4597 43253 4644
rect 43053 4563 43069 4597
rect 43237 4563 43253 4597
rect 43053 4547 43253 4563
rect 43425 4597 43625 4644
rect 43425 4563 43441 4597
rect 43609 4563 43625 4597
rect 43425 4547 43625 4563
rect 40821 4489 41021 4505
rect 40821 4455 40837 4489
rect 41005 4455 41021 4489
rect 40821 4408 41021 4455
rect 41193 4489 41393 4505
rect 41193 4455 41209 4489
rect 41377 4455 41393 4489
rect 41193 4408 41393 4455
rect 41565 4489 41765 4505
rect 41565 4455 41581 4489
rect 41749 4455 41765 4489
rect 41565 4408 41765 4455
rect 41937 4489 42137 4505
rect 41937 4455 41953 4489
rect 42121 4455 42137 4489
rect 41937 4408 42137 4455
rect 42309 4489 42509 4505
rect 42309 4455 42325 4489
rect 42493 4455 42509 4489
rect 42309 4408 42509 4455
rect 42681 4489 42881 4505
rect 42681 4455 42697 4489
rect 42865 4455 42881 4489
rect 42681 4408 42881 4455
rect 43053 4489 43253 4505
rect 43053 4455 43069 4489
rect 43237 4455 43253 4489
rect 43053 4408 43253 4455
rect 43425 4489 43625 4505
rect 43425 4455 43441 4489
rect 43609 4455 43625 4489
rect 43425 4408 43625 4455
rect 40821 3561 41021 3608
rect 40821 3527 40837 3561
rect 41005 3527 41021 3561
rect 40821 3511 41021 3527
rect 41193 3561 41393 3608
rect 41193 3527 41209 3561
rect 41377 3527 41393 3561
rect 41193 3511 41393 3527
rect 41565 3561 41765 3608
rect 41565 3527 41581 3561
rect 41749 3527 41765 3561
rect 41565 3511 41765 3527
rect 41937 3561 42137 3608
rect 41937 3527 41953 3561
rect 42121 3527 42137 3561
rect 41937 3511 42137 3527
rect 42309 3561 42509 3608
rect 42309 3527 42325 3561
rect 42493 3527 42509 3561
rect 42309 3511 42509 3527
rect 42681 3561 42881 3608
rect 42681 3527 42697 3561
rect 42865 3527 42881 3561
rect 42681 3511 42881 3527
rect 43053 3561 43253 3608
rect 43053 3527 43069 3561
rect 43237 3527 43253 3561
rect 43053 3511 43253 3527
rect 43425 3561 43625 3608
rect 43425 3527 43441 3561
rect 43609 3527 43625 3561
rect 43425 3511 43625 3527
rect 40821 3453 41021 3469
rect 40821 3419 40837 3453
rect 41005 3419 41021 3453
rect 40821 3372 41021 3419
rect 41193 3453 41393 3469
rect 41193 3419 41209 3453
rect 41377 3419 41393 3453
rect 41193 3372 41393 3419
rect 41565 3453 41765 3469
rect 41565 3419 41581 3453
rect 41749 3419 41765 3453
rect 41565 3372 41765 3419
rect 41937 3453 42137 3469
rect 41937 3419 41953 3453
rect 42121 3419 42137 3453
rect 41937 3372 42137 3419
rect 42309 3453 42509 3469
rect 42309 3419 42325 3453
rect 42493 3419 42509 3453
rect 42309 3372 42509 3419
rect 42681 3453 42881 3469
rect 42681 3419 42697 3453
rect 42865 3419 42881 3453
rect 42681 3372 42881 3419
rect 43053 3453 43253 3469
rect 43053 3419 43069 3453
rect 43237 3419 43253 3453
rect 43053 3372 43253 3419
rect 43425 3453 43625 3469
rect 43425 3419 43441 3453
rect 43609 3419 43625 3453
rect 43425 3372 43625 3419
rect 40821 2525 41021 2572
rect 40821 2491 40837 2525
rect 41005 2491 41021 2525
rect 40821 2475 41021 2491
rect 41193 2525 41393 2572
rect 41193 2491 41209 2525
rect 41377 2491 41393 2525
rect 41193 2475 41393 2491
rect 41565 2525 41765 2572
rect 41565 2491 41581 2525
rect 41749 2491 41765 2525
rect 41565 2475 41765 2491
rect 41937 2525 42137 2572
rect 41937 2491 41953 2525
rect 42121 2491 42137 2525
rect 41937 2475 42137 2491
rect 42309 2525 42509 2572
rect 42309 2491 42325 2525
rect 42493 2491 42509 2525
rect 42309 2475 42509 2491
rect 42681 2525 42881 2572
rect 42681 2491 42697 2525
rect 42865 2491 42881 2525
rect 42681 2475 42881 2491
rect 43053 2525 43253 2572
rect 43053 2491 43069 2525
rect 43237 2491 43253 2525
rect 43053 2475 43253 2491
rect 43425 2525 43625 2572
rect 43425 2491 43441 2525
rect 43609 2491 43625 2525
rect 43425 2475 43625 2491
rect 40821 1867 41021 1883
rect 40821 1833 40837 1867
rect 41005 1833 41021 1867
rect 40821 1795 41021 1833
rect 41193 1867 41393 1883
rect 41193 1833 41209 1867
rect 41377 1833 41393 1867
rect 41193 1795 41393 1833
rect 41565 1867 41765 1883
rect 41565 1833 41581 1867
rect 41749 1833 41765 1867
rect 41565 1795 41765 1833
rect 41937 1867 42137 1883
rect 41937 1833 41953 1867
rect 42121 1833 42137 1867
rect 41937 1795 42137 1833
rect 42309 1867 42509 1883
rect 42309 1833 42325 1867
rect 42493 1833 42509 1867
rect 42309 1795 42509 1833
rect 42681 1867 42881 1883
rect 42681 1833 42697 1867
rect 42865 1833 42881 1867
rect 42681 1795 42881 1833
rect 43053 1867 43253 1883
rect 43053 1833 43069 1867
rect 43237 1833 43253 1867
rect 43053 1795 43253 1833
rect 43425 1867 43625 1883
rect 43425 1833 43441 1867
rect 43609 1833 43625 1867
rect 43425 1795 43625 1833
rect 43797 1867 43997 1883
rect 43797 1833 43813 1867
rect 43981 1833 43997 1867
rect 43797 1795 43997 1833
rect 44169 1867 44369 1883
rect 44169 1833 44185 1867
rect 44353 1833 44369 1867
rect 44169 1795 44369 1833
rect 44541 1867 44741 1883
rect 44541 1833 44557 1867
rect 44725 1833 44741 1867
rect 44541 1795 44741 1833
rect 44913 1867 45113 1883
rect 44913 1833 44929 1867
rect 45097 1833 45113 1867
rect 44913 1795 45113 1833
rect 45285 1867 45485 1883
rect 45285 1833 45301 1867
rect 45469 1833 45485 1867
rect 45285 1795 45485 1833
rect 45657 1867 45857 1883
rect 45657 1833 45673 1867
rect 45841 1833 45857 1867
rect 45657 1795 45857 1833
rect 46029 1867 46229 1883
rect 46029 1833 46045 1867
rect 46213 1833 46229 1867
rect 46029 1795 46229 1833
rect 46401 1867 46601 1883
rect 46401 1833 46417 1867
rect 46585 1833 46601 1867
rect 46401 1795 46601 1833
rect 46773 1867 46973 1883
rect 46773 1833 46789 1867
rect 46957 1833 46973 1867
rect 46773 1795 46973 1833
rect 47145 1867 47345 1883
rect 47145 1833 47161 1867
rect 47329 1833 47345 1867
rect 47145 1795 47345 1833
rect 47517 1867 47717 1883
rect 47517 1833 47533 1867
rect 47701 1833 47717 1867
rect 47517 1795 47717 1833
rect 47889 1867 48089 1883
rect 47889 1833 47905 1867
rect 48073 1833 48089 1867
rect 47889 1795 48089 1833
rect 48261 1867 48461 1883
rect 48261 1833 48277 1867
rect 48445 1833 48461 1867
rect 48261 1795 48461 1833
rect 48633 1867 48833 1883
rect 48633 1833 48649 1867
rect 48817 1833 48833 1867
rect 48633 1795 48833 1833
rect 49005 1867 49205 1883
rect 49005 1833 49021 1867
rect 49189 1833 49205 1867
rect 49005 1795 49205 1833
rect 49377 1867 49577 1883
rect 49377 1833 49393 1867
rect 49561 1833 49577 1867
rect 49377 1795 49577 1833
rect 40821 1557 41021 1595
rect 40821 1523 40837 1557
rect 41005 1523 41021 1557
rect 40821 1507 41021 1523
rect 41193 1557 41393 1595
rect 41193 1523 41209 1557
rect 41377 1523 41393 1557
rect 41193 1507 41393 1523
rect 41565 1557 41765 1595
rect 41565 1523 41581 1557
rect 41749 1523 41765 1557
rect 41565 1507 41765 1523
rect 41937 1557 42137 1595
rect 41937 1523 41953 1557
rect 42121 1523 42137 1557
rect 41937 1507 42137 1523
rect 42309 1557 42509 1595
rect 42309 1523 42325 1557
rect 42493 1523 42509 1557
rect 42309 1507 42509 1523
rect 42681 1557 42881 1595
rect 42681 1523 42697 1557
rect 42865 1523 42881 1557
rect 42681 1507 42881 1523
rect 43053 1557 43253 1595
rect 43053 1523 43069 1557
rect 43237 1523 43253 1557
rect 43053 1507 43253 1523
rect 43425 1557 43625 1595
rect 43425 1523 43441 1557
rect 43609 1523 43625 1557
rect 43425 1507 43625 1523
rect 43797 1557 43997 1595
rect 43797 1523 43813 1557
rect 43981 1523 43997 1557
rect 43797 1507 43997 1523
rect 44169 1557 44369 1595
rect 44169 1523 44185 1557
rect 44353 1523 44369 1557
rect 44169 1507 44369 1523
rect 44541 1557 44741 1595
rect 44541 1523 44557 1557
rect 44725 1523 44741 1557
rect 44541 1507 44741 1523
rect 44913 1557 45113 1595
rect 44913 1523 44929 1557
rect 45097 1523 45113 1557
rect 44913 1507 45113 1523
rect 45285 1557 45485 1595
rect 45285 1523 45301 1557
rect 45469 1523 45485 1557
rect 45285 1507 45485 1523
rect 45657 1557 45857 1595
rect 45657 1523 45673 1557
rect 45841 1523 45857 1557
rect 45657 1507 45857 1523
rect 46029 1557 46229 1595
rect 46029 1523 46045 1557
rect 46213 1523 46229 1557
rect 46029 1507 46229 1523
rect 46401 1557 46601 1595
rect 46401 1523 46417 1557
rect 46585 1523 46601 1557
rect 46401 1507 46601 1523
rect 46773 1557 46973 1595
rect 46773 1523 46789 1557
rect 46957 1523 46973 1557
rect 46773 1507 46973 1523
rect 47145 1557 47345 1595
rect 47145 1523 47161 1557
rect 47329 1523 47345 1557
rect 47145 1507 47345 1523
rect 47517 1557 47717 1595
rect 47517 1523 47533 1557
rect 47701 1523 47717 1557
rect 47517 1507 47717 1523
rect 47889 1557 48089 1595
rect 47889 1523 47905 1557
rect 48073 1523 48089 1557
rect 47889 1507 48089 1523
rect 48261 1557 48461 1595
rect 48261 1523 48277 1557
rect 48445 1523 48461 1557
rect 48261 1507 48461 1523
rect 48633 1557 48833 1595
rect 48633 1523 48649 1557
rect 48817 1523 48833 1557
rect 48633 1507 48833 1523
rect 49005 1557 49205 1595
rect 49005 1523 49021 1557
rect 49189 1523 49205 1557
rect 49005 1507 49205 1523
rect 49377 1557 49577 1595
rect 49377 1523 49393 1557
rect 49561 1523 49577 1557
rect 49377 1507 49577 1523
rect 40821 1449 41021 1465
rect 40821 1415 40837 1449
rect 41005 1415 41021 1449
rect 40821 1377 41021 1415
rect 41193 1449 41393 1465
rect 41193 1415 41209 1449
rect 41377 1415 41393 1449
rect 41193 1377 41393 1415
rect 41565 1449 41765 1465
rect 41565 1415 41581 1449
rect 41749 1415 41765 1449
rect 41565 1377 41765 1415
rect 41937 1449 42137 1465
rect 41937 1415 41953 1449
rect 42121 1415 42137 1449
rect 41937 1377 42137 1415
rect 42309 1449 42509 1465
rect 42309 1415 42325 1449
rect 42493 1415 42509 1449
rect 42309 1377 42509 1415
rect 42681 1449 42881 1465
rect 42681 1415 42697 1449
rect 42865 1415 42881 1449
rect 42681 1377 42881 1415
rect 43053 1449 43253 1465
rect 43053 1415 43069 1449
rect 43237 1415 43253 1449
rect 43053 1377 43253 1415
rect 43425 1449 43625 1465
rect 43425 1415 43441 1449
rect 43609 1415 43625 1449
rect 43425 1377 43625 1415
rect 43797 1449 43997 1465
rect 43797 1415 43813 1449
rect 43981 1415 43997 1449
rect 43797 1377 43997 1415
rect 44169 1449 44369 1465
rect 44169 1415 44185 1449
rect 44353 1415 44369 1449
rect 44169 1377 44369 1415
rect 44541 1449 44741 1465
rect 44541 1415 44557 1449
rect 44725 1415 44741 1449
rect 44541 1377 44741 1415
rect 44913 1449 45113 1465
rect 44913 1415 44929 1449
rect 45097 1415 45113 1449
rect 44913 1377 45113 1415
rect 45285 1449 45485 1465
rect 45285 1415 45301 1449
rect 45469 1415 45485 1449
rect 45285 1377 45485 1415
rect 45657 1449 45857 1465
rect 45657 1415 45673 1449
rect 45841 1415 45857 1449
rect 45657 1377 45857 1415
rect 46029 1449 46229 1465
rect 46029 1415 46045 1449
rect 46213 1415 46229 1449
rect 46029 1377 46229 1415
rect 46401 1449 46601 1465
rect 46401 1415 46417 1449
rect 46585 1415 46601 1449
rect 46401 1377 46601 1415
rect 46773 1449 46973 1465
rect 46773 1415 46789 1449
rect 46957 1415 46973 1449
rect 46773 1377 46973 1415
rect 47145 1449 47345 1465
rect 47145 1415 47161 1449
rect 47329 1415 47345 1449
rect 47145 1377 47345 1415
rect 47517 1449 47717 1465
rect 47517 1415 47533 1449
rect 47701 1415 47717 1449
rect 47517 1377 47717 1415
rect 47889 1449 48089 1465
rect 47889 1415 47905 1449
rect 48073 1415 48089 1449
rect 47889 1377 48089 1415
rect 48261 1449 48461 1465
rect 48261 1415 48277 1449
rect 48445 1415 48461 1449
rect 48261 1377 48461 1415
rect 48633 1449 48833 1465
rect 48633 1415 48649 1449
rect 48817 1415 48833 1449
rect 48633 1377 48833 1415
rect 49005 1449 49205 1465
rect 49005 1415 49021 1449
rect 49189 1415 49205 1449
rect 49005 1377 49205 1415
rect 49377 1449 49577 1465
rect 49377 1415 49393 1449
rect 49561 1415 49577 1449
rect 49377 1377 49577 1415
rect 40821 1139 41021 1177
rect 40821 1105 40837 1139
rect 41005 1105 41021 1139
rect 40821 1089 41021 1105
rect 41193 1139 41393 1177
rect 41193 1105 41209 1139
rect 41377 1105 41393 1139
rect 41193 1089 41393 1105
rect 41565 1139 41765 1177
rect 41565 1105 41581 1139
rect 41749 1105 41765 1139
rect 41565 1089 41765 1105
rect 41937 1139 42137 1177
rect 41937 1105 41953 1139
rect 42121 1105 42137 1139
rect 41937 1089 42137 1105
rect 42309 1139 42509 1177
rect 42309 1105 42325 1139
rect 42493 1105 42509 1139
rect 42309 1089 42509 1105
rect 42681 1139 42881 1177
rect 42681 1105 42697 1139
rect 42865 1105 42881 1139
rect 42681 1089 42881 1105
rect 43053 1139 43253 1177
rect 43053 1105 43069 1139
rect 43237 1105 43253 1139
rect 43053 1089 43253 1105
rect 43425 1139 43625 1177
rect 43425 1105 43441 1139
rect 43609 1105 43625 1139
rect 43425 1089 43625 1105
rect 43797 1139 43997 1177
rect 43797 1105 43813 1139
rect 43981 1105 43997 1139
rect 43797 1089 43997 1105
rect 44169 1139 44369 1177
rect 44169 1105 44185 1139
rect 44353 1105 44369 1139
rect 44169 1089 44369 1105
rect 44541 1139 44741 1177
rect 44541 1105 44557 1139
rect 44725 1105 44741 1139
rect 44541 1089 44741 1105
rect 44913 1139 45113 1177
rect 44913 1105 44929 1139
rect 45097 1105 45113 1139
rect 44913 1089 45113 1105
rect 45285 1139 45485 1177
rect 45285 1105 45301 1139
rect 45469 1105 45485 1139
rect 45285 1089 45485 1105
rect 45657 1139 45857 1177
rect 45657 1105 45673 1139
rect 45841 1105 45857 1139
rect 45657 1089 45857 1105
rect 46029 1139 46229 1177
rect 46029 1105 46045 1139
rect 46213 1105 46229 1139
rect 46029 1089 46229 1105
rect 46401 1139 46601 1177
rect 46401 1105 46417 1139
rect 46585 1105 46601 1139
rect 46401 1089 46601 1105
rect 46773 1139 46973 1177
rect 46773 1105 46789 1139
rect 46957 1105 46973 1139
rect 46773 1089 46973 1105
rect 47145 1139 47345 1177
rect 47145 1105 47161 1139
rect 47329 1105 47345 1139
rect 47145 1089 47345 1105
rect 47517 1139 47717 1177
rect 47517 1105 47533 1139
rect 47701 1105 47717 1139
rect 47517 1089 47717 1105
rect 47889 1139 48089 1177
rect 47889 1105 47905 1139
rect 48073 1105 48089 1139
rect 47889 1089 48089 1105
rect 48261 1139 48461 1177
rect 48261 1105 48277 1139
rect 48445 1105 48461 1139
rect 48261 1089 48461 1105
rect 48633 1139 48833 1177
rect 48633 1105 48649 1139
rect 48817 1105 48833 1139
rect 48633 1089 48833 1105
rect 49005 1139 49205 1177
rect 49005 1105 49021 1139
rect 49189 1105 49205 1139
rect 49005 1089 49205 1105
rect 49377 1139 49577 1177
rect 49377 1105 49393 1139
rect 49561 1105 49577 1139
rect 49377 1089 49577 1105
rect 40821 1031 41021 1047
rect 40821 997 40837 1031
rect 41005 997 41021 1031
rect 40821 959 41021 997
rect 41193 1031 41393 1047
rect 41193 997 41209 1031
rect 41377 997 41393 1031
rect 41193 959 41393 997
rect 41565 1031 41765 1047
rect 41565 997 41581 1031
rect 41749 997 41765 1031
rect 41565 959 41765 997
rect 41937 1031 42137 1047
rect 41937 997 41953 1031
rect 42121 997 42137 1031
rect 41937 959 42137 997
rect 42309 1031 42509 1047
rect 42309 997 42325 1031
rect 42493 997 42509 1031
rect 42309 959 42509 997
rect 42681 1031 42881 1047
rect 42681 997 42697 1031
rect 42865 997 42881 1031
rect 42681 959 42881 997
rect 43053 1031 43253 1047
rect 43053 997 43069 1031
rect 43237 997 43253 1031
rect 43053 959 43253 997
rect 43425 1031 43625 1047
rect 43425 997 43441 1031
rect 43609 997 43625 1031
rect 43425 959 43625 997
rect 43797 1031 43997 1047
rect 43797 997 43813 1031
rect 43981 997 43997 1031
rect 43797 959 43997 997
rect 44169 1031 44369 1047
rect 44169 997 44185 1031
rect 44353 997 44369 1031
rect 44169 959 44369 997
rect 44541 1031 44741 1047
rect 44541 997 44557 1031
rect 44725 997 44741 1031
rect 44541 959 44741 997
rect 44913 1031 45113 1047
rect 44913 997 44929 1031
rect 45097 997 45113 1031
rect 44913 959 45113 997
rect 45285 1031 45485 1047
rect 45285 997 45301 1031
rect 45469 997 45485 1031
rect 45285 959 45485 997
rect 45657 1031 45857 1047
rect 45657 997 45673 1031
rect 45841 997 45857 1031
rect 45657 959 45857 997
rect 46029 1031 46229 1047
rect 46029 997 46045 1031
rect 46213 997 46229 1031
rect 46029 959 46229 997
rect 46401 1031 46601 1047
rect 46401 997 46417 1031
rect 46585 997 46601 1031
rect 46401 959 46601 997
rect 46773 1031 46973 1047
rect 46773 997 46789 1031
rect 46957 997 46973 1031
rect 46773 959 46973 997
rect 47145 1031 47345 1047
rect 47145 997 47161 1031
rect 47329 997 47345 1031
rect 47145 959 47345 997
rect 47517 1031 47717 1047
rect 47517 997 47533 1031
rect 47701 997 47717 1031
rect 47517 959 47717 997
rect 47889 1031 48089 1047
rect 47889 997 47905 1031
rect 48073 997 48089 1031
rect 47889 959 48089 997
rect 48261 1031 48461 1047
rect 48261 997 48277 1031
rect 48445 997 48461 1031
rect 48261 959 48461 997
rect 48633 1031 48833 1047
rect 48633 997 48649 1031
rect 48817 997 48833 1031
rect 48633 959 48833 997
rect 49005 1031 49205 1047
rect 49005 997 49021 1031
rect 49189 997 49205 1031
rect 49005 959 49205 997
rect 49377 1031 49577 1047
rect 49377 997 49393 1031
rect 49561 997 49577 1031
rect 49377 959 49577 997
rect 40821 721 41021 759
rect 40821 687 40837 721
rect 41005 687 41021 721
rect 40821 671 41021 687
rect 41193 721 41393 759
rect 41193 687 41209 721
rect 41377 687 41393 721
rect 41193 671 41393 687
rect 41565 721 41765 759
rect 41565 687 41581 721
rect 41749 687 41765 721
rect 41565 671 41765 687
rect 41937 721 42137 759
rect 41937 687 41953 721
rect 42121 687 42137 721
rect 41937 671 42137 687
rect 42309 721 42509 759
rect 42309 687 42325 721
rect 42493 687 42509 721
rect 42309 671 42509 687
rect 42681 721 42881 759
rect 42681 687 42697 721
rect 42865 687 42881 721
rect 42681 671 42881 687
rect 43053 721 43253 759
rect 43053 687 43069 721
rect 43237 687 43253 721
rect 43053 671 43253 687
rect 43425 721 43625 759
rect 43425 687 43441 721
rect 43609 687 43625 721
rect 43425 671 43625 687
rect 43797 721 43997 759
rect 43797 687 43813 721
rect 43981 687 43997 721
rect 43797 671 43997 687
rect 44169 721 44369 759
rect 44169 687 44185 721
rect 44353 687 44369 721
rect 44169 671 44369 687
rect 44541 721 44741 759
rect 44541 687 44557 721
rect 44725 687 44741 721
rect 44541 671 44741 687
rect 44913 721 45113 759
rect 44913 687 44929 721
rect 45097 687 45113 721
rect 44913 671 45113 687
rect 45285 721 45485 759
rect 45285 687 45301 721
rect 45469 687 45485 721
rect 45285 671 45485 687
rect 45657 721 45857 759
rect 45657 687 45673 721
rect 45841 687 45857 721
rect 45657 671 45857 687
rect 46029 721 46229 759
rect 46029 687 46045 721
rect 46213 687 46229 721
rect 46029 671 46229 687
rect 46401 721 46601 759
rect 46401 687 46417 721
rect 46585 687 46601 721
rect 46401 671 46601 687
rect 46773 721 46973 759
rect 46773 687 46789 721
rect 46957 687 46973 721
rect 46773 671 46973 687
rect 47145 721 47345 759
rect 47145 687 47161 721
rect 47329 687 47345 721
rect 47145 671 47345 687
rect 47517 721 47717 759
rect 47517 687 47533 721
rect 47701 687 47717 721
rect 47517 671 47717 687
rect 47889 721 48089 759
rect 47889 687 47905 721
rect 48073 687 48089 721
rect 47889 671 48089 687
rect 48261 721 48461 759
rect 48261 687 48277 721
rect 48445 687 48461 721
rect 48261 671 48461 687
rect 48633 721 48833 759
rect 48633 687 48649 721
rect 48817 687 48833 721
rect 48633 671 48833 687
rect 49005 721 49205 759
rect 49005 687 49021 721
rect 49189 687 49205 721
rect 49005 671 49205 687
rect 49377 721 49577 759
rect 49377 687 49393 721
rect 49561 687 49577 721
rect 49377 671 49577 687
rect 40821 613 41021 629
rect 40821 579 40837 613
rect 41005 579 41021 613
rect 40821 541 41021 579
rect 41193 613 41393 629
rect 41193 579 41209 613
rect 41377 579 41393 613
rect 41193 541 41393 579
rect 41565 613 41765 629
rect 41565 579 41581 613
rect 41749 579 41765 613
rect 41565 541 41765 579
rect 41937 613 42137 629
rect 41937 579 41953 613
rect 42121 579 42137 613
rect 41937 541 42137 579
rect 42309 613 42509 629
rect 42309 579 42325 613
rect 42493 579 42509 613
rect 42309 541 42509 579
rect 42681 613 42881 629
rect 42681 579 42697 613
rect 42865 579 42881 613
rect 42681 541 42881 579
rect 43053 613 43253 629
rect 43053 579 43069 613
rect 43237 579 43253 613
rect 43053 541 43253 579
rect 43425 613 43625 629
rect 43425 579 43441 613
rect 43609 579 43625 613
rect 43425 541 43625 579
rect 43797 613 43997 629
rect 43797 579 43813 613
rect 43981 579 43997 613
rect 43797 541 43997 579
rect 44169 613 44369 629
rect 44169 579 44185 613
rect 44353 579 44369 613
rect 44169 541 44369 579
rect 44541 613 44741 629
rect 44541 579 44557 613
rect 44725 579 44741 613
rect 44541 541 44741 579
rect 44913 613 45113 629
rect 44913 579 44929 613
rect 45097 579 45113 613
rect 44913 541 45113 579
rect 45285 613 45485 629
rect 45285 579 45301 613
rect 45469 579 45485 613
rect 45285 541 45485 579
rect 45657 613 45857 629
rect 45657 579 45673 613
rect 45841 579 45857 613
rect 45657 541 45857 579
rect 46029 613 46229 629
rect 46029 579 46045 613
rect 46213 579 46229 613
rect 46029 541 46229 579
rect 46401 613 46601 629
rect 46401 579 46417 613
rect 46585 579 46601 613
rect 46401 541 46601 579
rect 46773 613 46973 629
rect 46773 579 46789 613
rect 46957 579 46973 613
rect 46773 541 46973 579
rect 47145 613 47345 629
rect 47145 579 47161 613
rect 47329 579 47345 613
rect 47145 541 47345 579
rect 47517 613 47717 629
rect 47517 579 47533 613
rect 47701 579 47717 613
rect 47517 541 47717 579
rect 47889 613 48089 629
rect 47889 579 47905 613
rect 48073 579 48089 613
rect 47889 541 48089 579
rect 48261 613 48461 629
rect 48261 579 48277 613
rect 48445 579 48461 613
rect 48261 541 48461 579
rect 48633 613 48833 629
rect 48633 579 48649 613
rect 48817 579 48833 613
rect 48633 541 48833 579
rect 49005 613 49205 629
rect 49005 579 49021 613
rect 49189 579 49205 613
rect 49005 541 49205 579
rect 49377 613 49577 629
rect 49377 579 49393 613
rect 49561 579 49577 613
rect 49377 541 49577 579
rect 40821 303 41021 341
rect 40821 269 40837 303
rect 41005 269 41021 303
rect 40821 253 41021 269
rect 41193 303 41393 341
rect 41193 269 41209 303
rect 41377 269 41393 303
rect 41193 253 41393 269
rect 41565 303 41765 341
rect 41565 269 41581 303
rect 41749 269 41765 303
rect 41565 253 41765 269
rect 41937 303 42137 341
rect 41937 269 41953 303
rect 42121 269 42137 303
rect 41937 253 42137 269
rect 42309 303 42509 341
rect 42309 269 42325 303
rect 42493 269 42509 303
rect 42309 253 42509 269
rect 42681 303 42881 341
rect 42681 269 42697 303
rect 42865 269 42881 303
rect 42681 253 42881 269
rect 43053 303 43253 341
rect 43053 269 43069 303
rect 43237 269 43253 303
rect 43053 253 43253 269
rect 43425 303 43625 341
rect 43425 269 43441 303
rect 43609 269 43625 303
rect 43425 253 43625 269
rect 43797 303 43997 341
rect 43797 269 43813 303
rect 43981 269 43997 303
rect 43797 253 43997 269
rect 44169 303 44369 341
rect 44169 269 44185 303
rect 44353 269 44369 303
rect 44169 253 44369 269
rect 44541 303 44741 341
rect 44541 269 44557 303
rect 44725 269 44741 303
rect 44541 253 44741 269
rect 44913 303 45113 341
rect 44913 269 44929 303
rect 45097 269 45113 303
rect 44913 253 45113 269
rect 45285 303 45485 341
rect 45285 269 45301 303
rect 45469 269 45485 303
rect 45285 253 45485 269
rect 45657 303 45857 341
rect 45657 269 45673 303
rect 45841 269 45857 303
rect 45657 253 45857 269
rect 46029 303 46229 341
rect 46029 269 46045 303
rect 46213 269 46229 303
rect 46029 253 46229 269
rect 46401 303 46601 341
rect 46401 269 46417 303
rect 46585 269 46601 303
rect 46401 253 46601 269
rect 46773 303 46973 341
rect 46773 269 46789 303
rect 46957 269 46973 303
rect 46773 253 46973 269
rect 47145 303 47345 341
rect 47145 269 47161 303
rect 47329 269 47345 303
rect 47145 253 47345 269
rect 47517 303 47717 341
rect 47517 269 47533 303
rect 47701 269 47717 303
rect 47517 253 47717 269
rect 47889 303 48089 341
rect 47889 269 47905 303
rect 48073 269 48089 303
rect 47889 253 48089 269
rect 48261 303 48461 341
rect 48261 269 48277 303
rect 48445 269 48461 303
rect 48261 253 48461 269
rect 48633 303 48833 341
rect 48633 269 48649 303
rect 48817 269 48833 303
rect 48633 253 48833 269
rect 49005 303 49205 341
rect 49005 269 49021 303
rect 49189 269 49205 303
rect 49005 253 49205 269
rect 49377 303 49577 341
rect 49377 269 49393 303
rect 49561 269 49577 303
rect 49377 253 49577 269
<< polycont >>
rect 40837 19562 41005 19596
rect 41209 19562 41377 19596
rect 41581 19562 41749 19596
rect 41953 19562 42121 19596
rect 42325 19562 42493 19596
rect 42697 19562 42865 19596
rect 43069 19562 43237 19596
rect 43441 19562 43609 19596
rect 43813 19562 43981 19596
rect 44185 19562 44353 19596
rect 44557 19562 44725 19596
rect 44929 19562 45097 19596
rect 45301 19562 45469 19596
rect 45673 19562 45841 19596
rect 46045 19562 46213 19596
rect 46417 19562 46585 19596
rect 46789 19562 46957 19596
rect 47161 19562 47329 19596
rect 47533 19562 47701 19596
rect 47905 19562 48073 19596
rect 48277 19562 48445 19596
rect 48649 19562 48817 19596
rect 49021 19562 49189 19596
rect 49393 19562 49561 19596
rect 40837 19252 41005 19286
rect 41209 19252 41377 19286
rect 41581 19252 41749 19286
rect 41953 19252 42121 19286
rect 42325 19252 42493 19286
rect 42697 19252 42865 19286
rect 43069 19252 43237 19286
rect 43441 19252 43609 19286
rect 43813 19252 43981 19286
rect 44185 19252 44353 19286
rect 44557 19252 44725 19286
rect 44929 19252 45097 19286
rect 45301 19252 45469 19286
rect 45673 19252 45841 19286
rect 46045 19252 46213 19286
rect 46417 19252 46585 19286
rect 46789 19252 46957 19286
rect 47161 19252 47329 19286
rect 47533 19252 47701 19286
rect 47905 19252 48073 19286
rect 48277 19252 48445 19286
rect 48649 19252 48817 19286
rect 49021 19252 49189 19286
rect 49393 19252 49561 19286
rect 40837 19144 41005 19178
rect 41209 19144 41377 19178
rect 41581 19144 41749 19178
rect 41953 19144 42121 19178
rect 42325 19144 42493 19178
rect 42697 19144 42865 19178
rect 43069 19144 43237 19178
rect 43441 19144 43609 19178
rect 43813 19144 43981 19178
rect 44185 19144 44353 19178
rect 44557 19144 44725 19178
rect 44929 19144 45097 19178
rect 45301 19144 45469 19178
rect 45673 19144 45841 19178
rect 46045 19144 46213 19178
rect 46417 19144 46585 19178
rect 46789 19144 46957 19178
rect 47161 19144 47329 19178
rect 47533 19144 47701 19178
rect 47905 19144 48073 19178
rect 48277 19144 48445 19178
rect 48649 19144 48817 19178
rect 49021 19144 49189 19178
rect 49393 19144 49561 19178
rect 40837 18834 41005 18868
rect 41209 18834 41377 18868
rect 41581 18834 41749 18868
rect 41953 18834 42121 18868
rect 42325 18834 42493 18868
rect 42697 18834 42865 18868
rect 43069 18834 43237 18868
rect 43441 18834 43609 18868
rect 43813 18834 43981 18868
rect 44185 18834 44353 18868
rect 44557 18834 44725 18868
rect 44929 18834 45097 18868
rect 45301 18834 45469 18868
rect 45673 18834 45841 18868
rect 46045 18834 46213 18868
rect 46417 18834 46585 18868
rect 46789 18834 46957 18868
rect 47161 18834 47329 18868
rect 47533 18834 47701 18868
rect 47905 18834 48073 18868
rect 48277 18834 48445 18868
rect 48649 18834 48817 18868
rect 49021 18834 49189 18868
rect 49393 18834 49561 18868
rect 40837 18726 41005 18760
rect 41209 18726 41377 18760
rect 41581 18726 41749 18760
rect 41953 18726 42121 18760
rect 42325 18726 42493 18760
rect 42697 18726 42865 18760
rect 43069 18726 43237 18760
rect 43441 18726 43609 18760
rect 43813 18726 43981 18760
rect 44185 18726 44353 18760
rect 44557 18726 44725 18760
rect 44929 18726 45097 18760
rect 45301 18726 45469 18760
rect 45673 18726 45841 18760
rect 46045 18726 46213 18760
rect 46417 18726 46585 18760
rect 46789 18726 46957 18760
rect 47161 18726 47329 18760
rect 47533 18726 47701 18760
rect 47905 18726 48073 18760
rect 48277 18726 48445 18760
rect 48649 18726 48817 18760
rect 49021 18726 49189 18760
rect 49393 18726 49561 18760
rect 40837 18416 41005 18450
rect 41209 18416 41377 18450
rect 41581 18416 41749 18450
rect 41953 18416 42121 18450
rect 42325 18416 42493 18450
rect 42697 18416 42865 18450
rect 43069 18416 43237 18450
rect 43441 18416 43609 18450
rect 43813 18416 43981 18450
rect 44185 18416 44353 18450
rect 44557 18416 44725 18450
rect 44929 18416 45097 18450
rect 45301 18416 45469 18450
rect 45673 18416 45841 18450
rect 46045 18416 46213 18450
rect 46417 18416 46585 18450
rect 46789 18416 46957 18450
rect 47161 18416 47329 18450
rect 47533 18416 47701 18450
rect 47905 18416 48073 18450
rect 48277 18416 48445 18450
rect 48649 18416 48817 18450
rect 49021 18416 49189 18450
rect 49393 18416 49561 18450
rect 40837 18308 41005 18342
rect 41209 18308 41377 18342
rect 41581 18308 41749 18342
rect 41953 18308 42121 18342
rect 42325 18308 42493 18342
rect 42697 18308 42865 18342
rect 43069 18308 43237 18342
rect 43441 18308 43609 18342
rect 43813 18308 43981 18342
rect 44185 18308 44353 18342
rect 44557 18308 44725 18342
rect 44929 18308 45097 18342
rect 45301 18308 45469 18342
rect 45673 18308 45841 18342
rect 46045 18308 46213 18342
rect 46417 18308 46585 18342
rect 46789 18308 46957 18342
rect 47161 18308 47329 18342
rect 47533 18308 47701 18342
rect 47905 18308 48073 18342
rect 48277 18308 48445 18342
rect 48649 18308 48817 18342
rect 49021 18308 49189 18342
rect 49393 18308 49561 18342
rect 40837 17998 41005 18032
rect 41209 17998 41377 18032
rect 41581 17998 41749 18032
rect 41953 17998 42121 18032
rect 42325 17998 42493 18032
rect 42697 17998 42865 18032
rect 43069 17998 43237 18032
rect 43441 17998 43609 18032
rect 43813 17998 43981 18032
rect 44185 17998 44353 18032
rect 44557 17998 44725 18032
rect 44929 17998 45097 18032
rect 45301 17998 45469 18032
rect 45673 17998 45841 18032
rect 46045 17998 46213 18032
rect 46417 17998 46585 18032
rect 46789 17998 46957 18032
rect 47161 17998 47329 18032
rect 47533 17998 47701 18032
rect 47905 17998 48073 18032
rect 48277 17998 48445 18032
rect 48649 17998 48817 18032
rect 49021 17998 49189 18032
rect 49393 17998 49561 18032
rect 40837 17340 41005 17374
rect 41209 17340 41377 17374
rect 41581 17340 41749 17374
rect 41953 17340 42121 17374
rect 42325 17340 42493 17374
rect 42697 17340 42865 17374
rect 43069 17340 43237 17374
rect 43441 17340 43609 17374
rect 40837 16412 41005 16446
rect 41209 16412 41377 16446
rect 41581 16412 41749 16446
rect 41953 16412 42121 16446
rect 42325 16412 42493 16446
rect 42697 16412 42865 16446
rect 43069 16412 43237 16446
rect 43441 16412 43609 16446
rect 40837 16304 41005 16338
rect 41209 16304 41377 16338
rect 41581 16304 41749 16338
rect 41953 16304 42121 16338
rect 42325 16304 42493 16338
rect 42697 16304 42865 16338
rect 43069 16304 43237 16338
rect 43441 16304 43609 16338
rect 40837 15376 41005 15410
rect 41209 15376 41377 15410
rect 41581 15376 41749 15410
rect 41953 15376 42121 15410
rect 42325 15376 42493 15410
rect 42697 15376 42865 15410
rect 43069 15376 43237 15410
rect 43441 15376 43609 15410
rect 40837 15268 41005 15302
rect 41209 15268 41377 15302
rect 41581 15268 41749 15302
rect 41953 15268 42121 15302
rect 42325 15268 42493 15302
rect 42697 15268 42865 15302
rect 43069 15268 43237 15302
rect 43441 15268 43609 15302
rect 40837 14340 41005 14374
rect 41209 14340 41377 14374
rect 41581 14340 41749 14374
rect 41953 14340 42121 14374
rect 42325 14340 42493 14374
rect 42697 14340 42865 14374
rect 43069 14340 43237 14374
rect 43441 14340 43609 14374
rect 40837 14232 41005 14266
rect 41209 14232 41377 14266
rect 41581 14232 41749 14266
rect 41953 14232 42121 14266
rect 42325 14232 42493 14266
rect 42697 14232 42865 14266
rect 43069 14232 43237 14266
rect 43441 14232 43609 14266
rect 40837 13304 41005 13338
rect 41209 13304 41377 13338
rect 41581 13304 41749 13338
rect 41953 13304 42121 13338
rect 42325 13304 42493 13338
rect 42697 13304 42865 13338
rect 43069 13304 43237 13338
rect 43441 13304 43609 13338
rect 39349 12716 39517 12750
rect 39721 12716 39889 12750
rect 40093 12716 40261 12750
rect 40465 12716 40633 12750
rect 40837 12716 41005 12750
rect 41209 12716 41377 12750
rect 41581 12716 41749 12750
rect 41953 12716 42121 12750
rect 42325 12716 42493 12750
rect 42697 12716 42865 12750
rect 43069 12716 43237 12750
rect 43441 12716 43609 12750
rect 43813 12716 43981 12750
rect 44185 12716 44353 12750
rect 44557 12716 44725 12750
rect 44929 12716 45097 12750
rect 45301 12716 45469 12750
rect 45673 12716 45841 12750
rect 46045 12716 46213 12750
rect 46417 12716 46585 12750
rect 46789 12716 46957 12750
rect 47161 12716 47329 12750
rect 47533 12716 47701 12750
rect 47905 12716 48073 12750
rect 48277 12716 48445 12750
rect 48649 12716 48817 12750
rect 49021 12716 49189 12750
rect 49393 12716 49561 12750
rect 49765 12716 49933 12750
rect 50137 12716 50305 12750
rect 50509 12716 50677 12750
rect 50881 12716 51049 12750
rect 39349 12188 39517 12222
rect 39721 12188 39889 12222
rect 40093 12188 40261 12222
rect 40465 12188 40633 12222
rect 40837 12188 41005 12222
rect 41209 12188 41377 12222
rect 41581 12188 41749 12222
rect 41953 12188 42121 12222
rect 42325 12188 42493 12222
rect 42697 12188 42865 12222
rect 43069 12188 43237 12222
rect 43441 12188 43609 12222
rect 43813 12188 43981 12222
rect 44185 12188 44353 12222
rect 44557 12188 44725 12222
rect 44929 12188 45097 12222
rect 45301 12188 45469 12222
rect 45673 12188 45841 12222
rect 46045 12188 46213 12222
rect 46417 12188 46585 12222
rect 46789 12188 46957 12222
rect 47161 12188 47329 12222
rect 47533 12188 47701 12222
rect 47905 12188 48073 12222
rect 48277 12188 48445 12222
rect 48649 12188 48817 12222
rect 49021 12188 49189 12222
rect 49393 12188 49561 12222
rect 49765 12188 49933 12222
rect 50137 12188 50305 12222
rect 50509 12188 50677 12222
rect 50881 12188 51049 12222
rect 39349 12080 39517 12114
rect 39721 12080 39889 12114
rect 40093 12080 40261 12114
rect 40465 12080 40633 12114
rect 40837 12080 41005 12114
rect 41209 12080 41377 12114
rect 41581 12080 41749 12114
rect 41953 12080 42121 12114
rect 42325 12080 42493 12114
rect 42697 12080 42865 12114
rect 43069 12080 43237 12114
rect 43441 12080 43609 12114
rect 43813 12080 43981 12114
rect 44185 12080 44353 12114
rect 44557 12080 44725 12114
rect 44929 12080 45097 12114
rect 45301 12080 45469 12114
rect 45673 12080 45841 12114
rect 46045 12080 46213 12114
rect 46417 12080 46585 12114
rect 46789 12080 46957 12114
rect 47161 12080 47329 12114
rect 47533 12080 47701 12114
rect 47905 12080 48073 12114
rect 48277 12080 48445 12114
rect 48649 12080 48817 12114
rect 49021 12080 49189 12114
rect 49393 12080 49561 12114
rect 49765 12080 49933 12114
rect 50137 12080 50305 12114
rect 50509 12080 50677 12114
rect 50881 12080 51049 12114
rect 39349 11552 39517 11586
rect 39721 11552 39889 11586
rect 40093 11552 40261 11586
rect 40465 11552 40633 11586
rect 40837 11552 41005 11586
rect 41209 11552 41377 11586
rect 41581 11552 41749 11586
rect 41953 11552 42121 11586
rect 42325 11552 42493 11586
rect 42697 11552 42865 11586
rect 43069 11552 43237 11586
rect 43441 11552 43609 11586
rect 43813 11552 43981 11586
rect 44185 11552 44353 11586
rect 44557 11552 44725 11586
rect 44929 11552 45097 11586
rect 45301 11552 45469 11586
rect 45673 11552 45841 11586
rect 46045 11552 46213 11586
rect 46417 11552 46585 11586
rect 46789 11552 46957 11586
rect 47161 11552 47329 11586
rect 47533 11552 47701 11586
rect 47905 11552 48073 11586
rect 48277 11552 48445 11586
rect 48649 11552 48817 11586
rect 49021 11552 49189 11586
rect 49393 11552 49561 11586
rect 49765 11552 49933 11586
rect 50137 11552 50305 11586
rect 50509 11552 50677 11586
rect 50881 11552 51049 11586
rect 39349 11444 39517 11478
rect 39721 11444 39889 11478
rect 40093 11444 40261 11478
rect 40465 11444 40633 11478
rect 40837 11444 41005 11478
rect 41209 11444 41377 11478
rect 41581 11444 41749 11478
rect 41953 11444 42121 11478
rect 42325 11444 42493 11478
rect 42697 11444 42865 11478
rect 43069 11444 43237 11478
rect 43441 11444 43609 11478
rect 43813 11444 43981 11478
rect 44185 11444 44353 11478
rect 44557 11444 44725 11478
rect 44929 11444 45097 11478
rect 45301 11444 45469 11478
rect 45673 11444 45841 11478
rect 46045 11444 46213 11478
rect 46417 11444 46585 11478
rect 46789 11444 46957 11478
rect 47161 11444 47329 11478
rect 47533 11444 47701 11478
rect 47905 11444 48073 11478
rect 48277 11444 48445 11478
rect 48649 11444 48817 11478
rect 49021 11444 49189 11478
rect 49393 11444 49561 11478
rect 49765 11444 49933 11478
rect 50137 11444 50305 11478
rect 50509 11444 50677 11478
rect 50881 11444 51049 11478
rect 39349 10916 39517 10950
rect 39721 10916 39889 10950
rect 40093 10916 40261 10950
rect 40465 10916 40633 10950
rect 40837 10916 41005 10950
rect 41209 10916 41377 10950
rect 41581 10916 41749 10950
rect 41953 10916 42121 10950
rect 42325 10916 42493 10950
rect 42697 10916 42865 10950
rect 43069 10916 43237 10950
rect 43441 10916 43609 10950
rect 43813 10916 43981 10950
rect 44185 10916 44353 10950
rect 44557 10916 44725 10950
rect 44929 10916 45097 10950
rect 45301 10916 45469 10950
rect 45673 10916 45841 10950
rect 46045 10916 46213 10950
rect 46417 10916 46585 10950
rect 46789 10916 46957 10950
rect 47161 10916 47329 10950
rect 47533 10916 47701 10950
rect 47905 10916 48073 10950
rect 48277 10916 48445 10950
rect 48649 10916 48817 10950
rect 49021 10916 49189 10950
rect 49393 10916 49561 10950
rect 49765 10916 49933 10950
rect 50137 10916 50305 10950
rect 50509 10916 50677 10950
rect 50881 10916 51049 10950
rect 39349 8915 39517 8949
rect 39721 8915 39889 8949
rect 40093 8915 40261 8949
rect 40465 8915 40633 8949
rect 40837 8915 41005 8949
rect 41209 8915 41377 8949
rect 41581 8915 41749 8949
rect 41953 8915 42121 8949
rect 42325 8915 42493 8949
rect 42697 8915 42865 8949
rect 43069 8915 43237 8949
rect 43441 8915 43609 8949
rect 43813 8915 43981 8949
rect 44185 8915 44353 8949
rect 44557 8915 44725 8949
rect 44929 8915 45097 8949
rect 45301 8915 45469 8949
rect 45673 8915 45841 8949
rect 46045 8915 46213 8949
rect 46417 8915 46585 8949
rect 46789 8915 46957 8949
rect 47161 8915 47329 8949
rect 47533 8915 47701 8949
rect 47905 8915 48073 8949
rect 48277 8915 48445 8949
rect 48649 8915 48817 8949
rect 49021 8915 49189 8949
rect 49393 8915 49561 8949
rect 49765 8915 49933 8949
rect 50137 8915 50305 8949
rect 50509 8915 50677 8949
rect 50881 8915 51049 8949
rect 39349 8387 39517 8421
rect 39721 8387 39889 8421
rect 40093 8387 40261 8421
rect 40465 8387 40633 8421
rect 40837 8387 41005 8421
rect 41209 8387 41377 8421
rect 41581 8387 41749 8421
rect 41953 8387 42121 8421
rect 42325 8387 42493 8421
rect 42697 8387 42865 8421
rect 43069 8387 43237 8421
rect 43441 8387 43609 8421
rect 43813 8387 43981 8421
rect 44185 8387 44353 8421
rect 44557 8387 44725 8421
rect 44929 8387 45097 8421
rect 45301 8387 45469 8421
rect 45673 8387 45841 8421
rect 46045 8387 46213 8421
rect 46417 8387 46585 8421
rect 46789 8387 46957 8421
rect 47161 8387 47329 8421
rect 47533 8387 47701 8421
rect 47905 8387 48073 8421
rect 48277 8387 48445 8421
rect 48649 8387 48817 8421
rect 49021 8387 49189 8421
rect 49393 8387 49561 8421
rect 49765 8387 49933 8421
rect 50137 8387 50305 8421
rect 50509 8387 50677 8421
rect 50881 8387 51049 8421
rect 39349 8279 39517 8313
rect 39721 8279 39889 8313
rect 40093 8279 40261 8313
rect 40465 8279 40633 8313
rect 40837 8279 41005 8313
rect 41209 8279 41377 8313
rect 41581 8279 41749 8313
rect 41953 8279 42121 8313
rect 42325 8279 42493 8313
rect 42697 8279 42865 8313
rect 43069 8279 43237 8313
rect 43441 8279 43609 8313
rect 43813 8279 43981 8313
rect 44185 8279 44353 8313
rect 44557 8279 44725 8313
rect 44929 8279 45097 8313
rect 45301 8279 45469 8313
rect 45673 8279 45841 8313
rect 46045 8279 46213 8313
rect 46417 8279 46585 8313
rect 46789 8279 46957 8313
rect 47161 8279 47329 8313
rect 47533 8279 47701 8313
rect 47905 8279 48073 8313
rect 48277 8279 48445 8313
rect 48649 8279 48817 8313
rect 49021 8279 49189 8313
rect 49393 8279 49561 8313
rect 49765 8279 49933 8313
rect 50137 8279 50305 8313
rect 50509 8279 50677 8313
rect 50881 8279 51049 8313
rect 39349 7751 39517 7785
rect 39721 7751 39889 7785
rect 40093 7751 40261 7785
rect 40465 7751 40633 7785
rect 40837 7751 41005 7785
rect 41209 7751 41377 7785
rect 41581 7751 41749 7785
rect 41953 7751 42121 7785
rect 42325 7751 42493 7785
rect 42697 7751 42865 7785
rect 43069 7751 43237 7785
rect 43441 7751 43609 7785
rect 43813 7751 43981 7785
rect 44185 7751 44353 7785
rect 44557 7751 44725 7785
rect 44929 7751 45097 7785
rect 45301 7751 45469 7785
rect 45673 7751 45841 7785
rect 46045 7751 46213 7785
rect 46417 7751 46585 7785
rect 46789 7751 46957 7785
rect 47161 7751 47329 7785
rect 47533 7751 47701 7785
rect 47905 7751 48073 7785
rect 48277 7751 48445 7785
rect 48649 7751 48817 7785
rect 49021 7751 49189 7785
rect 49393 7751 49561 7785
rect 49765 7751 49933 7785
rect 50137 7751 50305 7785
rect 50509 7751 50677 7785
rect 50881 7751 51049 7785
rect 39349 7643 39517 7677
rect 39721 7643 39889 7677
rect 40093 7643 40261 7677
rect 40465 7643 40633 7677
rect 40837 7643 41005 7677
rect 41209 7643 41377 7677
rect 41581 7643 41749 7677
rect 41953 7643 42121 7677
rect 42325 7643 42493 7677
rect 42697 7643 42865 7677
rect 43069 7643 43237 7677
rect 43441 7643 43609 7677
rect 43813 7643 43981 7677
rect 44185 7643 44353 7677
rect 44557 7643 44725 7677
rect 44929 7643 45097 7677
rect 45301 7643 45469 7677
rect 45673 7643 45841 7677
rect 46045 7643 46213 7677
rect 46417 7643 46585 7677
rect 46789 7643 46957 7677
rect 47161 7643 47329 7677
rect 47533 7643 47701 7677
rect 47905 7643 48073 7677
rect 48277 7643 48445 7677
rect 48649 7643 48817 7677
rect 49021 7643 49189 7677
rect 49393 7643 49561 7677
rect 49765 7643 49933 7677
rect 50137 7643 50305 7677
rect 50509 7643 50677 7677
rect 50881 7643 51049 7677
rect 39349 7115 39517 7149
rect 39721 7115 39889 7149
rect 40093 7115 40261 7149
rect 40465 7115 40633 7149
rect 40837 7115 41005 7149
rect 41209 7115 41377 7149
rect 41581 7115 41749 7149
rect 41953 7115 42121 7149
rect 42325 7115 42493 7149
rect 42697 7115 42865 7149
rect 43069 7115 43237 7149
rect 43441 7115 43609 7149
rect 43813 7115 43981 7149
rect 44185 7115 44353 7149
rect 44557 7115 44725 7149
rect 44929 7115 45097 7149
rect 45301 7115 45469 7149
rect 45673 7115 45841 7149
rect 46045 7115 46213 7149
rect 46417 7115 46585 7149
rect 46789 7115 46957 7149
rect 47161 7115 47329 7149
rect 47533 7115 47701 7149
rect 47905 7115 48073 7149
rect 48277 7115 48445 7149
rect 48649 7115 48817 7149
rect 49021 7115 49189 7149
rect 49393 7115 49561 7149
rect 49765 7115 49933 7149
rect 50137 7115 50305 7149
rect 50509 7115 50677 7149
rect 50881 7115 51049 7149
rect 40837 6527 41005 6561
rect 41209 6527 41377 6561
rect 41581 6527 41749 6561
rect 41953 6527 42121 6561
rect 42325 6527 42493 6561
rect 42697 6527 42865 6561
rect 43069 6527 43237 6561
rect 43441 6527 43609 6561
rect 40837 5599 41005 5633
rect 41209 5599 41377 5633
rect 41581 5599 41749 5633
rect 41953 5599 42121 5633
rect 42325 5599 42493 5633
rect 42697 5599 42865 5633
rect 43069 5599 43237 5633
rect 43441 5599 43609 5633
rect 40837 5491 41005 5525
rect 41209 5491 41377 5525
rect 41581 5491 41749 5525
rect 41953 5491 42121 5525
rect 42325 5491 42493 5525
rect 42697 5491 42865 5525
rect 43069 5491 43237 5525
rect 43441 5491 43609 5525
rect 40837 4563 41005 4597
rect 41209 4563 41377 4597
rect 41581 4563 41749 4597
rect 41953 4563 42121 4597
rect 42325 4563 42493 4597
rect 42697 4563 42865 4597
rect 43069 4563 43237 4597
rect 43441 4563 43609 4597
rect 40837 4455 41005 4489
rect 41209 4455 41377 4489
rect 41581 4455 41749 4489
rect 41953 4455 42121 4489
rect 42325 4455 42493 4489
rect 42697 4455 42865 4489
rect 43069 4455 43237 4489
rect 43441 4455 43609 4489
rect 40837 3527 41005 3561
rect 41209 3527 41377 3561
rect 41581 3527 41749 3561
rect 41953 3527 42121 3561
rect 42325 3527 42493 3561
rect 42697 3527 42865 3561
rect 43069 3527 43237 3561
rect 43441 3527 43609 3561
rect 40837 3419 41005 3453
rect 41209 3419 41377 3453
rect 41581 3419 41749 3453
rect 41953 3419 42121 3453
rect 42325 3419 42493 3453
rect 42697 3419 42865 3453
rect 43069 3419 43237 3453
rect 43441 3419 43609 3453
rect 40837 2491 41005 2525
rect 41209 2491 41377 2525
rect 41581 2491 41749 2525
rect 41953 2491 42121 2525
rect 42325 2491 42493 2525
rect 42697 2491 42865 2525
rect 43069 2491 43237 2525
rect 43441 2491 43609 2525
rect 40837 1833 41005 1867
rect 41209 1833 41377 1867
rect 41581 1833 41749 1867
rect 41953 1833 42121 1867
rect 42325 1833 42493 1867
rect 42697 1833 42865 1867
rect 43069 1833 43237 1867
rect 43441 1833 43609 1867
rect 43813 1833 43981 1867
rect 44185 1833 44353 1867
rect 44557 1833 44725 1867
rect 44929 1833 45097 1867
rect 45301 1833 45469 1867
rect 45673 1833 45841 1867
rect 46045 1833 46213 1867
rect 46417 1833 46585 1867
rect 46789 1833 46957 1867
rect 47161 1833 47329 1867
rect 47533 1833 47701 1867
rect 47905 1833 48073 1867
rect 48277 1833 48445 1867
rect 48649 1833 48817 1867
rect 49021 1833 49189 1867
rect 49393 1833 49561 1867
rect 40837 1523 41005 1557
rect 41209 1523 41377 1557
rect 41581 1523 41749 1557
rect 41953 1523 42121 1557
rect 42325 1523 42493 1557
rect 42697 1523 42865 1557
rect 43069 1523 43237 1557
rect 43441 1523 43609 1557
rect 43813 1523 43981 1557
rect 44185 1523 44353 1557
rect 44557 1523 44725 1557
rect 44929 1523 45097 1557
rect 45301 1523 45469 1557
rect 45673 1523 45841 1557
rect 46045 1523 46213 1557
rect 46417 1523 46585 1557
rect 46789 1523 46957 1557
rect 47161 1523 47329 1557
rect 47533 1523 47701 1557
rect 47905 1523 48073 1557
rect 48277 1523 48445 1557
rect 48649 1523 48817 1557
rect 49021 1523 49189 1557
rect 49393 1523 49561 1557
rect 40837 1415 41005 1449
rect 41209 1415 41377 1449
rect 41581 1415 41749 1449
rect 41953 1415 42121 1449
rect 42325 1415 42493 1449
rect 42697 1415 42865 1449
rect 43069 1415 43237 1449
rect 43441 1415 43609 1449
rect 43813 1415 43981 1449
rect 44185 1415 44353 1449
rect 44557 1415 44725 1449
rect 44929 1415 45097 1449
rect 45301 1415 45469 1449
rect 45673 1415 45841 1449
rect 46045 1415 46213 1449
rect 46417 1415 46585 1449
rect 46789 1415 46957 1449
rect 47161 1415 47329 1449
rect 47533 1415 47701 1449
rect 47905 1415 48073 1449
rect 48277 1415 48445 1449
rect 48649 1415 48817 1449
rect 49021 1415 49189 1449
rect 49393 1415 49561 1449
rect 40837 1105 41005 1139
rect 41209 1105 41377 1139
rect 41581 1105 41749 1139
rect 41953 1105 42121 1139
rect 42325 1105 42493 1139
rect 42697 1105 42865 1139
rect 43069 1105 43237 1139
rect 43441 1105 43609 1139
rect 43813 1105 43981 1139
rect 44185 1105 44353 1139
rect 44557 1105 44725 1139
rect 44929 1105 45097 1139
rect 45301 1105 45469 1139
rect 45673 1105 45841 1139
rect 46045 1105 46213 1139
rect 46417 1105 46585 1139
rect 46789 1105 46957 1139
rect 47161 1105 47329 1139
rect 47533 1105 47701 1139
rect 47905 1105 48073 1139
rect 48277 1105 48445 1139
rect 48649 1105 48817 1139
rect 49021 1105 49189 1139
rect 49393 1105 49561 1139
rect 40837 997 41005 1031
rect 41209 997 41377 1031
rect 41581 997 41749 1031
rect 41953 997 42121 1031
rect 42325 997 42493 1031
rect 42697 997 42865 1031
rect 43069 997 43237 1031
rect 43441 997 43609 1031
rect 43813 997 43981 1031
rect 44185 997 44353 1031
rect 44557 997 44725 1031
rect 44929 997 45097 1031
rect 45301 997 45469 1031
rect 45673 997 45841 1031
rect 46045 997 46213 1031
rect 46417 997 46585 1031
rect 46789 997 46957 1031
rect 47161 997 47329 1031
rect 47533 997 47701 1031
rect 47905 997 48073 1031
rect 48277 997 48445 1031
rect 48649 997 48817 1031
rect 49021 997 49189 1031
rect 49393 997 49561 1031
rect 40837 687 41005 721
rect 41209 687 41377 721
rect 41581 687 41749 721
rect 41953 687 42121 721
rect 42325 687 42493 721
rect 42697 687 42865 721
rect 43069 687 43237 721
rect 43441 687 43609 721
rect 43813 687 43981 721
rect 44185 687 44353 721
rect 44557 687 44725 721
rect 44929 687 45097 721
rect 45301 687 45469 721
rect 45673 687 45841 721
rect 46045 687 46213 721
rect 46417 687 46585 721
rect 46789 687 46957 721
rect 47161 687 47329 721
rect 47533 687 47701 721
rect 47905 687 48073 721
rect 48277 687 48445 721
rect 48649 687 48817 721
rect 49021 687 49189 721
rect 49393 687 49561 721
rect 40837 579 41005 613
rect 41209 579 41377 613
rect 41581 579 41749 613
rect 41953 579 42121 613
rect 42325 579 42493 613
rect 42697 579 42865 613
rect 43069 579 43237 613
rect 43441 579 43609 613
rect 43813 579 43981 613
rect 44185 579 44353 613
rect 44557 579 44725 613
rect 44929 579 45097 613
rect 45301 579 45469 613
rect 45673 579 45841 613
rect 46045 579 46213 613
rect 46417 579 46585 613
rect 46789 579 46957 613
rect 47161 579 47329 613
rect 47533 579 47701 613
rect 47905 579 48073 613
rect 48277 579 48445 613
rect 48649 579 48817 613
rect 49021 579 49189 613
rect 49393 579 49561 613
rect 40837 269 41005 303
rect 41209 269 41377 303
rect 41581 269 41749 303
rect 41953 269 42121 303
rect 42325 269 42493 303
rect 42697 269 42865 303
rect 43069 269 43237 303
rect 43441 269 43609 303
rect 43813 269 43981 303
rect 44185 269 44353 303
rect 44557 269 44725 303
rect 44929 269 45097 303
rect 45301 269 45469 303
rect 45673 269 45841 303
rect 46045 269 46213 303
rect 46417 269 46585 303
rect 46789 269 46957 303
rect 47161 269 47329 303
rect 47533 269 47701 303
rect 47905 269 48073 303
rect 48277 269 48445 303
rect 48649 269 48817 303
rect 49021 269 49189 303
rect 49393 269 49561 303
<< xpolycontact >>
rect 45955 16020 46025 16452
rect 45955 15488 46025 15920
rect 39505 6308 39575 6740
rect 39505 4876 39575 5308
rect 39823 6308 39893 6740
rect 39823 4876 39893 5308
rect 44661 5668 44731 6100
rect 44661 4236 44731 4668
rect 44979 5668 45049 6100
rect 44979 4236 45049 4668
rect 45955 3945 46025 4377
rect 45955 3413 46025 3845
<< xpolyres >>
rect 45955 15920 46025 16020
rect 39505 5308 39575 6308
rect 39823 5308 39893 6308
rect 44661 4668 44731 5668
rect 44979 4668 45049 5668
rect 45955 3845 46025 3945
<< locali >>
rect 40661 19664 40757 19698
rect 49641 19664 49737 19698
rect 40661 19602 40695 19664
rect 49703 19602 49737 19664
rect 40821 19562 40837 19596
rect 41005 19562 41021 19596
rect 41193 19562 41209 19596
rect 41377 19562 41393 19596
rect 41565 19562 41581 19596
rect 41749 19562 41765 19596
rect 41937 19562 41953 19596
rect 42121 19562 42137 19596
rect 42309 19562 42325 19596
rect 42493 19562 42509 19596
rect 42681 19562 42697 19596
rect 42865 19562 42881 19596
rect 43053 19562 43069 19596
rect 43237 19562 43253 19596
rect 43425 19562 43441 19596
rect 43609 19562 43625 19596
rect 43797 19562 43813 19596
rect 43981 19562 43997 19596
rect 44169 19562 44185 19596
rect 44353 19562 44369 19596
rect 44541 19562 44557 19596
rect 44725 19562 44741 19596
rect 44913 19562 44929 19596
rect 45097 19562 45113 19596
rect 45285 19562 45301 19596
rect 45469 19562 45485 19596
rect 45657 19562 45673 19596
rect 45841 19562 45857 19596
rect 46029 19562 46045 19596
rect 46213 19562 46229 19596
rect 46401 19562 46417 19596
rect 46585 19562 46601 19596
rect 46773 19562 46789 19596
rect 46957 19562 46973 19596
rect 47145 19562 47161 19596
rect 47329 19562 47345 19596
rect 47517 19562 47533 19596
rect 47701 19562 47717 19596
rect 47889 19562 47905 19596
rect 48073 19562 48089 19596
rect 48261 19562 48277 19596
rect 48445 19562 48461 19596
rect 48633 19562 48649 19596
rect 48817 19562 48833 19596
rect 49005 19562 49021 19596
rect 49189 19562 49205 19596
rect 49377 19562 49393 19596
rect 49561 19562 49577 19596
rect 40775 19512 40809 19528
rect 40775 19320 40809 19336
rect 41033 19512 41067 19528
rect 41033 19320 41067 19336
rect 41147 19512 41181 19528
rect 41147 19320 41181 19336
rect 41405 19512 41439 19528
rect 41405 19320 41439 19336
rect 41519 19512 41553 19528
rect 41519 19320 41553 19336
rect 41777 19512 41811 19528
rect 41777 19320 41811 19336
rect 41891 19512 41925 19528
rect 41891 19320 41925 19336
rect 42149 19512 42183 19528
rect 42149 19320 42183 19336
rect 42263 19512 42297 19528
rect 42263 19320 42297 19336
rect 42521 19512 42555 19528
rect 42521 19320 42555 19336
rect 42635 19512 42669 19528
rect 42635 19320 42669 19336
rect 42893 19512 42927 19528
rect 42893 19320 42927 19336
rect 43007 19512 43041 19528
rect 43007 19320 43041 19336
rect 43265 19512 43299 19528
rect 43265 19320 43299 19336
rect 43379 19512 43413 19528
rect 43379 19320 43413 19336
rect 43637 19512 43671 19528
rect 43637 19320 43671 19336
rect 43751 19512 43785 19528
rect 43751 19320 43785 19336
rect 44009 19512 44043 19528
rect 44009 19320 44043 19336
rect 44123 19512 44157 19528
rect 44123 19320 44157 19336
rect 44381 19512 44415 19528
rect 44381 19320 44415 19336
rect 44495 19512 44529 19528
rect 44495 19320 44529 19336
rect 44753 19512 44787 19528
rect 44753 19320 44787 19336
rect 44867 19512 44901 19528
rect 44867 19320 44901 19336
rect 45125 19512 45159 19528
rect 45125 19320 45159 19336
rect 45239 19512 45273 19528
rect 45239 19320 45273 19336
rect 45497 19512 45531 19528
rect 45497 19320 45531 19336
rect 45611 19512 45645 19528
rect 45611 19320 45645 19336
rect 45869 19512 45903 19528
rect 45869 19320 45903 19336
rect 45983 19512 46017 19528
rect 45983 19320 46017 19336
rect 46241 19512 46275 19528
rect 46241 19320 46275 19336
rect 46355 19512 46389 19528
rect 46355 19320 46389 19336
rect 46613 19512 46647 19528
rect 46613 19320 46647 19336
rect 46727 19512 46761 19528
rect 46727 19320 46761 19336
rect 46985 19512 47019 19528
rect 46985 19320 47019 19336
rect 47099 19512 47133 19528
rect 47099 19320 47133 19336
rect 47357 19512 47391 19528
rect 47357 19320 47391 19336
rect 47471 19512 47505 19528
rect 47471 19320 47505 19336
rect 47729 19512 47763 19528
rect 47729 19320 47763 19336
rect 47843 19512 47877 19528
rect 47843 19320 47877 19336
rect 48101 19512 48135 19528
rect 48101 19320 48135 19336
rect 48215 19512 48249 19528
rect 48215 19320 48249 19336
rect 48473 19512 48507 19528
rect 48473 19320 48507 19336
rect 48587 19512 48621 19528
rect 48587 19320 48621 19336
rect 48845 19512 48879 19528
rect 48845 19320 48879 19336
rect 48959 19512 48993 19528
rect 48959 19320 48993 19336
rect 49217 19512 49251 19528
rect 49217 19320 49251 19336
rect 49331 19512 49365 19528
rect 49331 19320 49365 19336
rect 49589 19512 49623 19528
rect 49589 19320 49623 19336
rect 40821 19252 40837 19286
rect 41005 19252 41021 19286
rect 41193 19252 41209 19286
rect 41377 19252 41393 19286
rect 41565 19252 41581 19286
rect 41749 19252 41765 19286
rect 41937 19252 41953 19286
rect 42121 19252 42137 19286
rect 42309 19252 42325 19286
rect 42493 19252 42509 19286
rect 42681 19252 42697 19286
rect 42865 19252 42881 19286
rect 43053 19252 43069 19286
rect 43237 19252 43253 19286
rect 43425 19252 43441 19286
rect 43609 19252 43625 19286
rect 43797 19252 43813 19286
rect 43981 19252 43997 19286
rect 44169 19252 44185 19286
rect 44353 19252 44369 19286
rect 44541 19252 44557 19286
rect 44725 19252 44741 19286
rect 44913 19252 44929 19286
rect 45097 19252 45113 19286
rect 45285 19252 45301 19286
rect 45469 19252 45485 19286
rect 45657 19252 45673 19286
rect 45841 19252 45857 19286
rect 46029 19252 46045 19286
rect 46213 19252 46229 19286
rect 46401 19252 46417 19286
rect 46585 19252 46601 19286
rect 46773 19252 46789 19286
rect 46957 19252 46973 19286
rect 47145 19252 47161 19286
rect 47329 19252 47345 19286
rect 47517 19252 47533 19286
rect 47701 19252 47717 19286
rect 47889 19252 47905 19286
rect 48073 19252 48089 19286
rect 48261 19252 48277 19286
rect 48445 19252 48461 19286
rect 48633 19252 48649 19286
rect 48817 19252 48833 19286
rect 49005 19252 49021 19286
rect 49189 19252 49205 19286
rect 49377 19252 49393 19286
rect 49561 19252 49577 19286
rect 40821 19144 40837 19178
rect 41005 19144 41021 19178
rect 41193 19144 41209 19178
rect 41377 19144 41393 19178
rect 41565 19144 41581 19178
rect 41749 19144 41765 19178
rect 41937 19144 41953 19178
rect 42121 19144 42137 19178
rect 42309 19144 42325 19178
rect 42493 19144 42509 19178
rect 42681 19144 42697 19178
rect 42865 19144 42881 19178
rect 43053 19144 43069 19178
rect 43237 19144 43253 19178
rect 43425 19144 43441 19178
rect 43609 19144 43625 19178
rect 43797 19144 43813 19178
rect 43981 19144 43997 19178
rect 44169 19144 44185 19178
rect 44353 19144 44369 19178
rect 44541 19144 44557 19178
rect 44725 19144 44741 19178
rect 44913 19144 44929 19178
rect 45097 19144 45113 19178
rect 45285 19144 45301 19178
rect 45469 19144 45485 19178
rect 45657 19144 45673 19178
rect 45841 19144 45857 19178
rect 46029 19144 46045 19178
rect 46213 19144 46229 19178
rect 46401 19144 46417 19178
rect 46585 19144 46601 19178
rect 46773 19144 46789 19178
rect 46957 19144 46973 19178
rect 47145 19144 47161 19178
rect 47329 19144 47345 19178
rect 47517 19144 47533 19178
rect 47701 19144 47717 19178
rect 47889 19144 47905 19178
rect 48073 19144 48089 19178
rect 48261 19144 48277 19178
rect 48445 19144 48461 19178
rect 48633 19144 48649 19178
rect 48817 19144 48833 19178
rect 49005 19144 49021 19178
rect 49189 19144 49205 19178
rect 49377 19144 49393 19178
rect 49561 19144 49577 19178
rect 40775 19094 40809 19110
rect 40775 18902 40809 18918
rect 41033 19094 41067 19110
rect 41033 18902 41067 18918
rect 41147 19094 41181 19110
rect 41147 18902 41181 18918
rect 41405 19094 41439 19110
rect 41405 18902 41439 18918
rect 41519 19094 41553 19110
rect 41519 18902 41553 18918
rect 41777 19094 41811 19110
rect 41777 18902 41811 18918
rect 41891 19094 41925 19110
rect 41891 18902 41925 18918
rect 42149 19094 42183 19110
rect 42149 18902 42183 18918
rect 42263 19094 42297 19110
rect 42263 18902 42297 18918
rect 42521 19094 42555 19110
rect 42521 18902 42555 18918
rect 42635 19094 42669 19110
rect 42635 18902 42669 18918
rect 42893 19094 42927 19110
rect 42893 18902 42927 18918
rect 43007 19094 43041 19110
rect 43007 18902 43041 18918
rect 43265 19094 43299 19110
rect 43265 18902 43299 18918
rect 43379 19094 43413 19110
rect 43379 18902 43413 18918
rect 43637 19094 43671 19110
rect 43637 18902 43671 18918
rect 43751 19094 43785 19110
rect 43751 18902 43785 18918
rect 44009 19094 44043 19110
rect 44009 18902 44043 18918
rect 44123 19094 44157 19110
rect 44123 18902 44157 18918
rect 44381 19094 44415 19110
rect 44381 18902 44415 18918
rect 44495 19094 44529 19110
rect 44495 18902 44529 18918
rect 44753 19094 44787 19110
rect 44753 18902 44787 18918
rect 44867 19094 44901 19110
rect 44867 18902 44901 18918
rect 45125 19094 45159 19110
rect 45125 18902 45159 18918
rect 45239 19094 45273 19110
rect 45239 18902 45273 18918
rect 45497 19094 45531 19110
rect 45497 18902 45531 18918
rect 45611 19094 45645 19110
rect 45611 18902 45645 18918
rect 45869 19094 45903 19110
rect 45869 18902 45903 18918
rect 45983 19094 46017 19110
rect 45983 18902 46017 18918
rect 46241 19094 46275 19110
rect 46241 18902 46275 18918
rect 46355 19094 46389 19110
rect 46355 18902 46389 18918
rect 46613 19094 46647 19110
rect 46613 18902 46647 18918
rect 46727 19094 46761 19110
rect 46727 18902 46761 18918
rect 46985 19094 47019 19110
rect 46985 18902 47019 18918
rect 47099 19094 47133 19110
rect 47099 18902 47133 18918
rect 47357 19094 47391 19110
rect 47357 18902 47391 18918
rect 47471 19094 47505 19110
rect 47471 18902 47505 18918
rect 47729 19094 47763 19110
rect 47729 18902 47763 18918
rect 47843 19094 47877 19110
rect 47843 18902 47877 18918
rect 48101 19094 48135 19110
rect 48101 18902 48135 18918
rect 48215 19094 48249 19110
rect 48215 18902 48249 18918
rect 48473 19094 48507 19110
rect 48473 18902 48507 18918
rect 48587 19094 48621 19110
rect 48587 18902 48621 18918
rect 48845 19094 48879 19110
rect 48845 18902 48879 18918
rect 48959 19094 48993 19110
rect 48959 18902 48993 18918
rect 49217 19094 49251 19110
rect 49217 18902 49251 18918
rect 49331 19094 49365 19110
rect 49331 18902 49365 18918
rect 49589 19094 49623 19110
rect 49589 18902 49623 18918
rect 40821 18834 40837 18868
rect 41005 18834 41021 18868
rect 41193 18834 41209 18868
rect 41377 18834 41393 18868
rect 41565 18834 41581 18868
rect 41749 18834 41765 18868
rect 41937 18834 41953 18868
rect 42121 18834 42137 18868
rect 42309 18834 42325 18868
rect 42493 18834 42509 18868
rect 42681 18834 42697 18868
rect 42865 18834 42881 18868
rect 43053 18834 43069 18868
rect 43237 18834 43253 18868
rect 43425 18834 43441 18868
rect 43609 18834 43625 18868
rect 43797 18834 43813 18868
rect 43981 18834 43997 18868
rect 44169 18834 44185 18868
rect 44353 18834 44369 18868
rect 44541 18834 44557 18868
rect 44725 18834 44741 18868
rect 44913 18834 44929 18868
rect 45097 18834 45113 18868
rect 45285 18834 45301 18868
rect 45469 18834 45485 18868
rect 45657 18834 45673 18868
rect 45841 18834 45857 18868
rect 46029 18834 46045 18868
rect 46213 18834 46229 18868
rect 46401 18834 46417 18868
rect 46585 18834 46601 18868
rect 46773 18834 46789 18868
rect 46957 18834 46973 18868
rect 47145 18834 47161 18868
rect 47329 18834 47345 18868
rect 47517 18834 47533 18868
rect 47701 18834 47717 18868
rect 47889 18834 47905 18868
rect 48073 18834 48089 18868
rect 48261 18834 48277 18868
rect 48445 18834 48461 18868
rect 48633 18834 48649 18868
rect 48817 18834 48833 18868
rect 49005 18834 49021 18868
rect 49189 18834 49205 18868
rect 49377 18834 49393 18868
rect 49561 18834 49577 18868
rect 40821 18726 40837 18760
rect 41005 18726 41021 18760
rect 41193 18726 41209 18760
rect 41377 18726 41393 18760
rect 41565 18726 41581 18760
rect 41749 18726 41765 18760
rect 41937 18726 41953 18760
rect 42121 18726 42137 18760
rect 42309 18726 42325 18760
rect 42493 18726 42509 18760
rect 42681 18726 42697 18760
rect 42865 18726 42881 18760
rect 43053 18726 43069 18760
rect 43237 18726 43253 18760
rect 43425 18726 43441 18760
rect 43609 18726 43625 18760
rect 43797 18726 43813 18760
rect 43981 18726 43997 18760
rect 44169 18726 44185 18760
rect 44353 18726 44369 18760
rect 44541 18726 44557 18760
rect 44725 18726 44741 18760
rect 44913 18726 44929 18760
rect 45097 18726 45113 18760
rect 45285 18726 45301 18760
rect 45469 18726 45485 18760
rect 45657 18726 45673 18760
rect 45841 18726 45857 18760
rect 46029 18726 46045 18760
rect 46213 18726 46229 18760
rect 46401 18726 46417 18760
rect 46585 18726 46601 18760
rect 46773 18726 46789 18760
rect 46957 18726 46973 18760
rect 47145 18726 47161 18760
rect 47329 18726 47345 18760
rect 47517 18726 47533 18760
rect 47701 18726 47717 18760
rect 47889 18726 47905 18760
rect 48073 18726 48089 18760
rect 48261 18726 48277 18760
rect 48445 18726 48461 18760
rect 48633 18726 48649 18760
rect 48817 18726 48833 18760
rect 49005 18726 49021 18760
rect 49189 18726 49205 18760
rect 49377 18726 49393 18760
rect 49561 18726 49577 18760
rect 40775 18676 40809 18692
rect 40775 18484 40809 18500
rect 41033 18676 41067 18692
rect 41033 18484 41067 18500
rect 41147 18676 41181 18692
rect 41147 18484 41181 18500
rect 41405 18676 41439 18692
rect 41405 18484 41439 18500
rect 41519 18676 41553 18692
rect 41519 18484 41553 18500
rect 41777 18676 41811 18692
rect 41777 18484 41811 18500
rect 41891 18676 41925 18692
rect 41891 18484 41925 18500
rect 42149 18676 42183 18692
rect 42149 18484 42183 18500
rect 42263 18676 42297 18692
rect 42263 18484 42297 18500
rect 42521 18676 42555 18692
rect 42521 18484 42555 18500
rect 42635 18676 42669 18692
rect 42635 18484 42669 18500
rect 42893 18676 42927 18692
rect 42893 18484 42927 18500
rect 43007 18676 43041 18692
rect 43007 18484 43041 18500
rect 43265 18676 43299 18692
rect 43265 18484 43299 18500
rect 43379 18676 43413 18692
rect 43379 18484 43413 18500
rect 43637 18676 43671 18692
rect 43637 18484 43671 18500
rect 43751 18676 43785 18692
rect 43751 18484 43785 18500
rect 44009 18676 44043 18692
rect 44009 18484 44043 18500
rect 44123 18676 44157 18692
rect 44123 18484 44157 18500
rect 44381 18676 44415 18692
rect 44381 18484 44415 18500
rect 44495 18676 44529 18692
rect 44495 18484 44529 18500
rect 44753 18676 44787 18692
rect 44753 18484 44787 18500
rect 44867 18676 44901 18692
rect 44867 18484 44901 18500
rect 45125 18676 45159 18692
rect 45125 18484 45159 18500
rect 45239 18676 45273 18692
rect 45239 18484 45273 18500
rect 45497 18676 45531 18692
rect 45497 18484 45531 18500
rect 45611 18676 45645 18692
rect 45611 18484 45645 18500
rect 45869 18676 45903 18692
rect 45869 18484 45903 18500
rect 45983 18676 46017 18692
rect 45983 18484 46017 18500
rect 46241 18676 46275 18692
rect 46241 18484 46275 18500
rect 46355 18676 46389 18692
rect 46355 18484 46389 18500
rect 46613 18676 46647 18692
rect 46613 18484 46647 18500
rect 46727 18676 46761 18692
rect 46727 18484 46761 18500
rect 46985 18676 47019 18692
rect 46985 18484 47019 18500
rect 47099 18676 47133 18692
rect 47099 18484 47133 18500
rect 47357 18676 47391 18692
rect 47357 18484 47391 18500
rect 47471 18676 47505 18692
rect 47471 18484 47505 18500
rect 47729 18676 47763 18692
rect 47729 18484 47763 18500
rect 47843 18676 47877 18692
rect 47843 18484 47877 18500
rect 48101 18676 48135 18692
rect 48101 18484 48135 18500
rect 48215 18676 48249 18692
rect 48215 18484 48249 18500
rect 48473 18676 48507 18692
rect 48473 18484 48507 18500
rect 48587 18676 48621 18692
rect 48587 18484 48621 18500
rect 48845 18676 48879 18692
rect 48845 18484 48879 18500
rect 48959 18676 48993 18692
rect 48959 18484 48993 18500
rect 49217 18676 49251 18692
rect 49217 18484 49251 18500
rect 49331 18676 49365 18692
rect 49331 18484 49365 18500
rect 49589 18676 49623 18692
rect 49589 18484 49623 18500
rect 40821 18416 40837 18450
rect 41005 18416 41021 18450
rect 41193 18416 41209 18450
rect 41377 18416 41393 18450
rect 41565 18416 41581 18450
rect 41749 18416 41765 18450
rect 41937 18416 41953 18450
rect 42121 18416 42137 18450
rect 42309 18416 42325 18450
rect 42493 18416 42509 18450
rect 42681 18416 42697 18450
rect 42865 18416 42881 18450
rect 43053 18416 43069 18450
rect 43237 18416 43253 18450
rect 43425 18416 43441 18450
rect 43609 18416 43625 18450
rect 43797 18416 43813 18450
rect 43981 18416 43997 18450
rect 44169 18416 44185 18450
rect 44353 18416 44369 18450
rect 44541 18416 44557 18450
rect 44725 18416 44741 18450
rect 44913 18416 44929 18450
rect 45097 18416 45113 18450
rect 45285 18416 45301 18450
rect 45469 18416 45485 18450
rect 45657 18416 45673 18450
rect 45841 18416 45857 18450
rect 46029 18416 46045 18450
rect 46213 18416 46229 18450
rect 46401 18416 46417 18450
rect 46585 18416 46601 18450
rect 46773 18416 46789 18450
rect 46957 18416 46973 18450
rect 47145 18416 47161 18450
rect 47329 18416 47345 18450
rect 47517 18416 47533 18450
rect 47701 18416 47717 18450
rect 47889 18416 47905 18450
rect 48073 18416 48089 18450
rect 48261 18416 48277 18450
rect 48445 18416 48461 18450
rect 48633 18416 48649 18450
rect 48817 18416 48833 18450
rect 49005 18416 49021 18450
rect 49189 18416 49205 18450
rect 49377 18416 49393 18450
rect 49561 18416 49577 18450
rect 40821 18308 40837 18342
rect 41005 18308 41021 18342
rect 41193 18308 41209 18342
rect 41377 18308 41393 18342
rect 41565 18308 41581 18342
rect 41749 18308 41765 18342
rect 41937 18308 41953 18342
rect 42121 18308 42137 18342
rect 42309 18308 42325 18342
rect 42493 18308 42509 18342
rect 42681 18308 42697 18342
rect 42865 18308 42881 18342
rect 43053 18308 43069 18342
rect 43237 18308 43253 18342
rect 43425 18308 43441 18342
rect 43609 18308 43625 18342
rect 43797 18308 43813 18342
rect 43981 18308 43997 18342
rect 44169 18308 44185 18342
rect 44353 18308 44369 18342
rect 44541 18308 44557 18342
rect 44725 18308 44741 18342
rect 44913 18308 44929 18342
rect 45097 18308 45113 18342
rect 45285 18308 45301 18342
rect 45469 18308 45485 18342
rect 45657 18308 45673 18342
rect 45841 18308 45857 18342
rect 46029 18308 46045 18342
rect 46213 18308 46229 18342
rect 46401 18308 46417 18342
rect 46585 18308 46601 18342
rect 46773 18308 46789 18342
rect 46957 18308 46973 18342
rect 47145 18308 47161 18342
rect 47329 18308 47345 18342
rect 47517 18308 47533 18342
rect 47701 18308 47717 18342
rect 47889 18308 47905 18342
rect 48073 18308 48089 18342
rect 48261 18308 48277 18342
rect 48445 18308 48461 18342
rect 48633 18308 48649 18342
rect 48817 18308 48833 18342
rect 49005 18308 49021 18342
rect 49189 18308 49205 18342
rect 49377 18308 49393 18342
rect 49561 18308 49577 18342
rect 40775 18258 40809 18274
rect 40775 18066 40809 18082
rect 41033 18258 41067 18274
rect 41033 18066 41067 18082
rect 41147 18258 41181 18274
rect 41147 18066 41181 18082
rect 41405 18258 41439 18274
rect 41405 18066 41439 18082
rect 41519 18258 41553 18274
rect 41519 18066 41553 18082
rect 41777 18258 41811 18274
rect 41777 18066 41811 18082
rect 41891 18258 41925 18274
rect 41891 18066 41925 18082
rect 42149 18258 42183 18274
rect 42149 18066 42183 18082
rect 42263 18258 42297 18274
rect 42263 18066 42297 18082
rect 42521 18258 42555 18274
rect 42521 18066 42555 18082
rect 42635 18258 42669 18274
rect 42635 18066 42669 18082
rect 42893 18258 42927 18274
rect 42893 18066 42927 18082
rect 43007 18258 43041 18274
rect 43007 18066 43041 18082
rect 43265 18258 43299 18274
rect 43265 18066 43299 18082
rect 43379 18258 43413 18274
rect 43379 18066 43413 18082
rect 43637 18258 43671 18274
rect 43637 18066 43671 18082
rect 43751 18258 43785 18274
rect 43751 18066 43785 18082
rect 44009 18258 44043 18274
rect 44009 18066 44043 18082
rect 44123 18258 44157 18274
rect 44123 18066 44157 18082
rect 44381 18258 44415 18274
rect 44381 18066 44415 18082
rect 44495 18258 44529 18274
rect 44495 18066 44529 18082
rect 44753 18258 44787 18274
rect 44753 18066 44787 18082
rect 44867 18258 44901 18274
rect 44867 18066 44901 18082
rect 45125 18258 45159 18274
rect 45125 18066 45159 18082
rect 45239 18258 45273 18274
rect 45239 18066 45273 18082
rect 45497 18258 45531 18274
rect 45497 18066 45531 18082
rect 45611 18258 45645 18274
rect 45611 18066 45645 18082
rect 45869 18258 45903 18274
rect 45869 18066 45903 18082
rect 45983 18258 46017 18274
rect 45983 18066 46017 18082
rect 46241 18258 46275 18274
rect 46241 18066 46275 18082
rect 46355 18258 46389 18274
rect 46355 18066 46389 18082
rect 46613 18258 46647 18274
rect 46613 18066 46647 18082
rect 46727 18258 46761 18274
rect 46727 18066 46761 18082
rect 46985 18258 47019 18274
rect 46985 18066 47019 18082
rect 47099 18258 47133 18274
rect 47099 18066 47133 18082
rect 47357 18258 47391 18274
rect 47357 18066 47391 18082
rect 47471 18258 47505 18274
rect 47471 18066 47505 18082
rect 47729 18258 47763 18274
rect 47729 18066 47763 18082
rect 47843 18258 47877 18274
rect 47843 18066 47877 18082
rect 48101 18258 48135 18274
rect 48101 18066 48135 18082
rect 48215 18258 48249 18274
rect 48215 18066 48249 18082
rect 48473 18258 48507 18274
rect 48473 18066 48507 18082
rect 48587 18258 48621 18274
rect 48587 18066 48621 18082
rect 48845 18258 48879 18274
rect 48845 18066 48879 18082
rect 48959 18258 48993 18274
rect 48959 18066 48993 18082
rect 49217 18258 49251 18274
rect 49217 18066 49251 18082
rect 49331 18258 49365 18274
rect 49331 18066 49365 18082
rect 49589 18258 49623 18274
rect 49589 18066 49623 18082
rect 40821 17998 40837 18032
rect 41005 17998 41021 18032
rect 41193 17998 41209 18032
rect 41377 17998 41393 18032
rect 41565 17998 41581 18032
rect 41749 17998 41765 18032
rect 41937 17998 41953 18032
rect 42121 17998 42137 18032
rect 42309 17998 42325 18032
rect 42493 17998 42509 18032
rect 42681 17998 42697 18032
rect 42865 17998 42881 18032
rect 43053 17998 43069 18032
rect 43237 17998 43253 18032
rect 43425 17998 43441 18032
rect 43609 17998 43625 18032
rect 43797 17998 43813 18032
rect 43981 17998 43997 18032
rect 44169 17998 44185 18032
rect 44353 17998 44369 18032
rect 44541 17998 44557 18032
rect 44725 17998 44741 18032
rect 44913 17998 44929 18032
rect 45097 17998 45113 18032
rect 45285 17998 45301 18032
rect 45469 17998 45485 18032
rect 45657 17998 45673 18032
rect 45841 17998 45857 18032
rect 46029 17998 46045 18032
rect 46213 17998 46229 18032
rect 46401 17998 46417 18032
rect 46585 17998 46601 18032
rect 46773 17998 46789 18032
rect 46957 17998 46973 18032
rect 47145 17998 47161 18032
rect 47329 17998 47345 18032
rect 47517 17998 47533 18032
rect 47701 17998 47717 18032
rect 47889 17998 47905 18032
rect 48073 17998 48089 18032
rect 48261 17998 48277 18032
rect 48445 17998 48461 18032
rect 48633 17998 48649 18032
rect 48817 17998 48833 18032
rect 49005 17998 49021 18032
rect 49189 17998 49205 18032
rect 49377 17998 49393 18032
rect 49561 17998 49577 18032
rect 40661 17930 40695 17992
rect 49703 17930 49737 17992
rect 40661 17896 40757 17930
rect 49641 17896 49737 17930
rect 40661 17442 40757 17476
rect 43689 17442 43785 17476
rect 40661 17380 40695 17442
rect 43751 17380 43785 17442
rect 40821 17340 40837 17374
rect 41005 17340 41021 17374
rect 41193 17340 41209 17374
rect 41377 17340 41393 17374
rect 41565 17340 41581 17374
rect 41749 17340 41765 17374
rect 41937 17340 41953 17374
rect 42121 17340 42137 17374
rect 42309 17340 42325 17374
rect 42493 17340 42509 17374
rect 42681 17340 42697 17374
rect 42865 17340 42881 17374
rect 43053 17340 43069 17374
rect 43237 17340 43253 17374
rect 43425 17340 43441 17374
rect 43609 17340 43625 17374
rect 40775 17281 40809 17297
rect 40775 16489 40809 16505
rect 41033 17281 41067 17297
rect 41033 16489 41067 16505
rect 41147 17281 41181 17297
rect 41147 16489 41181 16505
rect 41405 17281 41439 17297
rect 41405 16489 41439 16505
rect 41519 17281 41553 17297
rect 41519 16489 41553 16505
rect 41777 17281 41811 17297
rect 41777 16489 41811 16505
rect 41891 17281 41925 17297
rect 41891 16489 41925 16505
rect 42149 17281 42183 17297
rect 42149 16489 42183 16505
rect 42263 17281 42297 17297
rect 42263 16489 42297 16505
rect 42521 17281 42555 17297
rect 42521 16489 42555 16505
rect 42635 17281 42669 17297
rect 42635 16489 42669 16505
rect 42893 17281 42927 17297
rect 42893 16489 42927 16505
rect 43007 17281 43041 17297
rect 43007 16489 43041 16505
rect 43265 17281 43299 17297
rect 43265 16489 43299 16505
rect 43379 17281 43413 17297
rect 43379 16489 43413 16505
rect 43637 17281 43671 17297
rect 43637 16489 43671 16505
rect 40821 16412 40837 16446
rect 41005 16412 41021 16446
rect 41193 16412 41209 16446
rect 41377 16412 41393 16446
rect 41565 16412 41581 16446
rect 41749 16412 41765 16446
rect 41937 16412 41953 16446
rect 42121 16412 42137 16446
rect 42309 16412 42325 16446
rect 42493 16412 42509 16446
rect 42681 16412 42697 16446
rect 42865 16412 42881 16446
rect 43053 16412 43069 16446
rect 43237 16412 43253 16446
rect 43425 16412 43441 16446
rect 43609 16412 43625 16446
rect 40821 16304 40837 16338
rect 41005 16304 41021 16338
rect 41193 16304 41209 16338
rect 41377 16304 41393 16338
rect 41565 16304 41581 16338
rect 41749 16304 41765 16338
rect 41937 16304 41953 16338
rect 42121 16304 42137 16338
rect 42309 16304 42325 16338
rect 42493 16304 42509 16338
rect 42681 16304 42697 16338
rect 42865 16304 42881 16338
rect 43053 16304 43069 16338
rect 43237 16304 43253 16338
rect 43425 16304 43441 16338
rect 43609 16304 43625 16338
rect 40775 16245 40809 16261
rect 40775 15453 40809 15469
rect 41033 16245 41067 16261
rect 41033 15453 41067 15469
rect 41147 16245 41181 16261
rect 41147 15453 41181 15469
rect 41405 16245 41439 16261
rect 41405 15453 41439 15469
rect 41519 16245 41553 16261
rect 41519 15453 41553 15469
rect 41777 16245 41811 16261
rect 41777 15453 41811 15469
rect 41891 16245 41925 16261
rect 41891 15453 41925 15469
rect 42149 16245 42183 16261
rect 42149 15453 42183 15469
rect 42263 16245 42297 16261
rect 42263 15453 42297 15469
rect 42521 16245 42555 16261
rect 42521 15453 42555 15469
rect 42635 16245 42669 16261
rect 42635 15453 42669 15469
rect 42893 16245 42927 16261
rect 42893 15453 42927 15469
rect 43007 16245 43041 16261
rect 43007 15453 43041 15469
rect 43265 16245 43299 16261
rect 43265 15453 43299 15469
rect 43379 16245 43413 16261
rect 43379 15453 43413 15469
rect 43637 16245 43671 16261
rect 43637 15453 43671 15469
rect 40821 15376 40837 15410
rect 41005 15376 41021 15410
rect 41193 15376 41209 15410
rect 41377 15376 41393 15410
rect 41565 15376 41581 15410
rect 41749 15376 41765 15410
rect 41937 15376 41953 15410
rect 42121 15376 42137 15410
rect 42309 15376 42325 15410
rect 42493 15376 42509 15410
rect 42681 15376 42697 15410
rect 42865 15376 42881 15410
rect 43053 15376 43069 15410
rect 43237 15376 43253 15410
rect 43425 15376 43441 15410
rect 43609 15376 43625 15410
rect 40821 15268 40837 15302
rect 41005 15268 41021 15302
rect 41193 15268 41209 15302
rect 41377 15268 41393 15302
rect 41565 15268 41581 15302
rect 41749 15268 41765 15302
rect 41937 15268 41953 15302
rect 42121 15268 42137 15302
rect 42309 15268 42325 15302
rect 42493 15268 42509 15302
rect 42681 15268 42697 15302
rect 42865 15268 42881 15302
rect 43053 15268 43069 15302
rect 43237 15268 43253 15302
rect 43425 15268 43441 15302
rect 43609 15268 43625 15302
rect 40775 15209 40809 15225
rect 40775 14417 40809 14433
rect 41033 15209 41067 15225
rect 41033 14417 41067 14433
rect 41147 15209 41181 15225
rect 41147 14417 41181 14433
rect 41405 15209 41439 15225
rect 41405 14417 41439 14433
rect 41519 15209 41553 15225
rect 41519 14417 41553 14433
rect 41777 15209 41811 15225
rect 41777 14417 41811 14433
rect 41891 15209 41925 15225
rect 41891 14417 41925 14433
rect 42149 15209 42183 15225
rect 42149 14417 42183 14433
rect 42263 15209 42297 15225
rect 42263 14417 42297 14433
rect 42521 15209 42555 15225
rect 42521 14417 42555 14433
rect 42635 15209 42669 15225
rect 42635 14417 42669 14433
rect 42893 15209 42927 15225
rect 42893 14417 42927 14433
rect 43007 15209 43041 15225
rect 43007 14417 43041 14433
rect 43265 15209 43299 15225
rect 43265 14417 43299 14433
rect 43379 15209 43413 15225
rect 43379 14417 43413 14433
rect 43637 15209 43671 15225
rect 43637 14417 43671 14433
rect 40821 14340 40837 14374
rect 41005 14340 41021 14374
rect 41193 14340 41209 14374
rect 41377 14340 41393 14374
rect 41565 14340 41581 14374
rect 41749 14340 41765 14374
rect 41937 14340 41953 14374
rect 42121 14340 42137 14374
rect 42309 14340 42325 14374
rect 42493 14340 42509 14374
rect 42681 14340 42697 14374
rect 42865 14340 42881 14374
rect 43053 14340 43069 14374
rect 43237 14340 43253 14374
rect 43425 14340 43441 14374
rect 43609 14340 43625 14374
rect 40821 14232 40837 14266
rect 41005 14232 41021 14266
rect 41193 14232 41209 14266
rect 41377 14232 41393 14266
rect 41565 14232 41581 14266
rect 41749 14232 41765 14266
rect 41937 14232 41953 14266
rect 42121 14232 42137 14266
rect 42309 14232 42325 14266
rect 42493 14232 42509 14266
rect 42681 14232 42697 14266
rect 42865 14232 42881 14266
rect 43053 14232 43069 14266
rect 43237 14232 43253 14266
rect 43425 14232 43441 14266
rect 43609 14232 43625 14266
rect 40775 14173 40809 14189
rect 40775 13381 40809 13397
rect 41033 14173 41067 14189
rect 41033 13381 41067 13397
rect 41147 14173 41181 14189
rect 41147 13381 41181 13397
rect 41405 14173 41439 14189
rect 41405 13381 41439 13397
rect 41519 14173 41553 14189
rect 41519 13381 41553 13397
rect 41777 14173 41811 14189
rect 41777 13381 41811 13397
rect 41891 14173 41925 14189
rect 41891 13381 41925 13397
rect 42149 14173 42183 14189
rect 42149 13381 42183 13397
rect 42263 14173 42297 14189
rect 42263 13381 42297 13397
rect 42521 14173 42555 14189
rect 42521 13381 42555 13397
rect 42635 14173 42669 14189
rect 42635 13381 42669 13397
rect 42893 14173 42927 14189
rect 42893 13381 42927 13397
rect 43007 14173 43041 14189
rect 43007 13381 43041 13397
rect 43265 14173 43299 14189
rect 43265 13381 43299 13397
rect 43379 14173 43413 14189
rect 43379 13381 43413 13397
rect 43637 14173 43671 14189
rect 43637 13381 43671 13397
rect 40821 13304 40837 13338
rect 41005 13304 41021 13338
rect 41193 13304 41209 13338
rect 41377 13304 41393 13338
rect 41565 13304 41581 13338
rect 41749 13304 41765 13338
rect 41937 13304 41953 13338
rect 42121 13304 42137 13338
rect 42309 13304 42325 13338
rect 42493 13304 42509 13338
rect 42681 13304 42697 13338
rect 42865 13304 42881 13338
rect 43053 13304 43069 13338
rect 43237 13304 43253 13338
rect 43425 13304 43441 13338
rect 43609 13304 43625 13338
rect 40661 13236 40695 13298
rect 45825 16548 45921 16582
rect 46059 16548 46155 16582
rect 45825 16486 45859 16548
rect 46121 16486 46155 16548
rect 45825 15392 45859 15454
rect 46121 15392 46155 15454
rect 45825 15358 45921 15392
rect 46059 15358 46155 15392
rect 43751 13236 43785 13298
rect 40661 13202 40746 13236
rect 43689 13202 43785 13236
rect 39173 12818 39269 12852
rect 51129 12818 51225 12852
rect 39173 12756 39207 12818
rect 51191 12756 51225 12818
rect 39333 12716 39349 12750
rect 39517 12716 39533 12750
rect 39705 12716 39721 12750
rect 39889 12716 39905 12750
rect 40077 12716 40093 12750
rect 40261 12716 40277 12750
rect 40449 12716 40465 12750
rect 40633 12716 40649 12750
rect 40821 12716 40837 12750
rect 41005 12716 41021 12750
rect 41193 12716 41209 12750
rect 41377 12716 41393 12750
rect 41565 12716 41581 12750
rect 41749 12716 41765 12750
rect 41937 12716 41953 12750
rect 42121 12716 42137 12750
rect 42309 12716 42325 12750
rect 42493 12716 42509 12750
rect 42681 12716 42697 12750
rect 42865 12716 42881 12750
rect 43053 12716 43069 12750
rect 43237 12716 43253 12750
rect 43425 12716 43441 12750
rect 43609 12716 43625 12750
rect 43797 12716 43813 12750
rect 43981 12716 43997 12750
rect 44169 12716 44185 12750
rect 44353 12716 44369 12750
rect 44541 12716 44557 12750
rect 44725 12716 44741 12750
rect 44913 12716 44929 12750
rect 45097 12716 45113 12750
rect 45285 12716 45301 12750
rect 45469 12716 45485 12750
rect 45657 12716 45673 12750
rect 45841 12716 45857 12750
rect 46029 12716 46045 12750
rect 46213 12716 46229 12750
rect 46401 12716 46417 12750
rect 46585 12716 46601 12750
rect 46773 12716 46789 12750
rect 46957 12716 46973 12750
rect 47145 12716 47161 12750
rect 47329 12716 47345 12750
rect 47517 12716 47533 12750
rect 47701 12716 47717 12750
rect 47889 12716 47905 12750
rect 48073 12716 48089 12750
rect 48261 12716 48277 12750
rect 48445 12716 48461 12750
rect 48633 12716 48649 12750
rect 48817 12716 48833 12750
rect 49005 12716 49021 12750
rect 49189 12716 49205 12750
rect 49377 12716 49393 12750
rect 49561 12716 49577 12750
rect 49749 12716 49765 12750
rect 49933 12716 49949 12750
rect 50121 12716 50137 12750
rect 50305 12716 50321 12750
rect 50493 12716 50509 12750
rect 50677 12716 50693 12750
rect 50865 12716 50881 12750
rect 51049 12716 51065 12750
rect 39287 12657 39321 12673
rect 39287 12265 39321 12281
rect 39545 12657 39579 12673
rect 39545 12265 39579 12281
rect 39659 12657 39693 12673
rect 39659 12265 39693 12281
rect 39917 12657 39951 12673
rect 39917 12265 39951 12281
rect 40031 12657 40065 12673
rect 40031 12265 40065 12281
rect 40289 12657 40323 12673
rect 40289 12265 40323 12281
rect 40403 12657 40437 12673
rect 40403 12265 40437 12281
rect 40661 12657 40695 12673
rect 40661 12265 40695 12281
rect 40775 12657 40809 12673
rect 40775 12265 40809 12281
rect 41033 12657 41067 12673
rect 41033 12265 41067 12281
rect 41147 12657 41181 12673
rect 41147 12265 41181 12281
rect 41405 12657 41439 12673
rect 41405 12265 41439 12281
rect 41519 12657 41553 12673
rect 41519 12265 41553 12281
rect 41777 12657 41811 12673
rect 41777 12265 41811 12281
rect 41891 12657 41925 12673
rect 41891 12265 41925 12281
rect 42149 12657 42183 12673
rect 42149 12265 42183 12281
rect 42263 12657 42297 12673
rect 42263 12265 42297 12281
rect 42521 12657 42555 12673
rect 42521 12265 42555 12281
rect 42635 12657 42669 12673
rect 42635 12265 42669 12281
rect 42893 12657 42927 12673
rect 42893 12265 42927 12281
rect 43007 12657 43041 12673
rect 43007 12265 43041 12281
rect 43265 12657 43299 12673
rect 43265 12265 43299 12281
rect 43379 12657 43413 12673
rect 43379 12265 43413 12281
rect 43637 12657 43671 12673
rect 43637 12265 43671 12281
rect 43751 12657 43785 12673
rect 43751 12265 43785 12281
rect 44009 12657 44043 12673
rect 44009 12265 44043 12281
rect 44123 12657 44157 12673
rect 44123 12265 44157 12281
rect 44381 12657 44415 12673
rect 44381 12265 44415 12281
rect 44495 12657 44529 12673
rect 44495 12265 44529 12281
rect 44753 12657 44787 12673
rect 44753 12265 44787 12281
rect 44867 12657 44901 12673
rect 44867 12265 44901 12281
rect 45125 12657 45159 12673
rect 45125 12265 45159 12281
rect 45239 12657 45273 12673
rect 45239 12265 45273 12281
rect 45497 12657 45531 12673
rect 45497 12265 45531 12281
rect 45611 12657 45645 12673
rect 45611 12265 45645 12281
rect 45869 12657 45903 12673
rect 45869 12265 45903 12281
rect 45983 12657 46017 12673
rect 45983 12265 46017 12281
rect 46241 12657 46275 12673
rect 46241 12265 46275 12281
rect 46355 12657 46389 12673
rect 46355 12265 46389 12281
rect 46613 12657 46647 12673
rect 46613 12265 46647 12281
rect 46727 12657 46761 12673
rect 46727 12265 46761 12281
rect 46985 12657 47019 12673
rect 46985 12265 47019 12281
rect 47099 12657 47133 12673
rect 47099 12265 47133 12281
rect 47357 12657 47391 12673
rect 47357 12265 47391 12281
rect 47471 12657 47505 12673
rect 47471 12265 47505 12281
rect 47729 12657 47763 12673
rect 47729 12265 47763 12281
rect 47843 12657 47877 12673
rect 47843 12265 47877 12281
rect 48101 12657 48135 12673
rect 48101 12265 48135 12281
rect 48215 12657 48249 12673
rect 48215 12265 48249 12281
rect 48473 12657 48507 12673
rect 48473 12265 48507 12281
rect 48587 12657 48621 12673
rect 48587 12265 48621 12281
rect 48845 12657 48879 12673
rect 48845 12265 48879 12281
rect 48959 12657 48993 12673
rect 48959 12265 48993 12281
rect 49217 12657 49251 12673
rect 49217 12265 49251 12281
rect 49331 12657 49365 12673
rect 49331 12265 49365 12281
rect 49589 12657 49623 12673
rect 49589 12265 49623 12281
rect 49703 12657 49737 12673
rect 49703 12265 49737 12281
rect 49961 12657 49995 12673
rect 49961 12265 49995 12281
rect 50075 12657 50109 12673
rect 50075 12265 50109 12281
rect 50333 12657 50367 12673
rect 50333 12265 50367 12281
rect 50447 12657 50481 12673
rect 50447 12265 50481 12281
rect 50705 12657 50739 12673
rect 50705 12265 50739 12281
rect 50819 12657 50853 12673
rect 50819 12265 50853 12281
rect 51077 12657 51111 12673
rect 51077 12265 51111 12281
rect 39333 12188 39349 12222
rect 39517 12188 39533 12222
rect 39705 12188 39721 12222
rect 39889 12188 39905 12222
rect 40077 12188 40093 12222
rect 40261 12188 40277 12222
rect 40449 12188 40465 12222
rect 40633 12188 40649 12222
rect 40821 12188 40837 12222
rect 41005 12188 41021 12222
rect 41193 12188 41209 12222
rect 41377 12188 41393 12222
rect 41565 12188 41581 12222
rect 41749 12188 41765 12222
rect 41937 12188 41953 12222
rect 42121 12188 42137 12222
rect 42309 12188 42325 12222
rect 42493 12188 42509 12222
rect 42681 12188 42697 12222
rect 42865 12188 42881 12222
rect 43053 12188 43069 12222
rect 43237 12188 43253 12222
rect 43425 12188 43441 12222
rect 43609 12188 43625 12222
rect 43797 12188 43813 12222
rect 43981 12188 43997 12222
rect 44169 12188 44185 12222
rect 44353 12188 44369 12222
rect 44541 12188 44557 12222
rect 44725 12188 44741 12222
rect 44913 12188 44929 12222
rect 45097 12188 45113 12222
rect 45285 12188 45301 12222
rect 45469 12188 45485 12222
rect 45657 12188 45673 12222
rect 45841 12188 45857 12222
rect 46029 12188 46045 12222
rect 46213 12188 46229 12222
rect 46401 12188 46417 12222
rect 46585 12188 46601 12222
rect 46773 12188 46789 12222
rect 46957 12188 46973 12222
rect 47145 12188 47161 12222
rect 47329 12188 47345 12222
rect 47517 12188 47533 12222
rect 47701 12188 47717 12222
rect 47889 12188 47905 12222
rect 48073 12188 48089 12222
rect 48261 12188 48277 12222
rect 48445 12188 48461 12222
rect 48633 12188 48649 12222
rect 48817 12188 48833 12222
rect 49005 12188 49021 12222
rect 49189 12188 49205 12222
rect 49377 12188 49393 12222
rect 49561 12188 49577 12222
rect 49749 12188 49765 12222
rect 49933 12188 49949 12222
rect 50121 12188 50137 12222
rect 50305 12188 50321 12222
rect 50493 12188 50509 12222
rect 50677 12188 50693 12222
rect 50865 12188 50881 12222
rect 51049 12188 51065 12222
rect 39333 12080 39349 12114
rect 39517 12080 39533 12114
rect 39705 12080 39721 12114
rect 39889 12080 39905 12114
rect 40077 12080 40093 12114
rect 40261 12080 40277 12114
rect 40449 12080 40465 12114
rect 40633 12080 40649 12114
rect 40821 12080 40837 12114
rect 41005 12080 41021 12114
rect 41193 12080 41209 12114
rect 41377 12080 41393 12114
rect 41565 12080 41581 12114
rect 41749 12080 41765 12114
rect 41937 12080 41953 12114
rect 42121 12080 42137 12114
rect 42309 12080 42325 12114
rect 42493 12080 42509 12114
rect 42681 12080 42697 12114
rect 42865 12080 42881 12114
rect 43053 12080 43069 12114
rect 43237 12080 43253 12114
rect 43425 12080 43441 12114
rect 43609 12080 43625 12114
rect 43797 12080 43813 12114
rect 43981 12080 43997 12114
rect 44169 12080 44185 12114
rect 44353 12080 44369 12114
rect 44541 12080 44557 12114
rect 44725 12080 44741 12114
rect 44913 12080 44929 12114
rect 45097 12080 45113 12114
rect 45285 12080 45301 12114
rect 45469 12080 45485 12114
rect 45657 12080 45673 12114
rect 45841 12080 45857 12114
rect 46029 12080 46045 12114
rect 46213 12080 46229 12114
rect 46401 12080 46417 12114
rect 46585 12080 46601 12114
rect 46773 12080 46789 12114
rect 46957 12080 46973 12114
rect 47145 12080 47161 12114
rect 47329 12080 47345 12114
rect 47517 12080 47533 12114
rect 47701 12080 47717 12114
rect 47889 12080 47905 12114
rect 48073 12080 48089 12114
rect 48261 12080 48277 12114
rect 48445 12080 48461 12114
rect 48633 12080 48649 12114
rect 48817 12080 48833 12114
rect 49005 12080 49021 12114
rect 49189 12080 49205 12114
rect 49377 12080 49393 12114
rect 49561 12080 49577 12114
rect 49749 12080 49765 12114
rect 49933 12080 49949 12114
rect 50121 12080 50137 12114
rect 50305 12080 50321 12114
rect 50493 12080 50509 12114
rect 50677 12080 50693 12114
rect 50865 12080 50881 12114
rect 51049 12080 51065 12114
rect 39287 12021 39321 12037
rect 39287 11629 39321 11645
rect 39545 12021 39579 12037
rect 39545 11629 39579 11645
rect 39659 12021 39693 12037
rect 39659 11629 39693 11645
rect 39917 12021 39951 12037
rect 39917 11629 39951 11645
rect 40031 12021 40065 12037
rect 40031 11629 40065 11645
rect 40289 12021 40323 12037
rect 40289 11629 40323 11645
rect 40403 12021 40437 12037
rect 40403 11629 40437 11645
rect 40661 12021 40695 12037
rect 40661 11629 40695 11645
rect 40775 12021 40809 12037
rect 40775 11629 40809 11645
rect 41033 12021 41067 12037
rect 41033 11629 41067 11645
rect 41147 12021 41181 12037
rect 41147 11629 41181 11645
rect 41405 12021 41439 12037
rect 41405 11629 41439 11645
rect 41519 12021 41553 12037
rect 41519 11629 41553 11645
rect 41777 12021 41811 12037
rect 41777 11629 41811 11645
rect 41891 12021 41925 12037
rect 41891 11629 41925 11645
rect 42149 12021 42183 12037
rect 42149 11629 42183 11645
rect 42263 12021 42297 12037
rect 42263 11629 42297 11645
rect 42521 12021 42555 12037
rect 42521 11629 42555 11645
rect 42635 12021 42669 12037
rect 42635 11629 42669 11645
rect 42893 12021 42927 12037
rect 42893 11629 42927 11645
rect 43007 12021 43041 12037
rect 43007 11629 43041 11645
rect 43265 12021 43299 12037
rect 43265 11629 43299 11645
rect 43379 12021 43413 12037
rect 43379 11629 43413 11645
rect 43637 12021 43671 12037
rect 43637 11629 43671 11645
rect 43751 12021 43785 12037
rect 43751 11629 43785 11645
rect 44009 12021 44043 12037
rect 44009 11629 44043 11645
rect 44123 12021 44157 12037
rect 44123 11629 44157 11645
rect 44381 12021 44415 12037
rect 44381 11629 44415 11645
rect 44495 12021 44529 12037
rect 44495 11629 44529 11645
rect 44753 12021 44787 12037
rect 44753 11629 44787 11645
rect 44867 12021 44901 12037
rect 44867 11629 44901 11645
rect 45125 12021 45159 12037
rect 45125 11629 45159 11645
rect 45239 12021 45273 12037
rect 45239 11629 45273 11645
rect 45497 12021 45531 12037
rect 45497 11629 45531 11645
rect 45611 12021 45645 12037
rect 45611 11629 45645 11645
rect 45869 12021 45903 12037
rect 45869 11629 45903 11645
rect 45983 12021 46017 12037
rect 45983 11629 46017 11645
rect 46241 12021 46275 12037
rect 46241 11629 46275 11645
rect 46355 12021 46389 12037
rect 46355 11629 46389 11645
rect 46613 12021 46647 12037
rect 46613 11629 46647 11645
rect 46727 12021 46761 12037
rect 46727 11629 46761 11645
rect 46985 12021 47019 12037
rect 46985 11629 47019 11645
rect 47099 12021 47133 12037
rect 47099 11629 47133 11645
rect 47357 12021 47391 12037
rect 47357 11629 47391 11645
rect 47471 12021 47505 12037
rect 47471 11629 47505 11645
rect 47729 12021 47763 12037
rect 47729 11629 47763 11645
rect 47843 12021 47877 12037
rect 47843 11629 47877 11645
rect 48101 12021 48135 12037
rect 48101 11629 48135 11645
rect 48215 12021 48249 12037
rect 48215 11629 48249 11645
rect 48473 12021 48507 12037
rect 48473 11629 48507 11645
rect 48587 12021 48621 12037
rect 48587 11629 48621 11645
rect 48845 12021 48879 12037
rect 48845 11629 48879 11645
rect 48959 12021 48993 12037
rect 48959 11629 48993 11645
rect 49217 12021 49251 12037
rect 49217 11629 49251 11645
rect 49331 12021 49365 12037
rect 49331 11629 49365 11645
rect 49589 12021 49623 12037
rect 49589 11629 49623 11645
rect 49703 12021 49737 12037
rect 49703 11629 49737 11645
rect 49961 12021 49995 12037
rect 49961 11629 49995 11645
rect 50075 12021 50109 12037
rect 50075 11629 50109 11645
rect 50333 12021 50367 12037
rect 50333 11629 50367 11645
rect 50447 12021 50481 12037
rect 50447 11629 50481 11645
rect 50705 12021 50739 12037
rect 50705 11629 50739 11645
rect 50819 12021 50853 12037
rect 50819 11629 50853 11645
rect 51077 12021 51111 12037
rect 51077 11629 51111 11645
rect 39333 11552 39349 11586
rect 39517 11552 39533 11586
rect 39705 11552 39721 11586
rect 39889 11552 39905 11586
rect 40077 11552 40093 11586
rect 40261 11552 40277 11586
rect 40449 11552 40465 11586
rect 40633 11552 40649 11586
rect 40821 11552 40837 11586
rect 41005 11552 41021 11586
rect 41193 11552 41209 11586
rect 41377 11552 41393 11586
rect 41565 11552 41581 11586
rect 41749 11552 41765 11586
rect 41937 11552 41953 11586
rect 42121 11552 42137 11586
rect 42309 11552 42325 11586
rect 42493 11552 42509 11586
rect 42681 11552 42697 11586
rect 42865 11552 42881 11586
rect 43053 11552 43069 11586
rect 43237 11552 43253 11586
rect 43425 11552 43441 11586
rect 43609 11552 43625 11586
rect 43797 11552 43813 11586
rect 43981 11552 43997 11586
rect 44169 11552 44185 11586
rect 44353 11552 44369 11586
rect 44541 11552 44557 11586
rect 44725 11552 44741 11586
rect 44913 11552 44929 11586
rect 45097 11552 45113 11586
rect 45285 11552 45301 11586
rect 45469 11552 45485 11586
rect 45657 11552 45673 11586
rect 45841 11552 45857 11586
rect 46029 11552 46045 11586
rect 46213 11552 46229 11586
rect 46401 11552 46417 11586
rect 46585 11552 46601 11586
rect 46773 11552 46789 11586
rect 46957 11552 46973 11586
rect 47145 11552 47161 11586
rect 47329 11552 47345 11586
rect 47517 11552 47533 11586
rect 47701 11552 47717 11586
rect 47889 11552 47905 11586
rect 48073 11552 48089 11586
rect 48261 11552 48277 11586
rect 48445 11552 48461 11586
rect 48633 11552 48649 11586
rect 48817 11552 48833 11586
rect 49005 11552 49021 11586
rect 49189 11552 49205 11586
rect 49377 11552 49393 11586
rect 49561 11552 49577 11586
rect 49749 11552 49765 11586
rect 49933 11552 49949 11586
rect 50121 11552 50137 11586
rect 50305 11552 50321 11586
rect 50493 11552 50509 11586
rect 50677 11552 50693 11586
rect 50865 11552 50881 11586
rect 51049 11552 51065 11586
rect 39333 11444 39349 11478
rect 39517 11444 39533 11478
rect 39705 11444 39721 11478
rect 39889 11444 39905 11478
rect 40077 11444 40093 11478
rect 40261 11444 40277 11478
rect 40449 11444 40465 11478
rect 40633 11444 40649 11478
rect 40821 11444 40837 11478
rect 41005 11444 41021 11478
rect 41193 11444 41209 11478
rect 41377 11444 41393 11478
rect 41565 11444 41581 11478
rect 41749 11444 41765 11478
rect 41937 11444 41953 11478
rect 42121 11444 42137 11478
rect 42309 11444 42325 11478
rect 42493 11444 42509 11478
rect 42681 11444 42697 11478
rect 42865 11444 42881 11478
rect 43053 11444 43069 11478
rect 43237 11444 43253 11478
rect 43425 11444 43441 11478
rect 43609 11444 43625 11478
rect 43797 11444 43813 11478
rect 43981 11444 43997 11478
rect 44169 11444 44185 11478
rect 44353 11444 44369 11478
rect 44541 11444 44557 11478
rect 44725 11444 44741 11478
rect 44913 11444 44929 11478
rect 45097 11444 45113 11478
rect 45285 11444 45301 11478
rect 45469 11444 45485 11478
rect 45657 11444 45673 11478
rect 45841 11444 45857 11478
rect 46029 11444 46045 11478
rect 46213 11444 46229 11478
rect 46401 11444 46417 11478
rect 46585 11444 46601 11478
rect 46773 11444 46789 11478
rect 46957 11444 46973 11478
rect 47145 11444 47161 11478
rect 47329 11444 47345 11478
rect 47517 11444 47533 11478
rect 47701 11444 47717 11478
rect 47889 11444 47905 11478
rect 48073 11444 48089 11478
rect 48261 11444 48277 11478
rect 48445 11444 48461 11478
rect 48633 11444 48649 11478
rect 48817 11444 48833 11478
rect 49005 11444 49021 11478
rect 49189 11444 49205 11478
rect 49377 11444 49393 11478
rect 49561 11444 49577 11478
rect 49749 11444 49765 11478
rect 49933 11444 49949 11478
rect 50121 11444 50137 11478
rect 50305 11444 50321 11478
rect 50493 11444 50509 11478
rect 50677 11444 50693 11478
rect 50865 11444 50881 11478
rect 51049 11444 51065 11478
rect 39287 11385 39321 11401
rect 39287 10993 39321 11009
rect 39545 11385 39579 11401
rect 39545 10993 39579 11009
rect 39659 11385 39693 11401
rect 39659 10993 39693 11009
rect 39917 11385 39951 11401
rect 39917 10993 39951 11009
rect 40031 11385 40065 11401
rect 40031 10993 40065 11009
rect 40289 11385 40323 11401
rect 40289 10993 40323 11009
rect 40403 11385 40437 11401
rect 40403 10993 40437 11009
rect 40661 11385 40695 11401
rect 40661 10993 40695 11009
rect 40775 11385 40809 11401
rect 40775 10993 40809 11009
rect 41033 11385 41067 11401
rect 41033 10993 41067 11009
rect 41147 11385 41181 11401
rect 41147 10993 41181 11009
rect 41405 11385 41439 11401
rect 41405 10993 41439 11009
rect 41519 11385 41553 11401
rect 41519 10993 41553 11009
rect 41777 11385 41811 11401
rect 41777 10993 41811 11009
rect 41891 11385 41925 11401
rect 41891 10993 41925 11009
rect 42149 11385 42183 11401
rect 42149 10993 42183 11009
rect 42263 11385 42297 11401
rect 42263 10993 42297 11009
rect 42521 11385 42555 11401
rect 42521 10993 42555 11009
rect 42635 11385 42669 11401
rect 42635 10993 42669 11009
rect 42893 11385 42927 11401
rect 42893 10993 42927 11009
rect 43007 11385 43041 11401
rect 43007 10993 43041 11009
rect 43265 11385 43299 11401
rect 43265 10993 43299 11009
rect 43379 11385 43413 11401
rect 43379 10993 43413 11009
rect 43637 11385 43671 11401
rect 43637 10993 43671 11009
rect 43751 11385 43785 11401
rect 43751 10993 43785 11009
rect 44009 11385 44043 11401
rect 44009 10993 44043 11009
rect 44123 11385 44157 11401
rect 44123 10993 44157 11009
rect 44381 11385 44415 11401
rect 44381 10993 44415 11009
rect 44495 11385 44529 11401
rect 44495 10993 44529 11009
rect 44753 11385 44787 11401
rect 44753 10993 44787 11009
rect 44867 11385 44901 11401
rect 44867 10993 44901 11009
rect 45125 11385 45159 11401
rect 45125 10993 45159 11009
rect 45239 11385 45273 11401
rect 45239 10993 45273 11009
rect 45497 11385 45531 11401
rect 45497 10993 45531 11009
rect 45611 11385 45645 11401
rect 45611 10993 45645 11009
rect 45869 11385 45903 11401
rect 45869 10993 45903 11009
rect 45983 11385 46017 11401
rect 45983 10993 46017 11009
rect 46241 11385 46275 11401
rect 46241 10993 46275 11009
rect 46355 11385 46389 11401
rect 46355 10993 46389 11009
rect 46613 11385 46647 11401
rect 46613 10993 46647 11009
rect 46727 11385 46761 11401
rect 46727 10993 46761 11009
rect 46985 11385 47019 11401
rect 46985 10993 47019 11009
rect 47099 11385 47133 11401
rect 47099 10993 47133 11009
rect 47357 11385 47391 11401
rect 47357 10993 47391 11009
rect 47471 11385 47505 11401
rect 47471 10993 47505 11009
rect 47729 11385 47763 11401
rect 47729 10993 47763 11009
rect 47843 11385 47877 11401
rect 47843 10993 47877 11009
rect 48101 11385 48135 11401
rect 48101 10993 48135 11009
rect 48215 11385 48249 11401
rect 48215 10993 48249 11009
rect 48473 11385 48507 11401
rect 48473 10993 48507 11009
rect 48587 11385 48621 11401
rect 48587 10993 48621 11009
rect 48845 11385 48879 11401
rect 48845 10993 48879 11009
rect 48959 11385 48993 11401
rect 48959 10993 48993 11009
rect 49217 11385 49251 11401
rect 49217 10993 49251 11009
rect 49331 11385 49365 11401
rect 49331 10993 49365 11009
rect 49589 11385 49623 11401
rect 49589 10993 49623 11009
rect 49703 11385 49737 11401
rect 49703 10993 49737 11009
rect 49961 11385 49995 11401
rect 49961 10993 49995 11009
rect 50075 11385 50109 11401
rect 50075 10993 50109 11009
rect 50333 11385 50367 11401
rect 50333 10993 50367 11009
rect 50447 11385 50481 11401
rect 50447 10993 50481 11009
rect 50705 11385 50739 11401
rect 50705 10993 50739 11009
rect 50819 11385 50853 11401
rect 50819 10993 50853 11009
rect 51077 11385 51111 11401
rect 51077 10993 51111 11009
rect 39333 10916 39349 10950
rect 39517 10916 39533 10950
rect 39705 10916 39721 10950
rect 39889 10916 39905 10950
rect 40077 10916 40093 10950
rect 40261 10916 40277 10950
rect 40449 10916 40465 10950
rect 40633 10916 40649 10950
rect 40821 10916 40837 10950
rect 41005 10916 41021 10950
rect 41193 10916 41209 10950
rect 41377 10916 41393 10950
rect 41565 10916 41581 10950
rect 41749 10916 41765 10950
rect 41937 10916 41953 10950
rect 42121 10916 42137 10950
rect 42309 10916 42325 10950
rect 42493 10916 42509 10950
rect 42681 10916 42697 10950
rect 42865 10916 42881 10950
rect 43053 10916 43069 10950
rect 43237 10916 43253 10950
rect 43425 10916 43441 10950
rect 43609 10916 43625 10950
rect 43797 10916 43813 10950
rect 43981 10916 43997 10950
rect 44169 10916 44185 10950
rect 44353 10916 44369 10950
rect 44541 10916 44557 10950
rect 44725 10916 44741 10950
rect 44913 10916 44929 10950
rect 45097 10916 45113 10950
rect 45285 10916 45301 10950
rect 45469 10916 45485 10950
rect 45657 10916 45673 10950
rect 45841 10916 45857 10950
rect 46029 10916 46045 10950
rect 46213 10916 46229 10950
rect 46401 10916 46417 10950
rect 46585 10916 46601 10950
rect 46773 10916 46789 10950
rect 46957 10916 46973 10950
rect 47145 10916 47161 10950
rect 47329 10916 47345 10950
rect 47517 10916 47533 10950
rect 47701 10916 47717 10950
rect 47889 10916 47905 10950
rect 48073 10916 48089 10950
rect 48261 10916 48277 10950
rect 48445 10916 48461 10950
rect 48633 10916 48649 10950
rect 48817 10916 48833 10950
rect 49005 10916 49021 10950
rect 49189 10916 49205 10950
rect 49377 10916 49393 10950
rect 49561 10916 49577 10950
rect 49749 10916 49765 10950
rect 49933 10916 49949 10950
rect 50121 10916 50137 10950
rect 50305 10916 50321 10950
rect 50493 10916 50509 10950
rect 50677 10916 50693 10950
rect 50865 10916 50881 10950
rect 51049 10916 51065 10950
rect 39173 10848 39207 10910
rect 51191 10848 51225 10910
rect 39173 10814 39269 10848
rect 51132 10814 51225 10848
rect 39173 9017 39269 9051
rect 51132 9017 51225 9051
rect 39173 8955 39207 9017
rect 51191 8955 51225 9017
rect 39333 8915 39349 8949
rect 39517 8915 39533 8949
rect 39705 8915 39721 8949
rect 39889 8915 39905 8949
rect 40077 8915 40093 8949
rect 40261 8915 40277 8949
rect 40449 8915 40465 8949
rect 40633 8915 40649 8949
rect 40821 8915 40837 8949
rect 41005 8915 41021 8949
rect 41193 8915 41209 8949
rect 41377 8915 41393 8949
rect 41565 8915 41581 8949
rect 41749 8915 41765 8949
rect 41937 8915 41953 8949
rect 42121 8915 42137 8949
rect 42309 8915 42325 8949
rect 42493 8915 42509 8949
rect 42681 8915 42697 8949
rect 42865 8915 42881 8949
rect 43053 8915 43069 8949
rect 43237 8915 43253 8949
rect 43425 8915 43441 8949
rect 43609 8915 43625 8949
rect 43797 8915 43813 8949
rect 43981 8915 43997 8949
rect 44169 8915 44185 8949
rect 44353 8915 44369 8949
rect 44541 8915 44557 8949
rect 44725 8915 44741 8949
rect 44913 8915 44929 8949
rect 45097 8915 45113 8949
rect 45285 8915 45301 8949
rect 45469 8915 45485 8949
rect 45657 8915 45673 8949
rect 45841 8915 45857 8949
rect 46029 8915 46045 8949
rect 46213 8915 46229 8949
rect 46401 8915 46417 8949
rect 46585 8915 46601 8949
rect 46773 8915 46789 8949
rect 46957 8915 46973 8949
rect 47145 8915 47161 8949
rect 47329 8915 47345 8949
rect 47517 8915 47533 8949
rect 47701 8915 47717 8949
rect 47889 8915 47905 8949
rect 48073 8915 48089 8949
rect 48261 8915 48277 8949
rect 48445 8915 48461 8949
rect 48633 8915 48649 8949
rect 48817 8915 48833 8949
rect 49005 8915 49021 8949
rect 49189 8915 49205 8949
rect 49377 8915 49393 8949
rect 49561 8915 49577 8949
rect 49749 8915 49765 8949
rect 49933 8915 49949 8949
rect 50121 8915 50137 8949
rect 50305 8915 50321 8949
rect 50493 8915 50509 8949
rect 50677 8915 50693 8949
rect 50865 8915 50881 8949
rect 51049 8915 51065 8949
rect 39287 8856 39321 8872
rect 39287 8464 39321 8480
rect 39545 8856 39579 8872
rect 39545 8464 39579 8480
rect 39659 8856 39693 8872
rect 39659 8464 39693 8480
rect 39917 8856 39951 8872
rect 39917 8464 39951 8480
rect 40031 8856 40065 8872
rect 40031 8464 40065 8480
rect 40289 8856 40323 8872
rect 40289 8464 40323 8480
rect 40403 8856 40437 8872
rect 40403 8464 40437 8480
rect 40661 8856 40695 8872
rect 40661 8464 40695 8480
rect 40775 8856 40809 8872
rect 40775 8464 40809 8480
rect 41033 8856 41067 8872
rect 41033 8464 41067 8480
rect 41147 8856 41181 8872
rect 41147 8464 41181 8480
rect 41405 8856 41439 8872
rect 41405 8464 41439 8480
rect 41519 8856 41553 8872
rect 41519 8464 41553 8480
rect 41777 8856 41811 8872
rect 41777 8464 41811 8480
rect 41891 8856 41925 8872
rect 41891 8464 41925 8480
rect 42149 8856 42183 8872
rect 42149 8464 42183 8480
rect 42263 8856 42297 8872
rect 42263 8464 42297 8480
rect 42521 8856 42555 8872
rect 42521 8464 42555 8480
rect 42635 8856 42669 8872
rect 42635 8464 42669 8480
rect 42893 8856 42927 8872
rect 42893 8464 42927 8480
rect 43007 8856 43041 8872
rect 43007 8464 43041 8480
rect 43265 8856 43299 8872
rect 43265 8464 43299 8480
rect 43379 8856 43413 8872
rect 43379 8464 43413 8480
rect 43637 8856 43671 8872
rect 43637 8464 43671 8480
rect 43751 8856 43785 8872
rect 43751 8464 43785 8480
rect 44009 8856 44043 8872
rect 44009 8464 44043 8480
rect 44123 8856 44157 8872
rect 44123 8464 44157 8480
rect 44381 8856 44415 8872
rect 44381 8464 44415 8480
rect 44495 8856 44529 8872
rect 44495 8464 44529 8480
rect 44753 8856 44787 8872
rect 44753 8464 44787 8480
rect 44867 8856 44901 8872
rect 44867 8464 44901 8480
rect 45125 8856 45159 8872
rect 45125 8464 45159 8480
rect 45239 8856 45273 8872
rect 45239 8464 45273 8480
rect 45497 8856 45531 8872
rect 45497 8464 45531 8480
rect 45611 8856 45645 8872
rect 45611 8464 45645 8480
rect 45869 8856 45903 8872
rect 45869 8464 45903 8480
rect 45983 8856 46017 8872
rect 45983 8464 46017 8480
rect 46241 8856 46275 8872
rect 46241 8464 46275 8480
rect 46355 8856 46389 8872
rect 46355 8464 46389 8480
rect 46613 8856 46647 8872
rect 46613 8464 46647 8480
rect 46727 8856 46761 8872
rect 46727 8464 46761 8480
rect 46985 8856 47019 8872
rect 46985 8464 47019 8480
rect 47099 8856 47133 8872
rect 47099 8464 47133 8480
rect 47357 8856 47391 8872
rect 47357 8464 47391 8480
rect 47471 8856 47505 8872
rect 47471 8464 47505 8480
rect 47729 8856 47763 8872
rect 47729 8464 47763 8480
rect 47843 8856 47877 8872
rect 47843 8464 47877 8480
rect 48101 8856 48135 8872
rect 48101 8464 48135 8480
rect 48215 8856 48249 8872
rect 48215 8464 48249 8480
rect 48473 8856 48507 8872
rect 48473 8464 48507 8480
rect 48587 8856 48621 8872
rect 48587 8464 48621 8480
rect 48845 8856 48879 8872
rect 48845 8464 48879 8480
rect 48959 8856 48993 8872
rect 48959 8464 48993 8480
rect 49217 8856 49251 8872
rect 49217 8464 49251 8480
rect 49331 8856 49365 8872
rect 49331 8464 49365 8480
rect 49589 8856 49623 8872
rect 49589 8464 49623 8480
rect 49703 8856 49737 8872
rect 49703 8464 49737 8480
rect 49961 8856 49995 8872
rect 49961 8464 49995 8480
rect 50075 8856 50109 8872
rect 50075 8464 50109 8480
rect 50333 8856 50367 8872
rect 50333 8464 50367 8480
rect 50447 8856 50481 8872
rect 50447 8464 50481 8480
rect 50705 8856 50739 8872
rect 50705 8464 50739 8480
rect 50819 8856 50853 8872
rect 50819 8464 50853 8480
rect 51077 8856 51111 8872
rect 51077 8464 51111 8480
rect 39333 8387 39349 8421
rect 39517 8387 39533 8421
rect 39705 8387 39721 8421
rect 39889 8387 39905 8421
rect 40077 8387 40093 8421
rect 40261 8387 40277 8421
rect 40449 8387 40465 8421
rect 40633 8387 40649 8421
rect 40821 8387 40837 8421
rect 41005 8387 41021 8421
rect 41193 8387 41209 8421
rect 41377 8387 41393 8421
rect 41565 8387 41581 8421
rect 41749 8387 41765 8421
rect 41937 8387 41953 8421
rect 42121 8387 42137 8421
rect 42309 8387 42325 8421
rect 42493 8387 42509 8421
rect 42681 8387 42697 8421
rect 42865 8387 42881 8421
rect 43053 8387 43069 8421
rect 43237 8387 43253 8421
rect 43425 8387 43441 8421
rect 43609 8387 43625 8421
rect 43797 8387 43813 8421
rect 43981 8387 43997 8421
rect 44169 8387 44185 8421
rect 44353 8387 44369 8421
rect 44541 8387 44557 8421
rect 44725 8387 44741 8421
rect 44913 8387 44929 8421
rect 45097 8387 45113 8421
rect 45285 8387 45301 8421
rect 45469 8387 45485 8421
rect 45657 8387 45673 8421
rect 45841 8387 45857 8421
rect 46029 8387 46045 8421
rect 46213 8387 46229 8421
rect 46401 8387 46417 8421
rect 46585 8387 46601 8421
rect 46773 8387 46789 8421
rect 46957 8387 46973 8421
rect 47145 8387 47161 8421
rect 47329 8387 47345 8421
rect 47517 8387 47533 8421
rect 47701 8387 47717 8421
rect 47889 8387 47905 8421
rect 48073 8387 48089 8421
rect 48261 8387 48277 8421
rect 48445 8387 48461 8421
rect 48633 8387 48649 8421
rect 48817 8387 48833 8421
rect 49005 8387 49021 8421
rect 49189 8387 49205 8421
rect 49377 8387 49393 8421
rect 49561 8387 49577 8421
rect 49749 8387 49765 8421
rect 49933 8387 49949 8421
rect 50121 8387 50137 8421
rect 50305 8387 50321 8421
rect 50493 8387 50509 8421
rect 50677 8387 50693 8421
rect 50865 8387 50881 8421
rect 51049 8387 51065 8421
rect 39333 8279 39349 8313
rect 39517 8279 39533 8313
rect 39705 8279 39721 8313
rect 39889 8279 39905 8313
rect 40077 8279 40093 8313
rect 40261 8279 40277 8313
rect 40449 8279 40465 8313
rect 40633 8279 40649 8313
rect 40821 8279 40837 8313
rect 41005 8279 41021 8313
rect 41193 8279 41209 8313
rect 41377 8279 41393 8313
rect 41565 8279 41581 8313
rect 41749 8279 41765 8313
rect 41937 8279 41953 8313
rect 42121 8279 42137 8313
rect 42309 8279 42325 8313
rect 42493 8279 42509 8313
rect 42681 8279 42697 8313
rect 42865 8279 42881 8313
rect 43053 8279 43069 8313
rect 43237 8279 43253 8313
rect 43425 8279 43441 8313
rect 43609 8279 43625 8313
rect 43797 8279 43813 8313
rect 43981 8279 43997 8313
rect 44169 8279 44185 8313
rect 44353 8279 44369 8313
rect 44541 8279 44557 8313
rect 44725 8279 44741 8313
rect 44913 8279 44929 8313
rect 45097 8279 45113 8313
rect 45285 8279 45301 8313
rect 45469 8279 45485 8313
rect 45657 8279 45673 8313
rect 45841 8279 45857 8313
rect 46029 8279 46045 8313
rect 46213 8279 46229 8313
rect 46401 8279 46417 8313
rect 46585 8279 46601 8313
rect 46773 8279 46789 8313
rect 46957 8279 46973 8313
rect 47145 8279 47161 8313
rect 47329 8279 47345 8313
rect 47517 8279 47533 8313
rect 47701 8279 47717 8313
rect 47889 8279 47905 8313
rect 48073 8279 48089 8313
rect 48261 8279 48277 8313
rect 48445 8279 48461 8313
rect 48633 8279 48649 8313
rect 48817 8279 48833 8313
rect 49005 8279 49021 8313
rect 49189 8279 49205 8313
rect 49377 8279 49393 8313
rect 49561 8279 49577 8313
rect 49749 8279 49765 8313
rect 49933 8279 49949 8313
rect 50121 8279 50137 8313
rect 50305 8279 50321 8313
rect 50493 8279 50509 8313
rect 50677 8279 50693 8313
rect 50865 8279 50881 8313
rect 51049 8279 51065 8313
rect 39287 8220 39321 8236
rect 39287 7828 39321 7844
rect 39545 8220 39579 8236
rect 39545 7828 39579 7844
rect 39659 8220 39693 8236
rect 39659 7828 39693 7844
rect 39917 8220 39951 8236
rect 39917 7828 39951 7844
rect 40031 8220 40065 8236
rect 40031 7828 40065 7844
rect 40289 8220 40323 8236
rect 40289 7828 40323 7844
rect 40403 8220 40437 8236
rect 40403 7828 40437 7844
rect 40661 8220 40695 8236
rect 40661 7828 40695 7844
rect 40775 8220 40809 8236
rect 40775 7828 40809 7844
rect 41033 8220 41067 8236
rect 41033 7828 41067 7844
rect 41147 8220 41181 8236
rect 41147 7828 41181 7844
rect 41405 8220 41439 8236
rect 41405 7828 41439 7844
rect 41519 8220 41553 8236
rect 41519 7828 41553 7844
rect 41777 8220 41811 8236
rect 41777 7828 41811 7844
rect 41891 8220 41925 8236
rect 41891 7828 41925 7844
rect 42149 8220 42183 8236
rect 42149 7828 42183 7844
rect 42263 8220 42297 8236
rect 42263 7828 42297 7844
rect 42521 8220 42555 8236
rect 42521 7828 42555 7844
rect 42635 8220 42669 8236
rect 42635 7828 42669 7844
rect 42893 8220 42927 8236
rect 42893 7828 42927 7844
rect 43007 8220 43041 8236
rect 43007 7828 43041 7844
rect 43265 8220 43299 8236
rect 43265 7828 43299 7844
rect 43379 8220 43413 8236
rect 43379 7828 43413 7844
rect 43637 8220 43671 8236
rect 43637 7828 43671 7844
rect 43751 8220 43785 8236
rect 43751 7828 43785 7844
rect 44009 8220 44043 8236
rect 44009 7828 44043 7844
rect 44123 8220 44157 8236
rect 44123 7828 44157 7844
rect 44381 8220 44415 8236
rect 44381 7828 44415 7844
rect 44495 8220 44529 8236
rect 44495 7828 44529 7844
rect 44753 8220 44787 8236
rect 44753 7828 44787 7844
rect 44867 8220 44901 8236
rect 44867 7828 44901 7844
rect 45125 8220 45159 8236
rect 45125 7828 45159 7844
rect 45239 8220 45273 8236
rect 45239 7828 45273 7844
rect 45497 8220 45531 8236
rect 45497 7828 45531 7844
rect 45611 8220 45645 8236
rect 45611 7828 45645 7844
rect 45869 8220 45903 8236
rect 45869 7828 45903 7844
rect 45983 8220 46017 8236
rect 45983 7828 46017 7844
rect 46241 8220 46275 8236
rect 46241 7828 46275 7844
rect 46355 8220 46389 8236
rect 46355 7828 46389 7844
rect 46613 8220 46647 8236
rect 46613 7828 46647 7844
rect 46727 8220 46761 8236
rect 46727 7828 46761 7844
rect 46985 8220 47019 8236
rect 46985 7828 47019 7844
rect 47099 8220 47133 8236
rect 47099 7828 47133 7844
rect 47357 8220 47391 8236
rect 47357 7828 47391 7844
rect 47471 8220 47505 8236
rect 47471 7828 47505 7844
rect 47729 8220 47763 8236
rect 47729 7828 47763 7844
rect 47843 8220 47877 8236
rect 47843 7828 47877 7844
rect 48101 8220 48135 8236
rect 48101 7828 48135 7844
rect 48215 8220 48249 8236
rect 48215 7828 48249 7844
rect 48473 8220 48507 8236
rect 48473 7828 48507 7844
rect 48587 8220 48621 8236
rect 48587 7828 48621 7844
rect 48845 8220 48879 8236
rect 48845 7828 48879 7844
rect 48959 8220 48993 8236
rect 48959 7828 48993 7844
rect 49217 8220 49251 8236
rect 49217 7828 49251 7844
rect 49331 8220 49365 8236
rect 49331 7828 49365 7844
rect 49589 8220 49623 8236
rect 49589 7828 49623 7844
rect 49703 8220 49737 8236
rect 49703 7828 49737 7844
rect 49961 8220 49995 8236
rect 49961 7828 49995 7844
rect 50075 8220 50109 8236
rect 50075 7828 50109 7844
rect 50333 8220 50367 8236
rect 50333 7828 50367 7844
rect 50447 8220 50481 8236
rect 50447 7828 50481 7844
rect 50705 8220 50739 8236
rect 50705 7828 50739 7844
rect 50819 8220 50853 8236
rect 50819 7828 50853 7844
rect 51077 8220 51111 8236
rect 51077 7828 51111 7844
rect 39333 7751 39349 7785
rect 39517 7751 39533 7785
rect 39705 7751 39721 7785
rect 39889 7751 39905 7785
rect 40077 7751 40093 7785
rect 40261 7751 40277 7785
rect 40449 7751 40465 7785
rect 40633 7751 40649 7785
rect 40821 7751 40837 7785
rect 41005 7751 41021 7785
rect 41193 7751 41209 7785
rect 41377 7751 41393 7785
rect 41565 7751 41581 7785
rect 41749 7751 41765 7785
rect 41937 7751 41953 7785
rect 42121 7751 42137 7785
rect 42309 7751 42325 7785
rect 42493 7751 42509 7785
rect 42681 7751 42697 7785
rect 42865 7751 42881 7785
rect 43053 7751 43069 7785
rect 43237 7751 43253 7785
rect 43425 7751 43441 7785
rect 43609 7751 43625 7785
rect 43797 7751 43813 7785
rect 43981 7751 43997 7785
rect 44169 7751 44185 7785
rect 44353 7751 44369 7785
rect 44541 7751 44557 7785
rect 44725 7751 44741 7785
rect 44913 7751 44929 7785
rect 45097 7751 45113 7785
rect 45285 7751 45301 7785
rect 45469 7751 45485 7785
rect 45657 7751 45673 7785
rect 45841 7751 45857 7785
rect 46029 7751 46045 7785
rect 46213 7751 46229 7785
rect 46401 7751 46417 7785
rect 46585 7751 46601 7785
rect 46773 7751 46789 7785
rect 46957 7751 46973 7785
rect 47145 7751 47161 7785
rect 47329 7751 47345 7785
rect 47517 7751 47533 7785
rect 47701 7751 47717 7785
rect 47889 7751 47905 7785
rect 48073 7751 48089 7785
rect 48261 7751 48277 7785
rect 48445 7751 48461 7785
rect 48633 7751 48649 7785
rect 48817 7751 48833 7785
rect 49005 7751 49021 7785
rect 49189 7751 49205 7785
rect 49377 7751 49393 7785
rect 49561 7751 49577 7785
rect 49749 7751 49765 7785
rect 49933 7751 49949 7785
rect 50121 7751 50137 7785
rect 50305 7751 50321 7785
rect 50493 7751 50509 7785
rect 50677 7751 50693 7785
rect 50865 7751 50881 7785
rect 51049 7751 51065 7785
rect 39333 7643 39349 7677
rect 39517 7643 39533 7677
rect 39705 7643 39721 7677
rect 39889 7643 39905 7677
rect 40077 7643 40093 7677
rect 40261 7643 40277 7677
rect 40449 7643 40465 7677
rect 40633 7643 40649 7677
rect 40821 7643 40837 7677
rect 41005 7643 41021 7677
rect 41193 7643 41209 7677
rect 41377 7643 41393 7677
rect 41565 7643 41581 7677
rect 41749 7643 41765 7677
rect 41937 7643 41953 7677
rect 42121 7643 42137 7677
rect 42309 7643 42325 7677
rect 42493 7643 42509 7677
rect 42681 7643 42697 7677
rect 42865 7643 42881 7677
rect 43053 7643 43069 7677
rect 43237 7643 43253 7677
rect 43425 7643 43441 7677
rect 43609 7643 43625 7677
rect 43797 7643 43813 7677
rect 43981 7643 43997 7677
rect 44169 7643 44185 7677
rect 44353 7643 44369 7677
rect 44541 7643 44557 7677
rect 44725 7643 44741 7677
rect 44913 7643 44929 7677
rect 45097 7643 45113 7677
rect 45285 7643 45301 7677
rect 45469 7643 45485 7677
rect 45657 7643 45673 7677
rect 45841 7643 45857 7677
rect 46029 7643 46045 7677
rect 46213 7643 46229 7677
rect 46401 7643 46417 7677
rect 46585 7643 46601 7677
rect 46773 7643 46789 7677
rect 46957 7643 46973 7677
rect 47145 7643 47161 7677
rect 47329 7643 47345 7677
rect 47517 7643 47533 7677
rect 47701 7643 47717 7677
rect 47889 7643 47905 7677
rect 48073 7643 48089 7677
rect 48261 7643 48277 7677
rect 48445 7643 48461 7677
rect 48633 7643 48649 7677
rect 48817 7643 48833 7677
rect 49005 7643 49021 7677
rect 49189 7643 49205 7677
rect 49377 7643 49393 7677
rect 49561 7643 49577 7677
rect 49749 7643 49765 7677
rect 49933 7643 49949 7677
rect 50121 7643 50137 7677
rect 50305 7643 50321 7677
rect 50493 7643 50509 7677
rect 50677 7643 50693 7677
rect 50865 7643 50881 7677
rect 51049 7643 51065 7677
rect 39287 7584 39321 7600
rect 39287 7192 39321 7208
rect 39545 7584 39579 7600
rect 39545 7192 39579 7208
rect 39659 7584 39693 7600
rect 39659 7192 39693 7208
rect 39917 7584 39951 7600
rect 39917 7192 39951 7208
rect 40031 7584 40065 7600
rect 40031 7192 40065 7208
rect 40289 7584 40323 7600
rect 40289 7192 40323 7208
rect 40403 7584 40437 7600
rect 40403 7192 40437 7208
rect 40661 7584 40695 7600
rect 40661 7192 40695 7208
rect 40775 7584 40809 7600
rect 40775 7192 40809 7208
rect 41033 7584 41067 7600
rect 41033 7192 41067 7208
rect 41147 7584 41181 7600
rect 41147 7192 41181 7208
rect 41405 7584 41439 7600
rect 41405 7192 41439 7208
rect 41519 7584 41553 7600
rect 41519 7192 41553 7208
rect 41777 7584 41811 7600
rect 41777 7192 41811 7208
rect 41891 7584 41925 7600
rect 41891 7192 41925 7208
rect 42149 7584 42183 7600
rect 42149 7192 42183 7208
rect 42263 7584 42297 7600
rect 42263 7192 42297 7208
rect 42521 7584 42555 7600
rect 42521 7192 42555 7208
rect 42635 7584 42669 7600
rect 42635 7192 42669 7208
rect 42893 7584 42927 7600
rect 42893 7192 42927 7208
rect 43007 7584 43041 7600
rect 43007 7192 43041 7208
rect 43265 7584 43299 7600
rect 43265 7192 43299 7208
rect 43379 7584 43413 7600
rect 43379 7192 43413 7208
rect 43637 7584 43671 7600
rect 43637 7192 43671 7208
rect 43751 7584 43785 7600
rect 43751 7192 43785 7208
rect 44009 7584 44043 7600
rect 44009 7192 44043 7208
rect 44123 7584 44157 7600
rect 44123 7192 44157 7208
rect 44381 7584 44415 7600
rect 44381 7192 44415 7208
rect 44495 7584 44529 7600
rect 44495 7192 44529 7208
rect 44753 7584 44787 7600
rect 44753 7192 44787 7208
rect 44867 7584 44901 7600
rect 44867 7192 44901 7208
rect 45125 7584 45159 7600
rect 45125 7192 45159 7208
rect 45239 7584 45273 7600
rect 45239 7192 45273 7208
rect 45497 7584 45531 7600
rect 45497 7192 45531 7208
rect 45611 7584 45645 7600
rect 45611 7192 45645 7208
rect 45869 7584 45903 7600
rect 45869 7192 45903 7208
rect 45983 7584 46017 7600
rect 45983 7192 46017 7208
rect 46241 7584 46275 7600
rect 46241 7192 46275 7208
rect 46355 7584 46389 7600
rect 46355 7192 46389 7208
rect 46613 7584 46647 7600
rect 46613 7192 46647 7208
rect 46727 7584 46761 7600
rect 46727 7192 46761 7208
rect 46985 7584 47019 7600
rect 46985 7192 47019 7208
rect 47099 7584 47133 7600
rect 47099 7192 47133 7208
rect 47357 7584 47391 7600
rect 47357 7192 47391 7208
rect 47471 7584 47505 7600
rect 47471 7192 47505 7208
rect 47729 7584 47763 7600
rect 47729 7192 47763 7208
rect 47843 7584 47877 7600
rect 47843 7192 47877 7208
rect 48101 7584 48135 7600
rect 48101 7192 48135 7208
rect 48215 7584 48249 7600
rect 48215 7192 48249 7208
rect 48473 7584 48507 7600
rect 48473 7192 48507 7208
rect 48587 7584 48621 7600
rect 48587 7192 48621 7208
rect 48845 7584 48879 7600
rect 48845 7192 48879 7208
rect 48959 7584 48993 7600
rect 48959 7192 48993 7208
rect 49217 7584 49251 7600
rect 49217 7192 49251 7208
rect 49331 7584 49365 7600
rect 49331 7192 49365 7208
rect 49589 7584 49623 7600
rect 49589 7192 49623 7208
rect 49703 7584 49737 7600
rect 49703 7192 49737 7208
rect 49961 7584 49995 7600
rect 49961 7192 49995 7208
rect 50075 7584 50109 7600
rect 50075 7192 50109 7208
rect 50333 7584 50367 7600
rect 50333 7192 50367 7208
rect 50447 7584 50481 7600
rect 50447 7192 50481 7208
rect 50705 7584 50739 7600
rect 50705 7192 50739 7208
rect 50819 7584 50853 7600
rect 50819 7192 50853 7208
rect 51077 7584 51111 7600
rect 51077 7192 51111 7208
rect 39333 7115 39349 7149
rect 39517 7115 39533 7149
rect 39705 7115 39721 7149
rect 39889 7115 39905 7149
rect 40077 7115 40093 7149
rect 40261 7115 40277 7149
rect 40449 7115 40465 7149
rect 40633 7115 40649 7149
rect 40821 7115 40837 7149
rect 41005 7115 41021 7149
rect 41193 7115 41209 7149
rect 41377 7115 41393 7149
rect 41565 7115 41581 7149
rect 41749 7115 41765 7149
rect 41937 7115 41953 7149
rect 42121 7115 42137 7149
rect 42309 7115 42325 7149
rect 42493 7115 42509 7149
rect 42681 7115 42697 7149
rect 42865 7115 42881 7149
rect 43053 7115 43069 7149
rect 43237 7115 43253 7149
rect 43425 7115 43441 7149
rect 43609 7115 43625 7149
rect 43797 7115 43813 7149
rect 43981 7115 43997 7149
rect 44169 7115 44185 7149
rect 44353 7115 44369 7149
rect 44541 7115 44557 7149
rect 44725 7115 44741 7149
rect 44913 7115 44929 7149
rect 45097 7115 45113 7149
rect 45285 7115 45301 7149
rect 45469 7115 45485 7149
rect 45657 7115 45673 7149
rect 45841 7115 45857 7149
rect 46029 7115 46045 7149
rect 46213 7115 46229 7149
rect 46401 7115 46417 7149
rect 46585 7115 46601 7149
rect 46773 7115 46789 7149
rect 46957 7115 46973 7149
rect 47145 7115 47161 7149
rect 47329 7115 47345 7149
rect 47517 7115 47533 7149
rect 47701 7115 47717 7149
rect 47889 7115 47905 7149
rect 48073 7115 48089 7149
rect 48261 7115 48277 7149
rect 48445 7115 48461 7149
rect 48633 7115 48649 7149
rect 48817 7115 48833 7149
rect 49005 7115 49021 7149
rect 49189 7115 49205 7149
rect 49377 7115 49393 7149
rect 49561 7115 49577 7149
rect 49749 7115 49765 7149
rect 49933 7115 49949 7149
rect 50121 7115 50137 7149
rect 50305 7115 50321 7149
rect 50493 7115 50509 7149
rect 50677 7115 50693 7149
rect 50865 7115 50881 7149
rect 51049 7115 51065 7149
rect 39173 7047 39207 7109
rect 51191 7047 51225 7109
rect 39173 7013 39269 7047
rect 51129 7013 51225 7047
rect 39375 6836 39471 6870
rect 39927 6836 40023 6870
rect 39375 6774 39409 6836
rect 39989 6774 40023 6836
rect 40661 6629 40746 6663
rect 43689 6629 43785 6663
rect 40661 6567 40695 6629
rect 39375 4780 39409 4842
rect 39989 4780 40023 4842
rect 39375 4746 39471 4780
rect 39927 4746 40023 4780
rect 43751 6567 43785 6629
rect 40821 6527 40837 6561
rect 41005 6527 41021 6561
rect 41193 6527 41209 6561
rect 41377 6527 41393 6561
rect 41565 6527 41581 6561
rect 41749 6527 41765 6561
rect 41937 6527 41953 6561
rect 42121 6527 42137 6561
rect 42309 6527 42325 6561
rect 42493 6527 42509 6561
rect 42681 6527 42697 6561
rect 42865 6527 42881 6561
rect 43053 6527 43069 6561
rect 43237 6527 43253 6561
rect 43425 6527 43441 6561
rect 43609 6527 43625 6561
rect 40775 6468 40809 6484
rect 40775 5676 40809 5692
rect 41033 6468 41067 6484
rect 41033 5676 41067 5692
rect 41147 6468 41181 6484
rect 41147 5676 41181 5692
rect 41405 6468 41439 6484
rect 41405 5676 41439 5692
rect 41519 6468 41553 6484
rect 41519 5676 41553 5692
rect 41777 6468 41811 6484
rect 41777 5676 41811 5692
rect 41891 6468 41925 6484
rect 41891 5676 41925 5692
rect 42149 6468 42183 6484
rect 42149 5676 42183 5692
rect 42263 6468 42297 6484
rect 42263 5676 42297 5692
rect 42521 6468 42555 6484
rect 42521 5676 42555 5692
rect 42635 6468 42669 6484
rect 42635 5676 42669 5692
rect 42893 6468 42927 6484
rect 42893 5676 42927 5692
rect 43007 6468 43041 6484
rect 43007 5676 43041 5692
rect 43265 6468 43299 6484
rect 43265 5676 43299 5692
rect 43379 6468 43413 6484
rect 43379 5676 43413 5692
rect 43637 6468 43671 6484
rect 43637 5676 43671 5692
rect 40821 5599 40837 5633
rect 41005 5599 41021 5633
rect 41193 5599 41209 5633
rect 41377 5599 41393 5633
rect 41565 5599 41581 5633
rect 41749 5599 41765 5633
rect 41937 5599 41953 5633
rect 42121 5599 42137 5633
rect 42309 5599 42325 5633
rect 42493 5599 42509 5633
rect 42681 5599 42697 5633
rect 42865 5599 42881 5633
rect 43053 5599 43069 5633
rect 43237 5599 43253 5633
rect 43425 5599 43441 5633
rect 43609 5599 43625 5633
rect 40821 5491 40837 5525
rect 41005 5491 41021 5525
rect 41193 5491 41209 5525
rect 41377 5491 41393 5525
rect 41565 5491 41581 5525
rect 41749 5491 41765 5525
rect 41937 5491 41953 5525
rect 42121 5491 42137 5525
rect 42309 5491 42325 5525
rect 42493 5491 42509 5525
rect 42681 5491 42697 5525
rect 42865 5491 42881 5525
rect 43053 5491 43069 5525
rect 43237 5491 43253 5525
rect 43425 5491 43441 5525
rect 43609 5491 43625 5525
rect 40775 5432 40809 5448
rect 40775 4640 40809 4656
rect 41033 5432 41067 5448
rect 41033 4640 41067 4656
rect 41147 5432 41181 5448
rect 41147 4640 41181 4656
rect 41405 5432 41439 5448
rect 41405 4640 41439 4656
rect 41519 5432 41553 5448
rect 41519 4640 41553 4656
rect 41777 5432 41811 5448
rect 41777 4640 41811 4656
rect 41891 5432 41925 5448
rect 41891 4640 41925 4656
rect 42149 5432 42183 5448
rect 42149 4640 42183 4656
rect 42263 5432 42297 5448
rect 42263 4640 42297 4656
rect 42521 5432 42555 5448
rect 42521 4640 42555 4656
rect 42635 5432 42669 5448
rect 42635 4640 42669 4656
rect 42893 5432 42927 5448
rect 42893 4640 42927 4656
rect 43007 5432 43041 5448
rect 43007 4640 43041 4656
rect 43265 5432 43299 5448
rect 43265 4640 43299 4656
rect 43379 5432 43413 5448
rect 43379 4640 43413 4656
rect 43637 5432 43671 5448
rect 43637 4640 43671 4656
rect 40821 4563 40837 4597
rect 41005 4563 41021 4597
rect 41193 4563 41209 4597
rect 41377 4563 41393 4597
rect 41565 4563 41581 4597
rect 41749 4563 41765 4597
rect 41937 4563 41953 4597
rect 42121 4563 42137 4597
rect 42309 4563 42325 4597
rect 42493 4563 42509 4597
rect 42681 4563 42697 4597
rect 42865 4563 42881 4597
rect 43053 4563 43069 4597
rect 43237 4563 43253 4597
rect 43425 4563 43441 4597
rect 43609 4563 43625 4597
rect 40821 4455 40837 4489
rect 41005 4455 41021 4489
rect 41193 4455 41209 4489
rect 41377 4455 41393 4489
rect 41565 4455 41581 4489
rect 41749 4455 41765 4489
rect 41937 4455 41953 4489
rect 42121 4455 42137 4489
rect 42309 4455 42325 4489
rect 42493 4455 42509 4489
rect 42681 4455 42697 4489
rect 42865 4455 42881 4489
rect 43053 4455 43069 4489
rect 43237 4455 43253 4489
rect 43425 4455 43441 4489
rect 43609 4455 43625 4489
rect 40775 4396 40809 4412
rect 40775 3604 40809 3620
rect 41033 4396 41067 4412
rect 41033 3604 41067 3620
rect 41147 4396 41181 4412
rect 41147 3604 41181 3620
rect 41405 4396 41439 4412
rect 41405 3604 41439 3620
rect 41519 4396 41553 4412
rect 41519 3604 41553 3620
rect 41777 4396 41811 4412
rect 41777 3604 41811 3620
rect 41891 4396 41925 4412
rect 41891 3604 41925 3620
rect 42149 4396 42183 4412
rect 42149 3604 42183 3620
rect 42263 4396 42297 4412
rect 42263 3604 42297 3620
rect 42521 4396 42555 4412
rect 42521 3604 42555 3620
rect 42635 4396 42669 4412
rect 42635 3604 42669 3620
rect 42893 4396 42927 4412
rect 42893 3604 42927 3620
rect 43007 4396 43041 4412
rect 43007 3604 43041 3620
rect 43265 4396 43299 4412
rect 43265 3604 43299 3620
rect 43379 4396 43413 4412
rect 43379 3604 43413 3620
rect 43637 4396 43671 4412
rect 43637 3604 43671 3620
rect 40821 3527 40837 3561
rect 41005 3527 41021 3561
rect 41193 3527 41209 3561
rect 41377 3527 41393 3561
rect 41565 3527 41581 3561
rect 41749 3527 41765 3561
rect 41937 3527 41953 3561
rect 42121 3527 42137 3561
rect 42309 3527 42325 3561
rect 42493 3527 42509 3561
rect 42681 3527 42697 3561
rect 42865 3527 42881 3561
rect 43053 3527 43069 3561
rect 43237 3527 43253 3561
rect 43425 3527 43441 3561
rect 43609 3527 43625 3561
rect 40821 3419 40837 3453
rect 41005 3419 41021 3453
rect 41193 3419 41209 3453
rect 41377 3419 41393 3453
rect 41565 3419 41581 3453
rect 41749 3419 41765 3453
rect 41937 3419 41953 3453
rect 42121 3419 42137 3453
rect 42309 3419 42325 3453
rect 42493 3419 42509 3453
rect 42681 3419 42697 3453
rect 42865 3419 42881 3453
rect 43053 3419 43069 3453
rect 43237 3419 43253 3453
rect 43425 3419 43441 3453
rect 43609 3419 43625 3453
rect 40775 3360 40809 3376
rect 40775 2568 40809 2584
rect 41033 3360 41067 3376
rect 41033 2568 41067 2584
rect 41147 3360 41181 3376
rect 41147 2568 41181 2584
rect 41405 3360 41439 3376
rect 41405 2568 41439 2584
rect 41519 3360 41553 3376
rect 41519 2568 41553 2584
rect 41777 3360 41811 3376
rect 41777 2568 41811 2584
rect 41891 3360 41925 3376
rect 41891 2568 41925 2584
rect 42149 3360 42183 3376
rect 42149 2568 42183 2584
rect 42263 3360 42297 3376
rect 42263 2568 42297 2584
rect 42521 3360 42555 3376
rect 42521 2568 42555 2584
rect 42635 3360 42669 3376
rect 42635 2568 42669 2584
rect 42893 3360 42927 3376
rect 42893 2568 42927 2584
rect 43007 3360 43041 3376
rect 43007 2568 43041 2584
rect 43265 3360 43299 3376
rect 43265 2568 43299 2584
rect 43379 3360 43413 3376
rect 43379 2568 43413 2584
rect 43637 3360 43671 3376
rect 43637 2568 43671 2584
rect 40821 2491 40837 2525
rect 41005 2491 41021 2525
rect 41193 2491 41209 2525
rect 41377 2491 41393 2525
rect 41565 2491 41581 2525
rect 41749 2491 41765 2525
rect 41937 2491 41953 2525
rect 42121 2491 42137 2525
rect 42309 2491 42325 2525
rect 42493 2491 42509 2525
rect 42681 2491 42697 2525
rect 42865 2491 42881 2525
rect 43053 2491 43069 2525
rect 43237 2491 43253 2525
rect 43425 2491 43441 2525
rect 43609 2491 43625 2525
rect 40661 2423 40695 2485
rect 44531 6196 44627 6230
rect 45083 6196 45179 6230
rect 44531 6134 44565 6196
rect 45145 6134 45179 6196
rect 44531 4140 44565 4202
rect 45825 4473 45921 4507
rect 46059 4473 46155 4507
rect 45825 4411 45859 4473
rect 46121 4411 46155 4473
rect 45145 4140 45179 4202
rect 44531 4106 44627 4140
rect 45083 4106 45179 4140
rect 45825 3317 45859 3379
rect 46121 3317 46155 3379
rect 45825 3283 45921 3317
rect 46059 3283 46155 3317
rect 43751 2423 43785 2485
rect 40661 2389 40757 2423
rect 43689 2389 43785 2423
rect 40661 1935 40757 1969
rect 49641 1935 49737 1969
rect 40661 1873 40695 1935
rect 49703 1873 49737 1935
rect 40821 1833 40837 1867
rect 41005 1833 41021 1867
rect 41193 1833 41209 1867
rect 41377 1833 41393 1867
rect 41565 1833 41581 1867
rect 41749 1833 41765 1867
rect 41937 1833 41953 1867
rect 42121 1833 42137 1867
rect 42309 1833 42325 1867
rect 42493 1833 42509 1867
rect 42681 1833 42697 1867
rect 42865 1833 42881 1867
rect 43053 1833 43069 1867
rect 43237 1833 43253 1867
rect 43425 1833 43441 1867
rect 43609 1833 43625 1867
rect 43797 1833 43813 1867
rect 43981 1833 43997 1867
rect 44169 1833 44185 1867
rect 44353 1833 44369 1867
rect 44541 1833 44557 1867
rect 44725 1833 44741 1867
rect 44913 1833 44929 1867
rect 45097 1833 45113 1867
rect 45285 1833 45301 1867
rect 45469 1833 45485 1867
rect 45657 1833 45673 1867
rect 45841 1833 45857 1867
rect 46029 1833 46045 1867
rect 46213 1833 46229 1867
rect 46401 1833 46417 1867
rect 46585 1833 46601 1867
rect 46773 1833 46789 1867
rect 46957 1833 46973 1867
rect 47145 1833 47161 1867
rect 47329 1833 47345 1867
rect 47517 1833 47533 1867
rect 47701 1833 47717 1867
rect 47889 1833 47905 1867
rect 48073 1833 48089 1867
rect 48261 1833 48277 1867
rect 48445 1833 48461 1867
rect 48633 1833 48649 1867
rect 48817 1833 48833 1867
rect 49005 1833 49021 1867
rect 49189 1833 49205 1867
rect 49377 1833 49393 1867
rect 49561 1833 49577 1867
rect 40775 1783 40809 1799
rect 40775 1591 40809 1607
rect 41033 1783 41067 1799
rect 41033 1591 41067 1607
rect 41147 1783 41181 1799
rect 41147 1591 41181 1607
rect 41405 1783 41439 1799
rect 41405 1591 41439 1607
rect 41519 1783 41553 1799
rect 41519 1591 41553 1607
rect 41777 1783 41811 1799
rect 41777 1591 41811 1607
rect 41891 1783 41925 1799
rect 41891 1591 41925 1607
rect 42149 1783 42183 1799
rect 42149 1591 42183 1607
rect 42263 1783 42297 1799
rect 42263 1591 42297 1607
rect 42521 1783 42555 1799
rect 42521 1591 42555 1607
rect 42635 1783 42669 1799
rect 42635 1591 42669 1607
rect 42893 1783 42927 1799
rect 42893 1591 42927 1607
rect 43007 1783 43041 1799
rect 43007 1591 43041 1607
rect 43265 1783 43299 1799
rect 43265 1591 43299 1607
rect 43379 1783 43413 1799
rect 43379 1591 43413 1607
rect 43637 1783 43671 1799
rect 43637 1591 43671 1607
rect 43751 1783 43785 1799
rect 43751 1591 43785 1607
rect 44009 1783 44043 1799
rect 44009 1591 44043 1607
rect 44123 1783 44157 1799
rect 44123 1591 44157 1607
rect 44381 1783 44415 1799
rect 44381 1591 44415 1607
rect 44495 1783 44529 1799
rect 44495 1591 44529 1607
rect 44753 1783 44787 1799
rect 44753 1591 44787 1607
rect 44867 1783 44901 1799
rect 44867 1591 44901 1607
rect 45125 1783 45159 1799
rect 45125 1591 45159 1607
rect 45239 1783 45273 1799
rect 45239 1591 45273 1607
rect 45497 1783 45531 1799
rect 45497 1591 45531 1607
rect 45611 1783 45645 1799
rect 45611 1591 45645 1607
rect 45869 1783 45903 1799
rect 45869 1591 45903 1607
rect 45983 1783 46017 1799
rect 45983 1591 46017 1607
rect 46241 1783 46275 1799
rect 46241 1591 46275 1607
rect 46355 1783 46389 1799
rect 46355 1591 46389 1607
rect 46613 1783 46647 1799
rect 46613 1591 46647 1607
rect 46727 1783 46761 1799
rect 46727 1591 46761 1607
rect 46985 1783 47019 1799
rect 46985 1591 47019 1607
rect 47099 1783 47133 1799
rect 47099 1591 47133 1607
rect 47357 1783 47391 1799
rect 47357 1591 47391 1607
rect 47471 1783 47505 1799
rect 47471 1591 47505 1607
rect 47729 1783 47763 1799
rect 47729 1591 47763 1607
rect 47843 1783 47877 1799
rect 47843 1591 47877 1607
rect 48101 1783 48135 1799
rect 48101 1591 48135 1607
rect 48215 1783 48249 1799
rect 48215 1591 48249 1607
rect 48473 1783 48507 1799
rect 48473 1591 48507 1607
rect 48587 1783 48621 1799
rect 48587 1591 48621 1607
rect 48845 1783 48879 1799
rect 48845 1591 48879 1607
rect 48959 1783 48993 1799
rect 48959 1591 48993 1607
rect 49217 1783 49251 1799
rect 49217 1591 49251 1607
rect 49331 1783 49365 1799
rect 49331 1591 49365 1607
rect 49589 1783 49623 1799
rect 49589 1591 49623 1607
rect 40821 1523 40837 1557
rect 41005 1523 41021 1557
rect 41193 1523 41209 1557
rect 41377 1523 41393 1557
rect 41565 1523 41581 1557
rect 41749 1523 41765 1557
rect 41937 1523 41953 1557
rect 42121 1523 42137 1557
rect 42309 1523 42325 1557
rect 42493 1523 42509 1557
rect 42681 1523 42697 1557
rect 42865 1523 42881 1557
rect 43053 1523 43069 1557
rect 43237 1523 43253 1557
rect 43425 1523 43441 1557
rect 43609 1523 43625 1557
rect 43797 1523 43813 1557
rect 43981 1523 43997 1557
rect 44169 1523 44185 1557
rect 44353 1523 44369 1557
rect 44541 1523 44557 1557
rect 44725 1523 44741 1557
rect 44913 1523 44929 1557
rect 45097 1523 45113 1557
rect 45285 1523 45301 1557
rect 45469 1523 45485 1557
rect 45657 1523 45673 1557
rect 45841 1523 45857 1557
rect 46029 1523 46045 1557
rect 46213 1523 46229 1557
rect 46401 1523 46417 1557
rect 46585 1523 46601 1557
rect 46773 1523 46789 1557
rect 46957 1523 46973 1557
rect 47145 1523 47161 1557
rect 47329 1523 47345 1557
rect 47517 1523 47533 1557
rect 47701 1523 47717 1557
rect 47889 1523 47905 1557
rect 48073 1523 48089 1557
rect 48261 1523 48277 1557
rect 48445 1523 48461 1557
rect 48633 1523 48649 1557
rect 48817 1523 48833 1557
rect 49005 1523 49021 1557
rect 49189 1523 49205 1557
rect 49377 1523 49393 1557
rect 49561 1523 49577 1557
rect 40821 1415 40837 1449
rect 41005 1415 41021 1449
rect 41193 1415 41209 1449
rect 41377 1415 41393 1449
rect 41565 1415 41581 1449
rect 41749 1415 41765 1449
rect 41937 1415 41953 1449
rect 42121 1415 42137 1449
rect 42309 1415 42325 1449
rect 42493 1415 42509 1449
rect 42681 1415 42697 1449
rect 42865 1415 42881 1449
rect 43053 1415 43069 1449
rect 43237 1415 43253 1449
rect 43425 1415 43441 1449
rect 43609 1415 43625 1449
rect 43797 1415 43813 1449
rect 43981 1415 43997 1449
rect 44169 1415 44185 1449
rect 44353 1415 44369 1449
rect 44541 1415 44557 1449
rect 44725 1415 44741 1449
rect 44913 1415 44929 1449
rect 45097 1415 45113 1449
rect 45285 1415 45301 1449
rect 45469 1415 45485 1449
rect 45657 1415 45673 1449
rect 45841 1415 45857 1449
rect 46029 1415 46045 1449
rect 46213 1415 46229 1449
rect 46401 1415 46417 1449
rect 46585 1415 46601 1449
rect 46773 1415 46789 1449
rect 46957 1415 46973 1449
rect 47145 1415 47161 1449
rect 47329 1415 47345 1449
rect 47517 1415 47533 1449
rect 47701 1415 47717 1449
rect 47889 1415 47905 1449
rect 48073 1415 48089 1449
rect 48261 1415 48277 1449
rect 48445 1415 48461 1449
rect 48633 1415 48649 1449
rect 48817 1415 48833 1449
rect 49005 1415 49021 1449
rect 49189 1415 49205 1449
rect 49377 1415 49393 1449
rect 49561 1415 49577 1449
rect 40775 1365 40809 1381
rect 40775 1173 40809 1189
rect 41033 1365 41067 1381
rect 41033 1173 41067 1189
rect 41147 1365 41181 1381
rect 41147 1173 41181 1189
rect 41405 1365 41439 1381
rect 41405 1173 41439 1189
rect 41519 1365 41553 1381
rect 41519 1173 41553 1189
rect 41777 1365 41811 1381
rect 41777 1173 41811 1189
rect 41891 1365 41925 1381
rect 41891 1173 41925 1189
rect 42149 1365 42183 1381
rect 42149 1173 42183 1189
rect 42263 1365 42297 1381
rect 42263 1173 42297 1189
rect 42521 1365 42555 1381
rect 42521 1173 42555 1189
rect 42635 1365 42669 1381
rect 42635 1173 42669 1189
rect 42893 1365 42927 1381
rect 42893 1173 42927 1189
rect 43007 1365 43041 1381
rect 43007 1173 43041 1189
rect 43265 1365 43299 1381
rect 43265 1173 43299 1189
rect 43379 1365 43413 1381
rect 43379 1173 43413 1189
rect 43637 1365 43671 1381
rect 43637 1173 43671 1189
rect 43751 1365 43785 1381
rect 43751 1173 43785 1189
rect 44009 1365 44043 1381
rect 44009 1173 44043 1189
rect 44123 1365 44157 1381
rect 44123 1173 44157 1189
rect 44381 1365 44415 1381
rect 44381 1173 44415 1189
rect 44495 1365 44529 1381
rect 44495 1173 44529 1189
rect 44753 1365 44787 1381
rect 44753 1173 44787 1189
rect 44867 1365 44901 1381
rect 44867 1173 44901 1189
rect 45125 1365 45159 1381
rect 45125 1173 45159 1189
rect 45239 1365 45273 1381
rect 45239 1173 45273 1189
rect 45497 1365 45531 1381
rect 45497 1173 45531 1189
rect 45611 1365 45645 1381
rect 45611 1173 45645 1189
rect 45869 1365 45903 1381
rect 45869 1173 45903 1189
rect 45983 1365 46017 1381
rect 45983 1173 46017 1189
rect 46241 1365 46275 1381
rect 46241 1173 46275 1189
rect 46355 1365 46389 1381
rect 46355 1173 46389 1189
rect 46613 1365 46647 1381
rect 46613 1173 46647 1189
rect 46727 1365 46761 1381
rect 46727 1173 46761 1189
rect 46985 1365 47019 1381
rect 46985 1173 47019 1189
rect 47099 1365 47133 1381
rect 47099 1173 47133 1189
rect 47357 1365 47391 1381
rect 47357 1173 47391 1189
rect 47471 1365 47505 1381
rect 47471 1173 47505 1189
rect 47729 1365 47763 1381
rect 47729 1173 47763 1189
rect 47843 1365 47877 1381
rect 47843 1173 47877 1189
rect 48101 1365 48135 1381
rect 48101 1173 48135 1189
rect 48215 1365 48249 1381
rect 48215 1173 48249 1189
rect 48473 1365 48507 1381
rect 48473 1173 48507 1189
rect 48587 1365 48621 1381
rect 48587 1173 48621 1189
rect 48845 1365 48879 1381
rect 48845 1173 48879 1189
rect 48959 1365 48993 1381
rect 48959 1173 48993 1189
rect 49217 1365 49251 1381
rect 49217 1173 49251 1189
rect 49331 1365 49365 1381
rect 49331 1173 49365 1189
rect 49589 1365 49623 1381
rect 49589 1173 49623 1189
rect 40821 1105 40837 1139
rect 41005 1105 41021 1139
rect 41193 1105 41209 1139
rect 41377 1105 41393 1139
rect 41565 1105 41581 1139
rect 41749 1105 41765 1139
rect 41937 1105 41953 1139
rect 42121 1105 42137 1139
rect 42309 1105 42325 1139
rect 42493 1105 42509 1139
rect 42681 1105 42697 1139
rect 42865 1105 42881 1139
rect 43053 1105 43069 1139
rect 43237 1105 43253 1139
rect 43425 1105 43441 1139
rect 43609 1105 43625 1139
rect 43797 1105 43813 1139
rect 43981 1105 43997 1139
rect 44169 1105 44185 1139
rect 44353 1105 44369 1139
rect 44541 1105 44557 1139
rect 44725 1105 44741 1139
rect 44913 1105 44929 1139
rect 45097 1105 45113 1139
rect 45285 1105 45301 1139
rect 45469 1105 45485 1139
rect 45657 1105 45673 1139
rect 45841 1105 45857 1139
rect 46029 1105 46045 1139
rect 46213 1105 46229 1139
rect 46401 1105 46417 1139
rect 46585 1105 46601 1139
rect 46773 1105 46789 1139
rect 46957 1105 46973 1139
rect 47145 1105 47161 1139
rect 47329 1105 47345 1139
rect 47517 1105 47533 1139
rect 47701 1105 47717 1139
rect 47889 1105 47905 1139
rect 48073 1105 48089 1139
rect 48261 1105 48277 1139
rect 48445 1105 48461 1139
rect 48633 1105 48649 1139
rect 48817 1105 48833 1139
rect 49005 1105 49021 1139
rect 49189 1105 49205 1139
rect 49377 1105 49393 1139
rect 49561 1105 49577 1139
rect 40821 997 40837 1031
rect 41005 997 41021 1031
rect 41193 997 41209 1031
rect 41377 997 41393 1031
rect 41565 997 41581 1031
rect 41749 997 41765 1031
rect 41937 997 41953 1031
rect 42121 997 42137 1031
rect 42309 997 42325 1031
rect 42493 997 42509 1031
rect 42681 997 42697 1031
rect 42865 997 42881 1031
rect 43053 997 43069 1031
rect 43237 997 43253 1031
rect 43425 997 43441 1031
rect 43609 997 43625 1031
rect 43797 997 43813 1031
rect 43981 997 43997 1031
rect 44169 997 44185 1031
rect 44353 997 44369 1031
rect 44541 997 44557 1031
rect 44725 997 44741 1031
rect 44913 997 44929 1031
rect 45097 997 45113 1031
rect 45285 997 45301 1031
rect 45469 997 45485 1031
rect 45657 997 45673 1031
rect 45841 997 45857 1031
rect 46029 997 46045 1031
rect 46213 997 46229 1031
rect 46401 997 46417 1031
rect 46585 997 46601 1031
rect 46773 997 46789 1031
rect 46957 997 46973 1031
rect 47145 997 47161 1031
rect 47329 997 47345 1031
rect 47517 997 47533 1031
rect 47701 997 47717 1031
rect 47889 997 47905 1031
rect 48073 997 48089 1031
rect 48261 997 48277 1031
rect 48445 997 48461 1031
rect 48633 997 48649 1031
rect 48817 997 48833 1031
rect 49005 997 49021 1031
rect 49189 997 49205 1031
rect 49377 997 49393 1031
rect 49561 997 49577 1031
rect 40775 947 40809 963
rect 40775 755 40809 771
rect 41033 947 41067 963
rect 41033 755 41067 771
rect 41147 947 41181 963
rect 41147 755 41181 771
rect 41405 947 41439 963
rect 41405 755 41439 771
rect 41519 947 41553 963
rect 41519 755 41553 771
rect 41777 947 41811 963
rect 41777 755 41811 771
rect 41891 947 41925 963
rect 41891 755 41925 771
rect 42149 947 42183 963
rect 42149 755 42183 771
rect 42263 947 42297 963
rect 42263 755 42297 771
rect 42521 947 42555 963
rect 42521 755 42555 771
rect 42635 947 42669 963
rect 42635 755 42669 771
rect 42893 947 42927 963
rect 42893 755 42927 771
rect 43007 947 43041 963
rect 43007 755 43041 771
rect 43265 947 43299 963
rect 43265 755 43299 771
rect 43379 947 43413 963
rect 43379 755 43413 771
rect 43637 947 43671 963
rect 43637 755 43671 771
rect 43751 947 43785 963
rect 43751 755 43785 771
rect 44009 947 44043 963
rect 44009 755 44043 771
rect 44123 947 44157 963
rect 44123 755 44157 771
rect 44381 947 44415 963
rect 44381 755 44415 771
rect 44495 947 44529 963
rect 44495 755 44529 771
rect 44753 947 44787 963
rect 44753 755 44787 771
rect 44867 947 44901 963
rect 44867 755 44901 771
rect 45125 947 45159 963
rect 45125 755 45159 771
rect 45239 947 45273 963
rect 45239 755 45273 771
rect 45497 947 45531 963
rect 45497 755 45531 771
rect 45611 947 45645 963
rect 45611 755 45645 771
rect 45869 947 45903 963
rect 45869 755 45903 771
rect 45983 947 46017 963
rect 45983 755 46017 771
rect 46241 947 46275 963
rect 46241 755 46275 771
rect 46355 947 46389 963
rect 46355 755 46389 771
rect 46613 947 46647 963
rect 46613 755 46647 771
rect 46727 947 46761 963
rect 46727 755 46761 771
rect 46985 947 47019 963
rect 46985 755 47019 771
rect 47099 947 47133 963
rect 47099 755 47133 771
rect 47357 947 47391 963
rect 47357 755 47391 771
rect 47471 947 47505 963
rect 47471 755 47505 771
rect 47729 947 47763 963
rect 47729 755 47763 771
rect 47843 947 47877 963
rect 47843 755 47877 771
rect 48101 947 48135 963
rect 48101 755 48135 771
rect 48215 947 48249 963
rect 48215 755 48249 771
rect 48473 947 48507 963
rect 48473 755 48507 771
rect 48587 947 48621 963
rect 48587 755 48621 771
rect 48845 947 48879 963
rect 48845 755 48879 771
rect 48959 947 48993 963
rect 48959 755 48993 771
rect 49217 947 49251 963
rect 49217 755 49251 771
rect 49331 947 49365 963
rect 49331 755 49365 771
rect 49589 947 49623 963
rect 49589 755 49623 771
rect 40821 687 40837 721
rect 41005 687 41021 721
rect 41193 687 41209 721
rect 41377 687 41393 721
rect 41565 687 41581 721
rect 41749 687 41765 721
rect 41937 687 41953 721
rect 42121 687 42137 721
rect 42309 687 42325 721
rect 42493 687 42509 721
rect 42681 687 42697 721
rect 42865 687 42881 721
rect 43053 687 43069 721
rect 43237 687 43253 721
rect 43425 687 43441 721
rect 43609 687 43625 721
rect 43797 687 43813 721
rect 43981 687 43997 721
rect 44169 687 44185 721
rect 44353 687 44369 721
rect 44541 687 44557 721
rect 44725 687 44741 721
rect 44913 687 44929 721
rect 45097 687 45113 721
rect 45285 687 45301 721
rect 45469 687 45485 721
rect 45657 687 45673 721
rect 45841 687 45857 721
rect 46029 687 46045 721
rect 46213 687 46229 721
rect 46401 687 46417 721
rect 46585 687 46601 721
rect 46773 687 46789 721
rect 46957 687 46973 721
rect 47145 687 47161 721
rect 47329 687 47345 721
rect 47517 687 47533 721
rect 47701 687 47717 721
rect 47889 687 47905 721
rect 48073 687 48089 721
rect 48261 687 48277 721
rect 48445 687 48461 721
rect 48633 687 48649 721
rect 48817 687 48833 721
rect 49005 687 49021 721
rect 49189 687 49205 721
rect 49377 687 49393 721
rect 49561 687 49577 721
rect 40821 579 40837 613
rect 41005 579 41021 613
rect 41193 579 41209 613
rect 41377 579 41393 613
rect 41565 579 41581 613
rect 41749 579 41765 613
rect 41937 579 41953 613
rect 42121 579 42137 613
rect 42309 579 42325 613
rect 42493 579 42509 613
rect 42681 579 42697 613
rect 42865 579 42881 613
rect 43053 579 43069 613
rect 43237 579 43253 613
rect 43425 579 43441 613
rect 43609 579 43625 613
rect 43797 579 43813 613
rect 43981 579 43997 613
rect 44169 579 44185 613
rect 44353 579 44369 613
rect 44541 579 44557 613
rect 44725 579 44741 613
rect 44913 579 44929 613
rect 45097 579 45113 613
rect 45285 579 45301 613
rect 45469 579 45485 613
rect 45657 579 45673 613
rect 45841 579 45857 613
rect 46029 579 46045 613
rect 46213 579 46229 613
rect 46401 579 46417 613
rect 46585 579 46601 613
rect 46773 579 46789 613
rect 46957 579 46973 613
rect 47145 579 47161 613
rect 47329 579 47345 613
rect 47517 579 47533 613
rect 47701 579 47717 613
rect 47889 579 47905 613
rect 48073 579 48089 613
rect 48261 579 48277 613
rect 48445 579 48461 613
rect 48633 579 48649 613
rect 48817 579 48833 613
rect 49005 579 49021 613
rect 49189 579 49205 613
rect 49377 579 49393 613
rect 49561 579 49577 613
rect 40775 529 40809 545
rect 40775 337 40809 353
rect 41033 529 41067 545
rect 41033 337 41067 353
rect 41147 529 41181 545
rect 41147 337 41181 353
rect 41405 529 41439 545
rect 41405 337 41439 353
rect 41519 529 41553 545
rect 41519 337 41553 353
rect 41777 529 41811 545
rect 41777 337 41811 353
rect 41891 529 41925 545
rect 41891 337 41925 353
rect 42149 529 42183 545
rect 42149 337 42183 353
rect 42263 529 42297 545
rect 42263 337 42297 353
rect 42521 529 42555 545
rect 42521 337 42555 353
rect 42635 529 42669 545
rect 42635 337 42669 353
rect 42893 529 42927 545
rect 42893 337 42927 353
rect 43007 529 43041 545
rect 43007 337 43041 353
rect 43265 529 43299 545
rect 43265 337 43299 353
rect 43379 529 43413 545
rect 43379 337 43413 353
rect 43637 529 43671 545
rect 43637 337 43671 353
rect 43751 529 43785 545
rect 43751 337 43785 353
rect 44009 529 44043 545
rect 44009 337 44043 353
rect 44123 529 44157 545
rect 44123 337 44157 353
rect 44381 529 44415 545
rect 44381 337 44415 353
rect 44495 529 44529 545
rect 44495 337 44529 353
rect 44753 529 44787 545
rect 44753 337 44787 353
rect 44867 529 44901 545
rect 44867 337 44901 353
rect 45125 529 45159 545
rect 45125 337 45159 353
rect 45239 529 45273 545
rect 45239 337 45273 353
rect 45497 529 45531 545
rect 45497 337 45531 353
rect 45611 529 45645 545
rect 45611 337 45645 353
rect 45869 529 45903 545
rect 45869 337 45903 353
rect 45983 529 46017 545
rect 45983 337 46017 353
rect 46241 529 46275 545
rect 46241 337 46275 353
rect 46355 529 46389 545
rect 46355 337 46389 353
rect 46613 529 46647 545
rect 46613 337 46647 353
rect 46727 529 46761 545
rect 46727 337 46761 353
rect 46985 529 47019 545
rect 46985 337 47019 353
rect 47099 529 47133 545
rect 47099 337 47133 353
rect 47357 529 47391 545
rect 47357 337 47391 353
rect 47471 529 47505 545
rect 47471 337 47505 353
rect 47729 529 47763 545
rect 47729 337 47763 353
rect 47843 529 47877 545
rect 47843 337 47877 353
rect 48101 529 48135 545
rect 48101 337 48135 353
rect 48215 529 48249 545
rect 48215 337 48249 353
rect 48473 529 48507 545
rect 48473 337 48507 353
rect 48587 529 48621 545
rect 48587 337 48621 353
rect 48845 529 48879 545
rect 48845 337 48879 353
rect 48959 529 48993 545
rect 48959 337 48993 353
rect 49217 529 49251 545
rect 49217 337 49251 353
rect 49331 529 49365 545
rect 49331 337 49365 353
rect 49589 529 49623 545
rect 49589 337 49623 353
rect 40821 269 40837 303
rect 41005 269 41021 303
rect 41193 269 41209 303
rect 41377 269 41393 303
rect 41565 269 41581 303
rect 41749 269 41765 303
rect 41937 269 41953 303
rect 42121 269 42137 303
rect 42309 269 42325 303
rect 42493 269 42509 303
rect 42681 269 42697 303
rect 42865 269 42881 303
rect 43053 269 43069 303
rect 43237 269 43253 303
rect 43425 269 43441 303
rect 43609 269 43625 303
rect 43797 269 43813 303
rect 43981 269 43997 303
rect 44169 269 44185 303
rect 44353 269 44369 303
rect 44541 269 44557 303
rect 44725 269 44741 303
rect 44913 269 44929 303
rect 45097 269 45113 303
rect 45285 269 45301 303
rect 45469 269 45485 303
rect 45657 269 45673 303
rect 45841 269 45857 303
rect 46029 269 46045 303
rect 46213 269 46229 303
rect 46401 269 46417 303
rect 46585 269 46601 303
rect 46773 269 46789 303
rect 46957 269 46973 303
rect 47145 269 47161 303
rect 47329 269 47345 303
rect 47517 269 47533 303
rect 47701 269 47717 303
rect 47889 269 47905 303
rect 48073 269 48089 303
rect 48261 269 48277 303
rect 48445 269 48461 303
rect 48633 269 48649 303
rect 48817 269 48833 303
rect 49005 269 49021 303
rect 49189 269 49205 303
rect 49377 269 49393 303
rect 49561 269 49577 303
rect 40661 201 40695 263
rect 49703 201 49737 263
rect 40661 167 40757 201
rect 49641 167 49737 201
<< viali >>
rect 40776 19698 40846 19723
rect 41444 19698 41514 19715
rect 42188 19698 42258 19715
rect 42932 19698 43002 19715
rect 43676 19698 43746 19715
rect 44420 19698 44490 19715
rect 45164 19698 45234 19715
rect 45908 19698 45978 19715
rect 46652 19698 46722 19715
rect 47396 19698 47466 19715
rect 48140 19698 48210 19715
rect 48884 19698 48954 19715
rect 49546 19698 49616 19719
rect 40776 19664 40846 19698
rect 41444 19664 41514 19698
rect 42188 19664 42258 19698
rect 42932 19664 43002 19698
rect 43676 19664 43746 19698
rect 44420 19664 44490 19698
rect 45164 19664 45234 19698
rect 45908 19664 45978 19698
rect 46652 19664 46722 19698
rect 47396 19664 47466 19698
rect 48140 19664 48210 19698
rect 48884 19664 48954 19698
rect 49546 19664 49616 19698
rect 40776 19653 40846 19664
rect 41444 19645 41514 19664
rect 42188 19645 42258 19664
rect 42932 19645 43002 19664
rect 43676 19645 43746 19664
rect 44420 19645 44490 19664
rect 45164 19645 45234 19664
rect 45908 19645 45978 19664
rect 46652 19645 46722 19664
rect 47396 19645 47466 19664
rect 48140 19645 48210 19664
rect 48884 19645 48954 19664
rect 49546 19649 49616 19664
rect 40837 19562 41005 19596
rect 41209 19562 41377 19596
rect 41581 19562 41749 19596
rect 41953 19562 42121 19596
rect 42325 19562 42493 19596
rect 42697 19562 42865 19596
rect 43069 19562 43237 19596
rect 43441 19562 43609 19596
rect 43813 19562 43981 19596
rect 44185 19562 44353 19596
rect 44557 19562 44725 19596
rect 44929 19562 45097 19596
rect 45301 19562 45469 19596
rect 45673 19562 45841 19596
rect 46045 19562 46213 19596
rect 46417 19562 46585 19596
rect 46789 19562 46957 19596
rect 47161 19562 47329 19596
rect 47533 19562 47701 19596
rect 47905 19562 48073 19596
rect 48277 19562 48445 19596
rect 48649 19562 48817 19596
rect 49021 19562 49189 19596
rect 49393 19562 49561 19596
rect 40775 19336 40809 19512
rect 41033 19336 41067 19512
rect 41147 19336 41181 19512
rect 41405 19336 41439 19512
rect 41519 19336 41553 19512
rect 41777 19336 41811 19512
rect 41891 19336 41925 19512
rect 42149 19336 42183 19512
rect 42263 19336 42297 19512
rect 42521 19336 42555 19512
rect 42635 19336 42669 19512
rect 42893 19336 42927 19512
rect 43007 19336 43041 19512
rect 43265 19336 43299 19512
rect 43379 19336 43413 19512
rect 43637 19336 43671 19512
rect 43751 19336 43785 19512
rect 44009 19336 44043 19512
rect 44123 19336 44157 19512
rect 44381 19336 44415 19512
rect 44495 19336 44529 19512
rect 44753 19336 44787 19512
rect 44867 19336 44901 19512
rect 45125 19336 45159 19512
rect 45239 19336 45273 19512
rect 45497 19336 45531 19512
rect 45611 19336 45645 19512
rect 45869 19336 45903 19512
rect 45983 19336 46017 19512
rect 46241 19336 46275 19512
rect 46355 19336 46389 19512
rect 46613 19336 46647 19512
rect 46727 19336 46761 19512
rect 46985 19336 47019 19512
rect 47099 19336 47133 19512
rect 47357 19336 47391 19512
rect 47471 19336 47505 19512
rect 47729 19336 47763 19512
rect 47843 19336 47877 19512
rect 48101 19336 48135 19512
rect 48215 19336 48249 19512
rect 48473 19336 48507 19512
rect 48587 19336 48621 19512
rect 48845 19336 48879 19512
rect 48959 19336 48993 19512
rect 49217 19336 49251 19512
rect 49331 19336 49365 19512
rect 49589 19336 49623 19512
rect 40837 19252 41005 19286
rect 41209 19252 41377 19286
rect 41581 19252 41749 19286
rect 41953 19252 42121 19286
rect 42325 19252 42493 19286
rect 42697 19252 42865 19286
rect 43069 19252 43237 19286
rect 43441 19252 43609 19286
rect 43813 19252 43981 19286
rect 44185 19252 44353 19286
rect 44557 19252 44725 19286
rect 44929 19252 45097 19286
rect 45301 19252 45469 19286
rect 45673 19252 45841 19286
rect 46045 19252 46213 19286
rect 46417 19252 46585 19286
rect 46789 19252 46957 19286
rect 47161 19252 47329 19286
rect 47533 19252 47701 19286
rect 47905 19252 48073 19286
rect 48277 19252 48445 19286
rect 48649 19252 48817 19286
rect 49021 19252 49189 19286
rect 49393 19252 49561 19286
rect 40837 19144 41005 19178
rect 41209 19144 41377 19178
rect 41581 19144 41749 19178
rect 41953 19144 42121 19178
rect 42325 19144 42493 19178
rect 42697 19144 42865 19178
rect 43069 19144 43237 19178
rect 43441 19144 43609 19178
rect 43813 19144 43981 19178
rect 44185 19144 44353 19178
rect 44557 19144 44725 19178
rect 44929 19144 45097 19178
rect 45301 19144 45469 19178
rect 45673 19144 45841 19178
rect 46045 19144 46213 19178
rect 46417 19144 46585 19178
rect 46789 19144 46957 19178
rect 47161 19144 47329 19178
rect 47533 19144 47701 19178
rect 47905 19144 48073 19178
rect 48277 19144 48445 19178
rect 48649 19144 48817 19178
rect 49021 19144 49189 19178
rect 49393 19144 49561 19178
rect 40775 18918 40809 19094
rect 41033 18918 41067 19094
rect 41147 18918 41181 19094
rect 41405 18918 41439 19094
rect 41519 18918 41553 19094
rect 41777 18918 41811 19094
rect 41891 18918 41925 19094
rect 42149 18918 42183 19094
rect 42263 18918 42297 19094
rect 42521 18918 42555 19094
rect 42635 18918 42669 19094
rect 42893 18918 42927 19094
rect 43007 18918 43041 19094
rect 43265 18918 43299 19094
rect 43379 18918 43413 19094
rect 43637 18918 43671 19094
rect 43751 18918 43785 19094
rect 44009 18918 44043 19094
rect 44123 18918 44157 19094
rect 44381 18918 44415 19094
rect 44495 18918 44529 19094
rect 44753 18918 44787 19094
rect 44867 18918 44901 19094
rect 45125 18918 45159 19094
rect 45239 18918 45273 19094
rect 45497 18918 45531 19094
rect 45611 18918 45645 19094
rect 45869 18918 45903 19094
rect 45983 18918 46017 19094
rect 46241 18918 46275 19094
rect 46355 18918 46389 19094
rect 46613 18918 46647 19094
rect 46727 18918 46761 19094
rect 46985 18918 47019 19094
rect 47099 18918 47133 19094
rect 47357 18918 47391 19094
rect 47471 18918 47505 19094
rect 47729 18918 47763 19094
rect 47843 18918 47877 19094
rect 48101 18918 48135 19094
rect 48215 18918 48249 19094
rect 48473 18918 48507 19094
rect 48587 18918 48621 19094
rect 48845 18918 48879 19094
rect 48959 18918 48993 19094
rect 49217 18918 49251 19094
rect 49331 18918 49365 19094
rect 49589 18918 49623 19094
rect 40837 18834 41005 18868
rect 41209 18834 41377 18868
rect 41581 18834 41749 18868
rect 41953 18834 42121 18868
rect 42325 18834 42493 18868
rect 42697 18834 42865 18868
rect 43069 18834 43237 18868
rect 43441 18834 43609 18868
rect 43813 18834 43981 18868
rect 44185 18834 44353 18868
rect 44557 18834 44725 18868
rect 44929 18834 45097 18868
rect 45301 18834 45469 18868
rect 45673 18834 45841 18868
rect 46045 18834 46213 18868
rect 46417 18834 46585 18868
rect 46789 18834 46957 18868
rect 47161 18834 47329 18868
rect 47533 18834 47701 18868
rect 47905 18834 48073 18868
rect 48277 18834 48445 18868
rect 48649 18834 48817 18868
rect 49021 18834 49189 18868
rect 49393 18834 49561 18868
rect 40837 18726 41005 18760
rect 41209 18726 41377 18760
rect 41581 18726 41749 18760
rect 41953 18726 42121 18760
rect 42325 18726 42493 18760
rect 42697 18726 42865 18760
rect 43069 18726 43237 18760
rect 43441 18726 43609 18760
rect 43813 18726 43981 18760
rect 44185 18726 44353 18760
rect 44557 18726 44725 18760
rect 44929 18726 45097 18760
rect 45301 18726 45469 18760
rect 45673 18726 45841 18760
rect 46045 18726 46213 18760
rect 46417 18726 46585 18760
rect 46789 18726 46957 18760
rect 47161 18726 47329 18760
rect 47533 18726 47701 18760
rect 47905 18726 48073 18760
rect 48277 18726 48445 18760
rect 48649 18726 48817 18760
rect 49021 18726 49189 18760
rect 49393 18726 49561 18760
rect 40775 18500 40809 18676
rect 41033 18500 41067 18676
rect 41147 18500 41181 18676
rect 41405 18500 41439 18676
rect 41519 18500 41553 18676
rect 41777 18500 41811 18676
rect 41891 18500 41925 18676
rect 42149 18500 42183 18676
rect 42263 18500 42297 18676
rect 42521 18500 42555 18676
rect 42635 18500 42669 18676
rect 42893 18500 42927 18676
rect 43007 18500 43041 18676
rect 43265 18500 43299 18676
rect 43379 18500 43413 18676
rect 43637 18500 43671 18676
rect 43751 18500 43785 18676
rect 44009 18500 44043 18676
rect 44123 18500 44157 18676
rect 44381 18500 44415 18676
rect 44495 18500 44529 18676
rect 44753 18500 44787 18676
rect 44867 18500 44901 18676
rect 45125 18500 45159 18676
rect 45239 18500 45273 18676
rect 45497 18500 45531 18676
rect 45611 18500 45645 18676
rect 45869 18500 45903 18676
rect 45983 18500 46017 18676
rect 46241 18500 46275 18676
rect 46355 18500 46389 18676
rect 46613 18500 46647 18676
rect 46727 18500 46761 18676
rect 46985 18500 47019 18676
rect 47099 18500 47133 18676
rect 47357 18500 47391 18676
rect 47471 18500 47505 18676
rect 47729 18500 47763 18676
rect 47843 18500 47877 18676
rect 48101 18500 48135 18676
rect 48215 18500 48249 18676
rect 48473 18500 48507 18676
rect 48587 18500 48621 18676
rect 48845 18500 48879 18676
rect 48959 18500 48993 18676
rect 49217 18500 49251 18676
rect 49331 18500 49365 18676
rect 49589 18500 49623 18676
rect 40837 18416 41005 18450
rect 41209 18416 41377 18450
rect 41581 18416 41749 18450
rect 41953 18416 42121 18450
rect 42325 18416 42493 18450
rect 42697 18416 42865 18450
rect 43069 18416 43237 18450
rect 43441 18416 43609 18450
rect 43813 18416 43981 18450
rect 44185 18416 44353 18450
rect 44557 18416 44725 18450
rect 44929 18416 45097 18450
rect 45301 18416 45469 18450
rect 45673 18416 45841 18450
rect 46045 18416 46213 18450
rect 46417 18416 46585 18450
rect 46789 18416 46957 18450
rect 47161 18416 47329 18450
rect 47533 18416 47701 18450
rect 47905 18416 48073 18450
rect 48277 18416 48445 18450
rect 48649 18416 48817 18450
rect 49021 18416 49189 18450
rect 49393 18416 49561 18450
rect 40837 18308 41005 18342
rect 41209 18308 41377 18342
rect 41581 18308 41749 18342
rect 41953 18308 42121 18342
rect 42325 18308 42493 18342
rect 42697 18308 42865 18342
rect 43069 18308 43237 18342
rect 43441 18308 43609 18342
rect 43813 18308 43981 18342
rect 44185 18308 44353 18342
rect 44557 18308 44725 18342
rect 44929 18308 45097 18342
rect 45301 18308 45469 18342
rect 45673 18308 45841 18342
rect 46045 18308 46213 18342
rect 46417 18308 46585 18342
rect 46789 18308 46957 18342
rect 47161 18308 47329 18342
rect 47533 18308 47701 18342
rect 47905 18308 48073 18342
rect 48277 18308 48445 18342
rect 48649 18308 48817 18342
rect 49021 18308 49189 18342
rect 49393 18308 49561 18342
rect 40775 18082 40809 18258
rect 41033 18082 41067 18258
rect 41147 18082 41181 18258
rect 41405 18082 41439 18258
rect 41519 18082 41553 18258
rect 41777 18082 41811 18258
rect 41891 18082 41925 18258
rect 42149 18082 42183 18258
rect 42263 18082 42297 18258
rect 42521 18082 42555 18258
rect 42635 18082 42669 18258
rect 42893 18082 42927 18258
rect 43007 18082 43041 18258
rect 43265 18082 43299 18258
rect 43379 18082 43413 18258
rect 43637 18082 43671 18258
rect 43751 18082 43785 18258
rect 44009 18082 44043 18258
rect 44123 18082 44157 18258
rect 44381 18082 44415 18258
rect 44495 18082 44529 18258
rect 44753 18082 44787 18258
rect 44867 18082 44901 18258
rect 45125 18082 45159 18258
rect 45239 18082 45273 18258
rect 45497 18082 45531 18258
rect 45611 18082 45645 18258
rect 45869 18082 45903 18258
rect 45983 18082 46017 18258
rect 46241 18082 46275 18258
rect 46355 18082 46389 18258
rect 46613 18082 46647 18258
rect 46727 18082 46761 18258
rect 46985 18082 47019 18258
rect 47099 18082 47133 18258
rect 47357 18082 47391 18258
rect 47471 18082 47505 18258
rect 47729 18082 47763 18258
rect 47843 18082 47877 18258
rect 48101 18082 48135 18258
rect 48215 18082 48249 18258
rect 48473 18082 48507 18258
rect 48587 18082 48621 18258
rect 48845 18082 48879 18258
rect 48959 18082 48993 18258
rect 49217 18082 49251 18258
rect 49331 18082 49365 18258
rect 49589 18082 49623 18258
rect 40837 17998 41005 18032
rect 41209 17998 41377 18032
rect 41581 17998 41749 18032
rect 41953 17998 42121 18032
rect 42325 17998 42493 18032
rect 42697 17998 42865 18032
rect 43069 17998 43237 18032
rect 43441 17998 43609 18032
rect 43813 17998 43981 18032
rect 44185 17998 44353 18032
rect 44557 17998 44725 18032
rect 44929 17998 45097 18032
rect 45301 17998 45469 18032
rect 45673 17998 45841 18032
rect 46045 17998 46213 18032
rect 46417 17998 46585 18032
rect 46789 17998 46957 18032
rect 47161 17998 47329 18032
rect 47533 17998 47701 18032
rect 47905 17998 48073 18032
rect 48277 17998 48445 18032
rect 48649 17998 48817 18032
rect 49021 17998 49189 18032
rect 49393 17998 49561 18032
rect 40837 17340 41005 17374
rect 41209 17340 41377 17374
rect 41581 17340 41749 17374
rect 41953 17340 42121 17374
rect 42325 17340 42493 17374
rect 42697 17340 42865 17374
rect 43069 17340 43237 17374
rect 43441 17340 43609 17374
rect 40775 16505 40809 17281
rect 41033 16505 41067 17281
rect 41147 16505 41181 17281
rect 41405 16505 41439 17281
rect 41519 16505 41553 17281
rect 41777 16505 41811 17281
rect 41891 16505 41925 17281
rect 42149 16505 42183 17281
rect 42263 16505 42297 17281
rect 42521 16505 42555 17281
rect 42635 16505 42669 17281
rect 42893 16505 42927 17281
rect 43007 16505 43041 17281
rect 43265 16505 43299 17281
rect 43379 16505 43413 17281
rect 43637 16505 43671 17281
rect 40837 16412 41005 16446
rect 41209 16412 41377 16446
rect 41581 16412 41749 16446
rect 41953 16412 42121 16446
rect 42325 16412 42493 16446
rect 42697 16412 42865 16446
rect 43069 16412 43237 16446
rect 43441 16412 43609 16446
rect 40837 16304 41005 16338
rect 41209 16304 41377 16338
rect 41581 16304 41749 16338
rect 41953 16304 42121 16338
rect 42325 16304 42493 16338
rect 42697 16304 42865 16338
rect 43069 16304 43237 16338
rect 43441 16304 43609 16338
rect 40775 15469 40809 16245
rect 41033 15469 41067 16245
rect 41147 15469 41181 16245
rect 41405 15469 41439 16245
rect 41519 15469 41553 16245
rect 41777 15469 41811 16245
rect 41891 15469 41925 16245
rect 42149 15469 42183 16245
rect 42263 15469 42297 16245
rect 42521 15469 42555 16245
rect 42635 15469 42669 16245
rect 42893 15469 42927 16245
rect 43007 15469 43041 16245
rect 43265 15469 43299 16245
rect 43379 15469 43413 16245
rect 43637 15469 43671 16245
rect 40837 15376 41005 15410
rect 41209 15376 41377 15410
rect 41581 15376 41749 15410
rect 41953 15376 42121 15410
rect 42325 15376 42493 15410
rect 42697 15376 42865 15410
rect 43069 15376 43237 15410
rect 43441 15376 43609 15410
rect 40837 15268 41005 15302
rect 41209 15268 41377 15302
rect 41581 15268 41749 15302
rect 41953 15268 42121 15302
rect 42325 15268 42493 15302
rect 42697 15268 42865 15302
rect 43069 15268 43237 15302
rect 43441 15268 43609 15302
rect 40775 14433 40809 15209
rect 41033 14433 41067 15209
rect 41147 14433 41181 15209
rect 41405 14433 41439 15209
rect 41519 14433 41553 15209
rect 41777 14433 41811 15209
rect 41891 14433 41925 15209
rect 42149 14433 42183 15209
rect 42263 14433 42297 15209
rect 42521 14433 42555 15209
rect 42635 14433 42669 15209
rect 42893 14433 42927 15209
rect 43007 14433 43041 15209
rect 43265 14433 43299 15209
rect 43379 14433 43413 15209
rect 43637 14433 43671 15209
rect 40837 14340 41005 14374
rect 41209 14340 41377 14374
rect 41581 14340 41749 14374
rect 41953 14340 42121 14374
rect 42325 14340 42493 14374
rect 42697 14340 42865 14374
rect 43069 14340 43237 14374
rect 43441 14340 43609 14374
rect 40837 14232 41005 14266
rect 41209 14232 41377 14266
rect 41581 14232 41749 14266
rect 41953 14232 42121 14266
rect 42325 14232 42493 14266
rect 42697 14232 42865 14266
rect 43069 14232 43237 14266
rect 43441 14232 43609 14266
rect 40775 13397 40809 14173
rect 41033 13397 41067 14173
rect 41147 13397 41181 14173
rect 41405 13397 41439 14173
rect 41519 13397 41553 14173
rect 41777 13397 41811 14173
rect 41891 13397 41925 14173
rect 42149 13397 42183 14173
rect 42263 13397 42297 14173
rect 42521 13397 42555 14173
rect 42635 13397 42669 14173
rect 42893 13397 42927 14173
rect 43007 13397 43041 14173
rect 43265 13397 43299 14173
rect 43379 13397 43413 14173
rect 43637 13397 43671 14173
rect 40837 13304 41005 13338
rect 41209 13304 41377 13338
rect 41581 13304 41749 13338
rect 41953 13304 42121 13338
rect 42325 13304 42493 13338
rect 42697 13304 42865 13338
rect 43069 13304 43237 13338
rect 43441 13304 43609 13338
rect 45813 16365 45825 16413
rect 45825 16365 45859 16413
rect 45859 16365 45867 16413
rect 45971 16037 46009 16434
rect 45813 15965 45825 16013
rect 45825 15965 45859 16013
rect 45859 15965 45867 16013
rect 45813 15565 45825 15613
rect 45825 15565 45859 15613
rect 45859 15565 45867 15613
rect 45971 15506 46009 15903
rect 40746 13236 40816 13255
rect 41118 13236 41188 13255
rect 41490 13236 41560 13255
rect 41862 13236 41932 13255
rect 42234 13236 42304 13255
rect 42606 13236 42676 13255
rect 42978 13236 43048 13255
rect 43350 13236 43420 13255
rect 43612 13236 43682 13255
rect 40746 13202 40757 13236
rect 40757 13202 40816 13236
rect 41118 13202 41188 13236
rect 41490 13202 41560 13236
rect 41862 13202 41932 13236
rect 42234 13202 42304 13236
rect 42606 13202 42676 13236
rect 42978 13202 43048 13236
rect 43350 13202 43420 13236
rect 43612 13202 43682 13236
rect 40746 13185 40816 13202
rect 41118 13185 41188 13202
rect 41490 13185 41560 13202
rect 41862 13185 41932 13202
rect 42234 13185 42304 13202
rect 42606 13185 42676 13202
rect 42978 13185 43048 13202
rect 43350 13185 43420 13202
rect 43612 13185 43682 13202
rect 39349 12716 39517 12750
rect 39721 12716 39889 12750
rect 40093 12716 40261 12750
rect 40465 12716 40633 12750
rect 40837 12716 41005 12750
rect 41209 12716 41377 12750
rect 41581 12716 41749 12750
rect 41953 12716 42121 12750
rect 42325 12716 42493 12750
rect 42697 12716 42865 12750
rect 43069 12716 43237 12750
rect 43441 12716 43609 12750
rect 43813 12716 43981 12750
rect 44185 12716 44353 12750
rect 44557 12716 44725 12750
rect 44929 12716 45097 12750
rect 45301 12716 45469 12750
rect 45673 12716 45841 12750
rect 46045 12716 46213 12750
rect 46417 12716 46585 12750
rect 46789 12716 46957 12750
rect 47161 12716 47329 12750
rect 47533 12716 47701 12750
rect 47905 12716 48073 12750
rect 48277 12716 48445 12750
rect 48649 12716 48817 12750
rect 49021 12716 49189 12750
rect 49393 12716 49561 12750
rect 49765 12716 49933 12750
rect 50137 12716 50305 12750
rect 50509 12716 50677 12750
rect 50881 12716 51049 12750
rect 39287 12281 39321 12657
rect 39545 12281 39579 12657
rect 39659 12281 39693 12657
rect 39917 12281 39951 12657
rect 40031 12281 40065 12657
rect 40289 12281 40323 12657
rect 40403 12281 40437 12657
rect 40661 12281 40695 12657
rect 40775 12281 40809 12657
rect 41033 12281 41067 12657
rect 41147 12281 41181 12657
rect 41405 12281 41439 12657
rect 41519 12281 41553 12657
rect 41777 12281 41811 12657
rect 41891 12281 41925 12657
rect 42149 12281 42183 12657
rect 42263 12281 42297 12657
rect 42521 12281 42555 12657
rect 42635 12281 42669 12657
rect 42893 12281 42927 12657
rect 43007 12281 43041 12657
rect 43265 12281 43299 12657
rect 43379 12281 43413 12657
rect 43637 12281 43671 12657
rect 43751 12281 43785 12657
rect 44009 12281 44043 12657
rect 44123 12281 44157 12657
rect 44381 12281 44415 12657
rect 44495 12281 44529 12657
rect 44753 12281 44787 12657
rect 44867 12281 44901 12657
rect 45125 12281 45159 12657
rect 45239 12281 45273 12657
rect 45497 12281 45531 12657
rect 45611 12281 45645 12657
rect 45869 12281 45903 12657
rect 45983 12281 46017 12657
rect 46241 12281 46275 12657
rect 46355 12281 46389 12657
rect 46613 12281 46647 12657
rect 46727 12281 46761 12657
rect 46985 12281 47019 12657
rect 47099 12281 47133 12657
rect 47357 12281 47391 12657
rect 47471 12281 47505 12657
rect 47729 12281 47763 12657
rect 47843 12281 47877 12657
rect 48101 12281 48135 12657
rect 48215 12281 48249 12657
rect 48473 12281 48507 12657
rect 48587 12281 48621 12657
rect 48845 12281 48879 12657
rect 48959 12281 48993 12657
rect 49217 12281 49251 12657
rect 49331 12281 49365 12657
rect 49589 12281 49623 12657
rect 49703 12281 49737 12657
rect 49961 12281 49995 12657
rect 50075 12281 50109 12657
rect 50333 12281 50367 12657
rect 50447 12281 50481 12657
rect 50705 12281 50739 12657
rect 50819 12281 50853 12657
rect 51077 12281 51111 12657
rect 39349 12188 39517 12222
rect 39721 12188 39889 12222
rect 40093 12188 40261 12222
rect 40465 12188 40633 12222
rect 40837 12188 41005 12222
rect 41209 12188 41377 12222
rect 41581 12188 41749 12222
rect 41953 12188 42121 12222
rect 42325 12188 42493 12222
rect 42697 12188 42865 12222
rect 43069 12188 43237 12222
rect 43441 12188 43609 12222
rect 43813 12188 43981 12222
rect 44185 12188 44353 12222
rect 44557 12188 44725 12222
rect 44929 12188 45097 12222
rect 45301 12188 45469 12222
rect 45673 12188 45841 12222
rect 46045 12188 46213 12222
rect 46417 12188 46585 12222
rect 46789 12188 46957 12222
rect 47161 12188 47329 12222
rect 47533 12188 47701 12222
rect 47905 12188 48073 12222
rect 48277 12188 48445 12222
rect 48649 12188 48817 12222
rect 49021 12188 49189 12222
rect 49393 12188 49561 12222
rect 49765 12188 49933 12222
rect 50137 12188 50305 12222
rect 50509 12188 50677 12222
rect 50881 12188 51049 12222
rect 39349 12080 39517 12114
rect 39721 12080 39889 12114
rect 40093 12080 40261 12114
rect 40465 12080 40633 12114
rect 40837 12080 41005 12114
rect 41209 12080 41377 12114
rect 41581 12080 41749 12114
rect 41953 12080 42121 12114
rect 42325 12080 42493 12114
rect 42697 12080 42865 12114
rect 43069 12080 43237 12114
rect 43441 12080 43609 12114
rect 43813 12080 43981 12114
rect 44185 12080 44353 12114
rect 44557 12080 44725 12114
rect 44929 12080 45097 12114
rect 45301 12080 45469 12114
rect 45673 12080 45841 12114
rect 46045 12080 46213 12114
rect 46417 12080 46585 12114
rect 46789 12080 46957 12114
rect 47161 12080 47329 12114
rect 47533 12080 47701 12114
rect 47905 12080 48073 12114
rect 48277 12080 48445 12114
rect 48649 12080 48817 12114
rect 49021 12080 49189 12114
rect 49393 12080 49561 12114
rect 49765 12080 49933 12114
rect 50137 12080 50305 12114
rect 50509 12080 50677 12114
rect 50881 12080 51049 12114
rect 39287 11645 39321 12021
rect 39545 11645 39579 12021
rect 39659 11645 39693 12021
rect 39917 11645 39951 12021
rect 40031 11645 40065 12021
rect 40289 11645 40323 12021
rect 40403 11645 40437 12021
rect 40661 11645 40695 12021
rect 40775 11645 40809 12021
rect 41033 11645 41067 12021
rect 41147 11645 41181 12021
rect 41405 11645 41439 12021
rect 41519 11645 41553 12021
rect 41777 11645 41811 12021
rect 41891 11645 41925 12021
rect 42149 11645 42183 12021
rect 42263 11645 42297 12021
rect 42521 11645 42555 12021
rect 42635 11645 42669 12021
rect 42893 11645 42927 12021
rect 43007 11645 43041 12021
rect 43265 11645 43299 12021
rect 43379 11645 43413 12021
rect 43637 11645 43671 12021
rect 43751 11645 43785 12021
rect 44009 11645 44043 12021
rect 44123 11645 44157 12021
rect 44381 11645 44415 12021
rect 44495 11645 44529 12021
rect 44753 11645 44787 12021
rect 44867 11645 44901 12021
rect 45125 11645 45159 12021
rect 45239 11645 45273 12021
rect 45497 11645 45531 12021
rect 45611 11645 45645 12021
rect 45869 11645 45903 12021
rect 45983 11645 46017 12021
rect 46241 11645 46275 12021
rect 46355 11645 46389 12021
rect 46613 11645 46647 12021
rect 46727 11645 46761 12021
rect 46985 11645 47019 12021
rect 47099 11645 47133 12021
rect 47357 11645 47391 12021
rect 47471 11645 47505 12021
rect 47729 11645 47763 12021
rect 47843 11645 47877 12021
rect 48101 11645 48135 12021
rect 48215 11645 48249 12021
rect 48473 11645 48507 12021
rect 48587 11645 48621 12021
rect 48845 11645 48879 12021
rect 48959 11645 48993 12021
rect 49217 11645 49251 12021
rect 49331 11645 49365 12021
rect 49589 11645 49623 12021
rect 49703 11645 49737 12021
rect 49961 11645 49995 12021
rect 50075 11645 50109 12021
rect 50333 11645 50367 12021
rect 50447 11645 50481 12021
rect 50705 11645 50739 12021
rect 50819 11645 50853 12021
rect 51077 11645 51111 12021
rect 39349 11552 39517 11586
rect 39721 11552 39889 11586
rect 40093 11552 40261 11586
rect 40465 11552 40633 11586
rect 40837 11552 41005 11586
rect 41209 11552 41377 11586
rect 41581 11552 41749 11586
rect 41953 11552 42121 11586
rect 42325 11552 42493 11586
rect 42697 11552 42865 11586
rect 43069 11552 43237 11586
rect 43441 11552 43609 11586
rect 43813 11552 43981 11586
rect 44185 11552 44353 11586
rect 44557 11552 44725 11586
rect 44929 11552 45097 11586
rect 45301 11552 45469 11586
rect 45673 11552 45841 11586
rect 46045 11552 46213 11586
rect 46417 11552 46585 11586
rect 46789 11552 46957 11586
rect 47161 11552 47329 11586
rect 47533 11552 47701 11586
rect 47905 11552 48073 11586
rect 48277 11552 48445 11586
rect 48649 11552 48817 11586
rect 49021 11552 49189 11586
rect 49393 11552 49561 11586
rect 49765 11552 49933 11586
rect 50137 11552 50305 11586
rect 50509 11552 50677 11586
rect 50881 11552 51049 11586
rect 39349 11444 39517 11478
rect 39721 11444 39889 11478
rect 40093 11444 40261 11478
rect 40465 11444 40633 11478
rect 40837 11444 41005 11478
rect 41209 11444 41377 11478
rect 41581 11444 41749 11478
rect 41953 11444 42121 11478
rect 42325 11444 42493 11478
rect 42697 11444 42865 11478
rect 43069 11444 43237 11478
rect 43441 11444 43609 11478
rect 43813 11444 43981 11478
rect 44185 11444 44353 11478
rect 44557 11444 44725 11478
rect 44929 11444 45097 11478
rect 45301 11444 45469 11478
rect 45673 11444 45841 11478
rect 46045 11444 46213 11478
rect 46417 11444 46585 11478
rect 46789 11444 46957 11478
rect 47161 11444 47329 11478
rect 47533 11444 47701 11478
rect 47905 11444 48073 11478
rect 48277 11444 48445 11478
rect 48649 11444 48817 11478
rect 49021 11444 49189 11478
rect 49393 11444 49561 11478
rect 49765 11444 49933 11478
rect 50137 11444 50305 11478
rect 50509 11444 50677 11478
rect 50881 11444 51049 11478
rect 39287 11009 39321 11385
rect 39545 11009 39579 11385
rect 39659 11009 39693 11385
rect 39917 11009 39951 11385
rect 40031 11009 40065 11385
rect 40289 11009 40323 11385
rect 40403 11009 40437 11385
rect 40661 11009 40695 11385
rect 40775 11009 40809 11385
rect 41033 11009 41067 11385
rect 41147 11009 41181 11385
rect 41405 11009 41439 11385
rect 41519 11009 41553 11385
rect 41777 11009 41811 11385
rect 41891 11009 41925 11385
rect 42149 11009 42183 11385
rect 42263 11009 42297 11385
rect 42521 11009 42555 11385
rect 42635 11009 42669 11385
rect 42893 11009 42927 11385
rect 43007 11009 43041 11385
rect 43265 11009 43299 11385
rect 43379 11009 43413 11385
rect 43637 11009 43671 11385
rect 43751 11009 43785 11385
rect 44009 11009 44043 11385
rect 44123 11009 44157 11385
rect 44381 11009 44415 11385
rect 44495 11009 44529 11385
rect 44753 11009 44787 11385
rect 44867 11009 44901 11385
rect 45125 11009 45159 11385
rect 45239 11009 45273 11385
rect 45497 11009 45531 11385
rect 45611 11009 45645 11385
rect 45869 11009 45903 11385
rect 45983 11009 46017 11385
rect 46241 11009 46275 11385
rect 46355 11009 46389 11385
rect 46613 11009 46647 11385
rect 46727 11009 46761 11385
rect 46985 11009 47019 11385
rect 47099 11009 47133 11385
rect 47357 11009 47391 11385
rect 47471 11009 47505 11385
rect 47729 11009 47763 11385
rect 47843 11009 47877 11385
rect 48101 11009 48135 11385
rect 48215 11009 48249 11385
rect 48473 11009 48507 11385
rect 48587 11009 48621 11385
rect 48845 11009 48879 11385
rect 48959 11009 48993 11385
rect 49217 11009 49251 11385
rect 49331 11009 49365 11385
rect 49589 11009 49623 11385
rect 49703 11009 49737 11385
rect 49961 11009 49995 11385
rect 50075 11009 50109 11385
rect 50333 11009 50367 11385
rect 50447 11009 50481 11385
rect 50705 11009 50739 11385
rect 50819 11009 50853 11385
rect 51077 11009 51111 11385
rect 39349 10916 39517 10950
rect 39721 10916 39889 10950
rect 40093 10916 40261 10950
rect 40465 10916 40633 10950
rect 40837 10916 41005 10950
rect 41209 10916 41377 10950
rect 41581 10916 41749 10950
rect 41953 10916 42121 10950
rect 42325 10916 42493 10950
rect 42697 10916 42865 10950
rect 43069 10916 43237 10950
rect 43441 10916 43609 10950
rect 43813 10916 43981 10950
rect 44185 10916 44353 10950
rect 44557 10916 44725 10950
rect 44929 10916 45097 10950
rect 45301 10916 45469 10950
rect 45673 10916 45841 10950
rect 46045 10916 46213 10950
rect 46417 10916 46585 10950
rect 46789 10916 46957 10950
rect 47161 10916 47329 10950
rect 47533 10916 47701 10950
rect 47905 10916 48073 10950
rect 48277 10916 48445 10950
rect 48649 10916 48817 10950
rect 49021 10916 49189 10950
rect 49393 10916 49561 10950
rect 49765 10916 49933 10950
rect 50137 10916 50305 10950
rect 50509 10916 50677 10950
rect 50881 10916 51049 10950
rect 39584 10848 39654 10867
rect 40328 10848 40398 10867
rect 41072 10848 41142 10867
rect 41816 10848 41886 10867
rect 42560 10848 42630 10867
rect 43304 10848 43374 10867
rect 44048 10848 44118 10867
rect 44792 10848 44862 10867
rect 45164 10848 45234 10867
rect 45908 10848 45978 10867
rect 46652 10848 46722 10867
rect 47396 10848 47466 10867
rect 48140 10848 48210 10867
rect 48884 10848 48954 10867
rect 49628 10848 49698 10867
rect 50372 10848 50442 10867
rect 51062 10848 51132 10867
rect 39584 10814 39654 10848
rect 40328 10814 40398 10848
rect 41072 10814 41142 10848
rect 41816 10814 41886 10848
rect 42560 10814 42630 10848
rect 43304 10814 43374 10848
rect 44048 10814 44118 10848
rect 44792 10814 44862 10848
rect 45164 10814 45234 10848
rect 45908 10814 45978 10848
rect 46652 10814 46722 10848
rect 47396 10814 47466 10848
rect 48140 10814 48210 10848
rect 48884 10814 48954 10848
rect 49628 10814 49698 10848
rect 50372 10814 50442 10848
rect 51062 10814 51129 10848
rect 51129 10814 51132 10848
rect 39584 10797 39654 10814
rect 40328 10797 40398 10814
rect 41072 10797 41142 10814
rect 41816 10797 41886 10814
rect 42560 10797 42630 10814
rect 43304 10797 43374 10814
rect 44048 10797 44118 10814
rect 44792 10797 44862 10814
rect 45164 10797 45234 10814
rect 45908 10797 45978 10814
rect 46652 10797 46722 10814
rect 47396 10797 47466 10814
rect 48140 10797 48210 10814
rect 48884 10797 48954 10814
rect 49628 10797 49698 10814
rect 50372 10797 50442 10814
rect 51062 10797 51132 10814
rect 39584 9051 39654 9068
rect 40328 9051 40398 9068
rect 41072 9051 41142 9068
rect 41816 9051 41886 9068
rect 42560 9051 42630 9068
rect 43304 9051 43374 9068
rect 44048 9051 44118 9068
rect 44792 9051 44862 9068
rect 45164 9051 45234 9068
rect 45908 9051 45978 9068
rect 46652 9051 46722 9068
rect 47396 9051 47466 9068
rect 48140 9051 48210 9068
rect 48884 9051 48954 9068
rect 49628 9051 49698 9068
rect 50372 9051 50442 9068
rect 51062 9051 51132 9068
rect 39584 9017 39654 9051
rect 40328 9017 40398 9051
rect 41072 9017 41142 9051
rect 41816 9017 41886 9051
rect 42560 9017 42630 9051
rect 43304 9017 43374 9051
rect 44048 9017 44118 9051
rect 44792 9017 44862 9051
rect 45164 9017 45234 9051
rect 45908 9017 45978 9051
rect 46652 9017 46722 9051
rect 47396 9017 47466 9051
rect 48140 9017 48210 9051
rect 48884 9017 48954 9051
rect 49628 9017 49698 9051
rect 50372 9017 50442 9051
rect 51062 9017 51129 9051
rect 51129 9017 51132 9051
rect 39584 8998 39654 9017
rect 40328 8998 40398 9017
rect 41072 8998 41142 9017
rect 41816 8998 41886 9017
rect 42560 8998 42630 9017
rect 43304 8998 43374 9017
rect 44048 8998 44118 9017
rect 44792 8998 44862 9017
rect 45164 8998 45234 9017
rect 45908 8998 45978 9017
rect 46652 8998 46722 9017
rect 47396 8998 47466 9017
rect 48140 8998 48210 9017
rect 48884 8998 48954 9017
rect 49628 8998 49698 9017
rect 50372 8998 50442 9017
rect 51062 8998 51132 9017
rect 39349 8915 39517 8949
rect 39721 8915 39889 8949
rect 40093 8915 40261 8949
rect 40465 8915 40633 8949
rect 40837 8915 41005 8949
rect 41209 8915 41377 8949
rect 41581 8915 41749 8949
rect 41953 8915 42121 8949
rect 42325 8915 42493 8949
rect 42697 8915 42865 8949
rect 43069 8915 43237 8949
rect 43441 8915 43609 8949
rect 43813 8915 43981 8949
rect 44185 8915 44353 8949
rect 44557 8915 44725 8949
rect 44929 8915 45097 8949
rect 45301 8915 45469 8949
rect 45673 8915 45841 8949
rect 46045 8915 46213 8949
rect 46417 8915 46585 8949
rect 46789 8915 46957 8949
rect 47161 8915 47329 8949
rect 47533 8915 47701 8949
rect 47905 8915 48073 8949
rect 48277 8915 48445 8949
rect 48649 8915 48817 8949
rect 49021 8915 49189 8949
rect 49393 8915 49561 8949
rect 49765 8915 49933 8949
rect 50137 8915 50305 8949
rect 50509 8915 50677 8949
rect 50881 8915 51049 8949
rect 39287 8480 39321 8856
rect 39545 8480 39579 8856
rect 39659 8480 39693 8856
rect 39917 8480 39951 8856
rect 40031 8480 40065 8856
rect 40289 8480 40323 8856
rect 40403 8480 40437 8856
rect 40661 8480 40695 8856
rect 40775 8480 40809 8856
rect 41033 8480 41067 8856
rect 41147 8480 41181 8856
rect 41405 8480 41439 8856
rect 41519 8480 41553 8856
rect 41777 8480 41811 8856
rect 41891 8480 41925 8856
rect 42149 8480 42183 8856
rect 42263 8480 42297 8856
rect 42521 8480 42555 8856
rect 42635 8480 42669 8856
rect 42893 8480 42927 8856
rect 43007 8480 43041 8856
rect 43265 8480 43299 8856
rect 43379 8480 43413 8856
rect 43637 8480 43671 8856
rect 43751 8480 43785 8856
rect 44009 8480 44043 8856
rect 44123 8480 44157 8856
rect 44381 8480 44415 8856
rect 44495 8480 44529 8856
rect 44753 8480 44787 8856
rect 44867 8480 44901 8856
rect 45125 8480 45159 8856
rect 45239 8480 45273 8856
rect 45497 8480 45531 8856
rect 45611 8480 45645 8856
rect 45869 8480 45903 8856
rect 45983 8480 46017 8856
rect 46241 8480 46275 8856
rect 46355 8480 46389 8856
rect 46613 8480 46647 8856
rect 46727 8480 46761 8856
rect 46985 8480 47019 8856
rect 47099 8480 47133 8856
rect 47357 8480 47391 8856
rect 47471 8480 47505 8856
rect 47729 8480 47763 8856
rect 47843 8480 47877 8856
rect 48101 8480 48135 8856
rect 48215 8480 48249 8856
rect 48473 8480 48507 8856
rect 48587 8480 48621 8856
rect 48845 8480 48879 8856
rect 48959 8480 48993 8856
rect 49217 8480 49251 8856
rect 49331 8480 49365 8856
rect 49589 8480 49623 8856
rect 49703 8480 49737 8856
rect 49961 8480 49995 8856
rect 50075 8480 50109 8856
rect 50333 8480 50367 8856
rect 50447 8480 50481 8856
rect 50705 8480 50739 8856
rect 50819 8480 50853 8856
rect 51077 8480 51111 8856
rect 39349 8387 39517 8421
rect 39721 8387 39889 8421
rect 40093 8387 40261 8421
rect 40465 8387 40633 8421
rect 40837 8387 41005 8421
rect 41209 8387 41377 8421
rect 41581 8387 41749 8421
rect 41953 8387 42121 8421
rect 42325 8387 42493 8421
rect 42697 8387 42865 8421
rect 43069 8387 43237 8421
rect 43441 8387 43609 8421
rect 43813 8387 43981 8421
rect 44185 8387 44353 8421
rect 44557 8387 44725 8421
rect 44929 8387 45097 8421
rect 45301 8387 45469 8421
rect 45673 8387 45841 8421
rect 46045 8387 46213 8421
rect 46417 8387 46585 8421
rect 46789 8387 46957 8421
rect 47161 8387 47329 8421
rect 47533 8387 47701 8421
rect 47905 8387 48073 8421
rect 48277 8387 48445 8421
rect 48649 8387 48817 8421
rect 49021 8387 49189 8421
rect 49393 8387 49561 8421
rect 49765 8387 49933 8421
rect 50137 8387 50305 8421
rect 50509 8387 50677 8421
rect 50881 8387 51049 8421
rect 39349 8279 39517 8313
rect 39721 8279 39889 8313
rect 40093 8279 40261 8313
rect 40465 8279 40633 8313
rect 40837 8279 41005 8313
rect 41209 8279 41377 8313
rect 41581 8279 41749 8313
rect 41953 8279 42121 8313
rect 42325 8279 42493 8313
rect 42697 8279 42865 8313
rect 43069 8279 43237 8313
rect 43441 8279 43609 8313
rect 43813 8279 43981 8313
rect 44185 8279 44353 8313
rect 44557 8279 44725 8313
rect 44929 8279 45097 8313
rect 45301 8279 45469 8313
rect 45673 8279 45841 8313
rect 46045 8279 46213 8313
rect 46417 8279 46585 8313
rect 46789 8279 46957 8313
rect 47161 8279 47329 8313
rect 47533 8279 47701 8313
rect 47905 8279 48073 8313
rect 48277 8279 48445 8313
rect 48649 8279 48817 8313
rect 49021 8279 49189 8313
rect 49393 8279 49561 8313
rect 49765 8279 49933 8313
rect 50137 8279 50305 8313
rect 50509 8279 50677 8313
rect 50881 8279 51049 8313
rect 39287 7844 39321 8220
rect 39545 7844 39579 8220
rect 39659 7844 39693 8220
rect 39917 7844 39951 8220
rect 40031 7844 40065 8220
rect 40289 7844 40323 8220
rect 40403 7844 40437 8220
rect 40661 7844 40695 8220
rect 40775 7844 40809 8220
rect 41033 7844 41067 8220
rect 41147 7844 41181 8220
rect 41405 7844 41439 8220
rect 41519 7844 41553 8220
rect 41777 7844 41811 8220
rect 41891 7844 41925 8220
rect 42149 7844 42183 8220
rect 42263 7844 42297 8220
rect 42521 7844 42555 8220
rect 42635 7844 42669 8220
rect 42893 7844 42927 8220
rect 43007 7844 43041 8220
rect 43265 7844 43299 8220
rect 43379 7844 43413 8220
rect 43637 7844 43671 8220
rect 43751 7844 43785 8220
rect 44009 7844 44043 8220
rect 44123 7844 44157 8220
rect 44381 7844 44415 8220
rect 44495 7844 44529 8220
rect 44753 7844 44787 8220
rect 44867 7844 44901 8220
rect 45125 7844 45159 8220
rect 45239 7844 45273 8220
rect 45497 7844 45531 8220
rect 45611 7844 45645 8220
rect 45869 7844 45903 8220
rect 45983 7844 46017 8220
rect 46241 7844 46275 8220
rect 46355 7844 46389 8220
rect 46613 7844 46647 8220
rect 46727 7844 46761 8220
rect 46985 7844 47019 8220
rect 47099 7844 47133 8220
rect 47357 7844 47391 8220
rect 47471 7844 47505 8220
rect 47729 7844 47763 8220
rect 47843 7844 47877 8220
rect 48101 7844 48135 8220
rect 48215 7844 48249 8220
rect 48473 7844 48507 8220
rect 48587 7844 48621 8220
rect 48845 7844 48879 8220
rect 48959 7844 48993 8220
rect 49217 7844 49251 8220
rect 49331 7844 49365 8220
rect 49589 7844 49623 8220
rect 49703 7844 49737 8220
rect 49961 7844 49995 8220
rect 50075 7844 50109 8220
rect 50333 7844 50367 8220
rect 50447 7844 50481 8220
rect 50705 7844 50739 8220
rect 50819 7844 50853 8220
rect 51077 7844 51111 8220
rect 39349 7751 39517 7785
rect 39721 7751 39889 7785
rect 40093 7751 40261 7785
rect 40465 7751 40633 7785
rect 40837 7751 41005 7785
rect 41209 7751 41377 7785
rect 41581 7751 41749 7785
rect 41953 7751 42121 7785
rect 42325 7751 42493 7785
rect 42697 7751 42865 7785
rect 43069 7751 43237 7785
rect 43441 7751 43609 7785
rect 43813 7751 43981 7785
rect 44185 7751 44353 7785
rect 44557 7751 44725 7785
rect 44929 7751 45097 7785
rect 45301 7751 45469 7785
rect 45673 7751 45841 7785
rect 46045 7751 46213 7785
rect 46417 7751 46585 7785
rect 46789 7751 46957 7785
rect 47161 7751 47329 7785
rect 47533 7751 47701 7785
rect 47905 7751 48073 7785
rect 48277 7751 48445 7785
rect 48649 7751 48817 7785
rect 49021 7751 49189 7785
rect 49393 7751 49561 7785
rect 49765 7751 49933 7785
rect 50137 7751 50305 7785
rect 50509 7751 50677 7785
rect 50881 7751 51049 7785
rect 39349 7643 39517 7677
rect 39721 7643 39889 7677
rect 40093 7643 40261 7677
rect 40465 7643 40633 7677
rect 40837 7643 41005 7677
rect 41209 7643 41377 7677
rect 41581 7643 41749 7677
rect 41953 7643 42121 7677
rect 42325 7643 42493 7677
rect 42697 7643 42865 7677
rect 43069 7643 43237 7677
rect 43441 7643 43609 7677
rect 43813 7643 43981 7677
rect 44185 7643 44353 7677
rect 44557 7643 44725 7677
rect 44929 7643 45097 7677
rect 45301 7643 45469 7677
rect 45673 7643 45841 7677
rect 46045 7643 46213 7677
rect 46417 7643 46585 7677
rect 46789 7643 46957 7677
rect 47161 7643 47329 7677
rect 47533 7643 47701 7677
rect 47905 7643 48073 7677
rect 48277 7643 48445 7677
rect 48649 7643 48817 7677
rect 49021 7643 49189 7677
rect 49393 7643 49561 7677
rect 49765 7643 49933 7677
rect 50137 7643 50305 7677
rect 50509 7643 50677 7677
rect 50881 7643 51049 7677
rect 39287 7208 39321 7584
rect 39545 7208 39579 7584
rect 39659 7208 39693 7584
rect 39917 7208 39951 7584
rect 40031 7208 40065 7584
rect 40289 7208 40323 7584
rect 40403 7208 40437 7584
rect 40661 7208 40695 7584
rect 40775 7208 40809 7584
rect 41033 7208 41067 7584
rect 41147 7208 41181 7584
rect 41405 7208 41439 7584
rect 41519 7208 41553 7584
rect 41777 7208 41811 7584
rect 41891 7208 41925 7584
rect 42149 7208 42183 7584
rect 42263 7208 42297 7584
rect 42521 7208 42555 7584
rect 42635 7208 42669 7584
rect 42893 7208 42927 7584
rect 43007 7208 43041 7584
rect 43265 7208 43299 7584
rect 43379 7208 43413 7584
rect 43637 7208 43671 7584
rect 43751 7208 43785 7584
rect 44009 7208 44043 7584
rect 44123 7208 44157 7584
rect 44381 7208 44415 7584
rect 44495 7208 44529 7584
rect 44753 7208 44787 7584
rect 44867 7208 44901 7584
rect 45125 7208 45159 7584
rect 45239 7208 45273 7584
rect 45497 7208 45531 7584
rect 45611 7208 45645 7584
rect 45869 7208 45903 7584
rect 45983 7208 46017 7584
rect 46241 7208 46275 7584
rect 46355 7208 46389 7584
rect 46613 7208 46647 7584
rect 46727 7208 46761 7584
rect 46985 7208 47019 7584
rect 47099 7208 47133 7584
rect 47357 7208 47391 7584
rect 47471 7208 47505 7584
rect 47729 7208 47763 7584
rect 47843 7208 47877 7584
rect 48101 7208 48135 7584
rect 48215 7208 48249 7584
rect 48473 7208 48507 7584
rect 48587 7208 48621 7584
rect 48845 7208 48879 7584
rect 48959 7208 48993 7584
rect 49217 7208 49251 7584
rect 49331 7208 49365 7584
rect 49589 7208 49623 7584
rect 49703 7208 49737 7584
rect 49961 7208 49995 7584
rect 50075 7208 50109 7584
rect 50333 7208 50367 7584
rect 50447 7208 50481 7584
rect 50705 7208 50739 7584
rect 50819 7208 50853 7584
rect 51077 7208 51111 7584
rect 39349 7115 39517 7149
rect 39721 7115 39889 7149
rect 40093 7115 40261 7149
rect 40465 7115 40633 7149
rect 40837 7115 41005 7149
rect 41209 7115 41377 7149
rect 41581 7115 41749 7149
rect 41953 7115 42121 7149
rect 42325 7115 42493 7149
rect 42697 7115 42865 7149
rect 43069 7115 43237 7149
rect 43441 7115 43609 7149
rect 43813 7115 43981 7149
rect 44185 7115 44353 7149
rect 44557 7115 44725 7149
rect 44929 7115 45097 7149
rect 45301 7115 45469 7149
rect 45673 7115 45841 7149
rect 46045 7115 46213 7149
rect 46417 7115 46585 7149
rect 46789 7115 46957 7149
rect 47161 7115 47329 7149
rect 47533 7115 47701 7149
rect 47905 7115 48073 7149
rect 48277 7115 48445 7149
rect 48649 7115 48817 7149
rect 49021 7115 49189 7149
rect 49393 7115 49561 7149
rect 49765 7115 49933 7149
rect 50137 7115 50305 7149
rect 50509 7115 50677 7149
rect 50881 7115 51049 7149
rect 39521 6325 39559 6722
rect 39839 6325 39877 6722
rect 40746 6663 40816 6680
rect 41118 6663 41188 6680
rect 41490 6663 41560 6680
rect 41862 6663 41932 6680
rect 42234 6663 42304 6680
rect 42606 6663 42676 6680
rect 42978 6663 43048 6680
rect 43350 6663 43420 6680
rect 43612 6663 43682 6680
rect 40746 6629 40757 6663
rect 40757 6629 40816 6663
rect 41118 6629 41188 6663
rect 41490 6629 41560 6663
rect 41862 6629 41932 6663
rect 42234 6629 42304 6663
rect 42606 6629 42676 6663
rect 42978 6629 43048 6663
rect 43350 6629 43420 6663
rect 43612 6629 43682 6663
rect 40746 6610 40816 6629
rect 41118 6610 41188 6629
rect 41490 6610 41560 6629
rect 41862 6610 41932 6629
rect 42234 6610 42304 6629
rect 42606 6610 42676 6629
rect 42978 6610 43048 6629
rect 43350 6610 43420 6629
rect 43612 6610 43682 6629
rect 39970 6153 39989 6219
rect 39989 6153 40023 6219
rect 40023 6153 40042 6219
rect 39970 5755 39989 5819
rect 39989 5755 40023 5819
rect 40023 5755 40042 5819
rect 39970 5355 39989 5419
rect 39989 5355 40023 5419
rect 40023 5355 40042 5419
rect 39521 4894 39559 5291
rect 39839 4894 39877 5291
rect 39970 4955 39989 5019
rect 39989 4955 40023 5019
rect 40023 4955 40042 5019
rect 40837 6527 41005 6561
rect 41209 6527 41377 6561
rect 41581 6527 41749 6561
rect 41953 6527 42121 6561
rect 42325 6527 42493 6561
rect 42697 6527 42865 6561
rect 43069 6527 43237 6561
rect 43441 6527 43609 6561
rect 40775 5692 40809 6468
rect 41033 5692 41067 6468
rect 41147 5692 41181 6468
rect 41405 5692 41439 6468
rect 41519 5692 41553 6468
rect 41777 5692 41811 6468
rect 41891 5692 41925 6468
rect 42149 5692 42183 6468
rect 42263 5692 42297 6468
rect 42521 5692 42555 6468
rect 42635 5692 42669 6468
rect 42893 5692 42927 6468
rect 43007 5692 43041 6468
rect 43265 5692 43299 6468
rect 43379 5692 43413 6468
rect 43637 5692 43671 6468
rect 40837 5599 41005 5633
rect 41209 5599 41377 5633
rect 41581 5599 41749 5633
rect 41953 5599 42121 5633
rect 42325 5599 42493 5633
rect 42697 5599 42865 5633
rect 43069 5599 43237 5633
rect 43441 5599 43609 5633
rect 40837 5491 41005 5525
rect 41209 5491 41377 5525
rect 41581 5491 41749 5525
rect 41953 5491 42121 5525
rect 42325 5491 42493 5525
rect 42697 5491 42865 5525
rect 43069 5491 43237 5525
rect 43441 5491 43609 5525
rect 40775 4656 40809 5432
rect 41033 4656 41067 5432
rect 41147 4656 41181 5432
rect 41405 4656 41439 5432
rect 41519 4656 41553 5432
rect 41777 4656 41811 5432
rect 41891 4656 41925 5432
rect 42149 4656 42183 5432
rect 42263 4656 42297 5432
rect 42521 4656 42555 5432
rect 42635 4656 42669 5432
rect 42893 4656 42927 5432
rect 43007 4656 43041 5432
rect 43265 4656 43299 5432
rect 43379 4656 43413 5432
rect 43637 4656 43671 5432
rect 40837 4563 41005 4597
rect 41209 4563 41377 4597
rect 41581 4563 41749 4597
rect 41953 4563 42121 4597
rect 42325 4563 42493 4597
rect 42697 4563 42865 4597
rect 43069 4563 43237 4597
rect 43441 4563 43609 4597
rect 40837 4455 41005 4489
rect 41209 4455 41377 4489
rect 41581 4455 41749 4489
rect 41953 4455 42121 4489
rect 42325 4455 42493 4489
rect 42697 4455 42865 4489
rect 43069 4455 43237 4489
rect 43441 4455 43609 4489
rect 40775 3620 40809 4396
rect 41033 3620 41067 4396
rect 41147 3620 41181 4396
rect 41405 3620 41439 4396
rect 41519 3620 41553 4396
rect 41777 3620 41811 4396
rect 41891 3620 41925 4396
rect 42149 3620 42183 4396
rect 42263 3620 42297 4396
rect 42521 3620 42555 4396
rect 42635 3620 42669 4396
rect 42893 3620 42927 4396
rect 43007 3620 43041 4396
rect 43265 3620 43299 4396
rect 43379 3620 43413 4396
rect 43637 3620 43671 4396
rect 40837 3527 41005 3561
rect 41209 3527 41377 3561
rect 41581 3527 41749 3561
rect 41953 3527 42121 3561
rect 42325 3527 42493 3561
rect 42697 3527 42865 3561
rect 43069 3527 43237 3561
rect 43441 3527 43609 3561
rect 40837 3419 41005 3453
rect 41209 3419 41377 3453
rect 41581 3419 41749 3453
rect 41953 3419 42121 3453
rect 42325 3419 42493 3453
rect 42697 3419 42865 3453
rect 43069 3419 43237 3453
rect 43441 3419 43609 3453
rect 40775 2584 40809 3360
rect 41033 2584 41067 3360
rect 41147 2584 41181 3360
rect 41405 2584 41439 3360
rect 41519 2584 41553 3360
rect 41777 2584 41811 3360
rect 41891 2584 41925 3360
rect 42149 2584 42183 3360
rect 42263 2584 42297 3360
rect 42521 2584 42555 3360
rect 42635 2584 42669 3360
rect 42893 2584 42927 3360
rect 43007 2584 43041 3360
rect 43265 2584 43299 3360
rect 43379 2584 43413 3360
rect 43637 2584 43671 3360
rect 40837 2491 41005 2525
rect 41209 2491 41377 2525
rect 41581 2491 41749 2525
rect 41953 2491 42121 2525
rect 42325 2491 42493 2525
rect 42697 2491 42865 2525
rect 43069 2491 43237 2525
rect 43441 2491 43609 2525
rect 44677 5685 44715 6082
rect 44512 5613 44531 5679
rect 44531 5613 44565 5679
rect 44565 5613 44584 5679
rect 44995 5685 45033 6082
rect 44512 5215 44531 5279
rect 44531 5215 44565 5279
rect 44565 5215 44584 5279
rect 44512 4815 44531 4879
rect 44531 4815 44565 4879
rect 44565 4815 44584 4879
rect 44512 4415 44531 4479
rect 44531 4415 44565 4479
rect 44565 4415 44584 4479
rect 44677 4254 44715 4651
rect 44995 4254 45033 4651
rect 45812 4186 45825 4240
rect 45825 4186 45859 4240
rect 45859 4186 45870 4240
rect 45971 3962 46009 4359
rect 45812 3786 45825 3840
rect 45825 3786 45859 3840
rect 45859 3786 45870 3840
rect 45812 3386 45825 3440
rect 45825 3386 45859 3440
rect 45859 3386 45870 3440
rect 45971 3431 46009 3828
rect 40837 1833 41005 1867
rect 41209 1833 41377 1867
rect 41581 1833 41749 1867
rect 41953 1833 42121 1867
rect 42325 1833 42493 1867
rect 42697 1833 42865 1867
rect 43069 1833 43237 1867
rect 43441 1833 43609 1867
rect 43813 1833 43981 1867
rect 44185 1833 44353 1867
rect 44557 1833 44725 1867
rect 44929 1833 45097 1867
rect 45301 1833 45469 1867
rect 45673 1833 45841 1867
rect 46045 1833 46213 1867
rect 46417 1833 46585 1867
rect 46789 1833 46957 1867
rect 47161 1833 47329 1867
rect 47533 1833 47701 1867
rect 47905 1833 48073 1867
rect 48277 1833 48445 1867
rect 48649 1833 48817 1867
rect 49021 1833 49189 1867
rect 49393 1833 49561 1867
rect 40775 1607 40809 1783
rect 41033 1607 41067 1783
rect 41147 1607 41181 1783
rect 41405 1607 41439 1783
rect 41519 1607 41553 1783
rect 41777 1607 41811 1783
rect 41891 1607 41925 1783
rect 42149 1607 42183 1783
rect 42263 1607 42297 1783
rect 42521 1607 42555 1783
rect 42635 1607 42669 1783
rect 42893 1607 42927 1783
rect 43007 1607 43041 1783
rect 43265 1607 43299 1783
rect 43379 1607 43413 1783
rect 43637 1607 43671 1783
rect 43751 1607 43785 1783
rect 44009 1607 44043 1783
rect 44123 1607 44157 1783
rect 44381 1607 44415 1783
rect 44495 1607 44529 1783
rect 44753 1607 44787 1783
rect 44867 1607 44901 1783
rect 45125 1607 45159 1783
rect 45239 1607 45273 1783
rect 45497 1607 45531 1783
rect 45611 1607 45645 1783
rect 45869 1607 45903 1783
rect 45983 1607 46017 1783
rect 46241 1607 46275 1783
rect 46355 1607 46389 1783
rect 46613 1607 46647 1783
rect 46727 1607 46761 1783
rect 46985 1607 47019 1783
rect 47099 1607 47133 1783
rect 47357 1607 47391 1783
rect 47471 1607 47505 1783
rect 47729 1607 47763 1783
rect 47843 1607 47877 1783
rect 48101 1607 48135 1783
rect 48215 1607 48249 1783
rect 48473 1607 48507 1783
rect 48587 1607 48621 1783
rect 48845 1607 48879 1783
rect 48959 1607 48993 1783
rect 49217 1607 49251 1783
rect 49331 1607 49365 1783
rect 49589 1607 49623 1783
rect 40837 1523 41005 1557
rect 41209 1523 41377 1557
rect 41581 1523 41749 1557
rect 41953 1523 42121 1557
rect 42325 1523 42493 1557
rect 42697 1523 42865 1557
rect 43069 1523 43237 1557
rect 43441 1523 43609 1557
rect 43813 1523 43981 1557
rect 44185 1523 44353 1557
rect 44557 1523 44725 1557
rect 44929 1523 45097 1557
rect 45301 1523 45469 1557
rect 45673 1523 45841 1557
rect 46045 1523 46213 1557
rect 46417 1523 46585 1557
rect 46789 1523 46957 1557
rect 47161 1523 47329 1557
rect 47533 1523 47701 1557
rect 47905 1523 48073 1557
rect 48277 1523 48445 1557
rect 48649 1523 48817 1557
rect 49021 1523 49189 1557
rect 49393 1523 49561 1557
rect 40837 1415 41005 1449
rect 41209 1415 41377 1449
rect 41581 1415 41749 1449
rect 41953 1415 42121 1449
rect 42325 1415 42493 1449
rect 42697 1415 42865 1449
rect 43069 1415 43237 1449
rect 43441 1415 43609 1449
rect 43813 1415 43981 1449
rect 44185 1415 44353 1449
rect 44557 1415 44725 1449
rect 44929 1415 45097 1449
rect 45301 1415 45469 1449
rect 45673 1415 45841 1449
rect 46045 1415 46213 1449
rect 46417 1415 46585 1449
rect 46789 1415 46957 1449
rect 47161 1415 47329 1449
rect 47533 1415 47701 1449
rect 47905 1415 48073 1449
rect 48277 1415 48445 1449
rect 48649 1415 48817 1449
rect 49021 1415 49189 1449
rect 49393 1415 49561 1449
rect 40775 1189 40809 1365
rect 41033 1189 41067 1365
rect 41147 1189 41181 1365
rect 41405 1189 41439 1365
rect 41519 1189 41553 1365
rect 41777 1189 41811 1365
rect 41891 1189 41925 1365
rect 42149 1189 42183 1365
rect 42263 1189 42297 1365
rect 42521 1189 42555 1365
rect 42635 1189 42669 1365
rect 42893 1189 42927 1365
rect 43007 1189 43041 1365
rect 43265 1189 43299 1365
rect 43379 1189 43413 1365
rect 43637 1189 43671 1365
rect 43751 1189 43785 1365
rect 44009 1189 44043 1365
rect 44123 1189 44157 1365
rect 44381 1189 44415 1365
rect 44495 1189 44529 1365
rect 44753 1189 44787 1365
rect 44867 1189 44901 1365
rect 45125 1189 45159 1365
rect 45239 1189 45273 1365
rect 45497 1189 45531 1365
rect 45611 1189 45645 1365
rect 45869 1189 45903 1365
rect 45983 1189 46017 1365
rect 46241 1189 46275 1365
rect 46355 1189 46389 1365
rect 46613 1189 46647 1365
rect 46727 1189 46761 1365
rect 46985 1189 47019 1365
rect 47099 1189 47133 1365
rect 47357 1189 47391 1365
rect 47471 1189 47505 1365
rect 47729 1189 47763 1365
rect 47843 1189 47877 1365
rect 48101 1189 48135 1365
rect 48215 1189 48249 1365
rect 48473 1189 48507 1365
rect 48587 1189 48621 1365
rect 48845 1189 48879 1365
rect 48959 1189 48993 1365
rect 49217 1189 49251 1365
rect 49331 1189 49365 1365
rect 49589 1189 49623 1365
rect 40837 1105 41005 1139
rect 41209 1105 41377 1139
rect 41581 1105 41749 1139
rect 41953 1105 42121 1139
rect 42325 1105 42493 1139
rect 42697 1105 42865 1139
rect 43069 1105 43237 1139
rect 43441 1105 43609 1139
rect 43813 1105 43981 1139
rect 44185 1105 44353 1139
rect 44557 1105 44725 1139
rect 44929 1105 45097 1139
rect 45301 1105 45469 1139
rect 45673 1105 45841 1139
rect 46045 1105 46213 1139
rect 46417 1105 46585 1139
rect 46789 1105 46957 1139
rect 47161 1105 47329 1139
rect 47533 1105 47701 1139
rect 47905 1105 48073 1139
rect 48277 1105 48445 1139
rect 48649 1105 48817 1139
rect 49021 1105 49189 1139
rect 49393 1105 49561 1139
rect 40837 997 41005 1031
rect 41209 997 41377 1031
rect 41581 997 41749 1031
rect 41953 997 42121 1031
rect 42325 997 42493 1031
rect 42697 997 42865 1031
rect 43069 997 43237 1031
rect 43441 997 43609 1031
rect 43813 997 43981 1031
rect 44185 997 44353 1031
rect 44557 997 44725 1031
rect 44929 997 45097 1031
rect 45301 997 45469 1031
rect 45673 997 45841 1031
rect 46045 997 46213 1031
rect 46417 997 46585 1031
rect 46789 997 46957 1031
rect 47161 997 47329 1031
rect 47533 997 47701 1031
rect 47905 997 48073 1031
rect 48277 997 48445 1031
rect 48649 997 48817 1031
rect 49021 997 49189 1031
rect 49393 997 49561 1031
rect 40775 771 40809 947
rect 41033 771 41067 947
rect 41147 771 41181 947
rect 41405 771 41439 947
rect 41519 771 41553 947
rect 41777 771 41811 947
rect 41891 771 41925 947
rect 42149 771 42183 947
rect 42263 771 42297 947
rect 42521 771 42555 947
rect 42635 771 42669 947
rect 42893 771 42927 947
rect 43007 771 43041 947
rect 43265 771 43299 947
rect 43379 771 43413 947
rect 43637 771 43671 947
rect 43751 771 43785 947
rect 44009 771 44043 947
rect 44123 771 44157 947
rect 44381 771 44415 947
rect 44495 771 44529 947
rect 44753 771 44787 947
rect 44867 771 44901 947
rect 45125 771 45159 947
rect 45239 771 45273 947
rect 45497 771 45531 947
rect 45611 771 45645 947
rect 45869 771 45903 947
rect 45983 771 46017 947
rect 46241 771 46275 947
rect 46355 771 46389 947
rect 46613 771 46647 947
rect 46727 771 46761 947
rect 46985 771 47019 947
rect 47099 771 47133 947
rect 47357 771 47391 947
rect 47471 771 47505 947
rect 47729 771 47763 947
rect 47843 771 47877 947
rect 48101 771 48135 947
rect 48215 771 48249 947
rect 48473 771 48507 947
rect 48587 771 48621 947
rect 48845 771 48879 947
rect 48959 771 48993 947
rect 49217 771 49251 947
rect 49331 771 49365 947
rect 49589 771 49623 947
rect 40837 687 41005 721
rect 41209 687 41377 721
rect 41581 687 41749 721
rect 41953 687 42121 721
rect 42325 687 42493 721
rect 42697 687 42865 721
rect 43069 687 43237 721
rect 43441 687 43609 721
rect 43813 687 43981 721
rect 44185 687 44353 721
rect 44557 687 44725 721
rect 44929 687 45097 721
rect 45301 687 45469 721
rect 45673 687 45841 721
rect 46045 687 46213 721
rect 46417 687 46585 721
rect 46789 687 46957 721
rect 47161 687 47329 721
rect 47533 687 47701 721
rect 47905 687 48073 721
rect 48277 687 48445 721
rect 48649 687 48817 721
rect 49021 687 49189 721
rect 49393 687 49561 721
rect 40837 579 41005 613
rect 41209 579 41377 613
rect 41581 579 41749 613
rect 41953 579 42121 613
rect 42325 579 42493 613
rect 42697 579 42865 613
rect 43069 579 43237 613
rect 43441 579 43609 613
rect 43813 579 43981 613
rect 44185 579 44353 613
rect 44557 579 44725 613
rect 44929 579 45097 613
rect 45301 579 45469 613
rect 45673 579 45841 613
rect 46045 579 46213 613
rect 46417 579 46585 613
rect 46789 579 46957 613
rect 47161 579 47329 613
rect 47533 579 47701 613
rect 47905 579 48073 613
rect 48277 579 48445 613
rect 48649 579 48817 613
rect 49021 579 49189 613
rect 49393 579 49561 613
rect 40775 353 40809 529
rect 41033 353 41067 529
rect 41147 353 41181 529
rect 41405 353 41439 529
rect 41519 353 41553 529
rect 41777 353 41811 529
rect 41891 353 41925 529
rect 42149 353 42183 529
rect 42263 353 42297 529
rect 42521 353 42555 529
rect 42635 353 42669 529
rect 42893 353 42927 529
rect 43007 353 43041 529
rect 43265 353 43299 529
rect 43379 353 43413 529
rect 43637 353 43671 529
rect 43751 353 43785 529
rect 44009 353 44043 529
rect 44123 353 44157 529
rect 44381 353 44415 529
rect 44495 353 44529 529
rect 44753 353 44787 529
rect 44867 353 44901 529
rect 45125 353 45159 529
rect 45239 353 45273 529
rect 45497 353 45531 529
rect 45611 353 45645 529
rect 45869 353 45903 529
rect 45983 353 46017 529
rect 46241 353 46275 529
rect 46355 353 46389 529
rect 46613 353 46647 529
rect 46727 353 46761 529
rect 46985 353 47019 529
rect 47099 353 47133 529
rect 47357 353 47391 529
rect 47471 353 47505 529
rect 47729 353 47763 529
rect 47843 353 47877 529
rect 48101 353 48135 529
rect 48215 353 48249 529
rect 48473 353 48507 529
rect 48587 353 48621 529
rect 48845 353 48879 529
rect 48959 353 48993 529
rect 49217 353 49251 529
rect 49331 353 49365 529
rect 49589 353 49623 529
rect 40837 269 41005 303
rect 41209 269 41377 303
rect 41581 269 41749 303
rect 41953 269 42121 303
rect 42325 269 42493 303
rect 42697 269 42865 303
rect 43069 269 43237 303
rect 43441 269 43609 303
rect 43813 269 43981 303
rect 44185 269 44353 303
rect 44557 269 44725 303
rect 44929 269 45097 303
rect 45301 269 45469 303
rect 45673 269 45841 303
rect 46045 269 46213 303
rect 46417 269 46585 303
rect 46789 269 46957 303
rect 47161 269 47329 303
rect 47533 269 47701 303
rect 47905 269 48073 303
rect 48277 269 48445 303
rect 48649 269 48817 303
rect 49021 269 49189 303
rect 49393 269 49561 303
rect 40776 201 40846 212
rect 41444 201 41514 220
rect 42188 201 42258 220
rect 42932 201 43002 220
rect 43676 201 43746 220
rect 44420 201 44490 220
rect 45164 201 45234 220
rect 45908 201 45978 220
rect 46652 201 46722 220
rect 47396 201 47466 220
rect 48140 201 48210 220
rect 48884 201 48954 220
rect 49546 201 49616 216
rect 40776 167 40846 201
rect 41444 167 41514 201
rect 42188 167 42258 201
rect 42932 167 43002 201
rect 43676 167 43746 201
rect 44420 167 44490 201
rect 45164 167 45234 201
rect 45908 167 45978 201
rect 46652 167 46722 201
rect 47396 167 47466 201
rect 48140 167 48210 201
rect 48884 167 48954 201
rect 49546 167 49616 201
rect 40776 142 40846 167
rect 41444 150 41514 167
rect 42188 150 42258 167
rect 42932 150 43002 167
rect 43676 150 43746 167
rect 44420 150 44490 167
rect 45164 150 45234 167
rect 45908 150 45978 167
rect 46652 150 46722 167
rect 47396 150 47466 167
rect 48140 150 48210 167
rect 48884 150 48954 167
rect 49546 146 49616 167
<< metal1 >>
rect 40646 19761 40656 19961
rect 40856 19761 40866 19961
rect 41370 19761 41380 19961
rect 41580 19761 41590 19961
rect 42114 19761 42124 19961
rect 42324 19761 42334 19961
rect 42858 19761 42868 19961
rect 43068 19761 43078 19961
rect 43602 19761 43612 19961
rect 43812 19761 43822 19961
rect 44346 19761 44356 19961
rect 44556 19761 44566 19961
rect 45090 19761 45100 19961
rect 45300 19761 45310 19961
rect 45834 19761 45844 19961
rect 46044 19761 46054 19961
rect 46578 19761 46588 19961
rect 46788 19761 46798 19961
rect 47322 19761 47332 19961
rect 47532 19761 47542 19961
rect 48066 19761 48076 19961
rect 48276 19761 48286 19961
rect 48810 19761 48820 19961
rect 49020 19761 49030 19961
rect 49554 19761 49564 19961
rect 49764 19761 49774 19961
rect 40720 19729 40794 19761
rect 40720 19723 40858 19729
rect 40720 19653 40776 19723
rect 40846 19653 40858 19723
rect 41450 19721 41508 19761
rect 42194 19721 42252 19761
rect 42938 19721 42996 19761
rect 43682 19721 43740 19761
rect 44426 19721 44484 19761
rect 45170 19721 45228 19761
rect 45914 19721 45972 19761
rect 46658 19721 46716 19761
rect 47402 19721 47460 19761
rect 48146 19721 48204 19761
rect 48890 19721 48948 19761
rect 49604 19749 49692 19761
rect 49604 19725 49678 19749
rect 40720 19647 40858 19653
rect 41432 19715 41526 19721
rect 40720 19524 40794 19647
rect 41432 19645 41444 19715
rect 41514 19645 41526 19715
rect 41432 19639 41526 19645
rect 42176 19715 42270 19721
rect 42176 19645 42188 19715
rect 42258 19645 42270 19715
rect 42176 19639 42270 19645
rect 42920 19715 43014 19721
rect 42920 19645 42932 19715
rect 43002 19645 43014 19715
rect 42920 19639 43014 19645
rect 43664 19715 43758 19721
rect 43664 19645 43676 19715
rect 43746 19645 43758 19715
rect 43664 19639 43758 19645
rect 44408 19715 44502 19721
rect 44408 19645 44420 19715
rect 44490 19645 44502 19715
rect 44408 19639 44502 19645
rect 45152 19715 45246 19721
rect 45152 19645 45164 19715
rect 45234 19645 45246 19715
rect 45152 19639 45246 19645
rect 45896 19715 45990 19721
rect 45896 19645 45908 19715
rect 45978 19645 45990 19715
rect 45896 19639 45990 19645
rect 46640 19715 46734 19721
rect 46640 19645 46652 19715
rect 46722 19645 46734 19715
rect 46640 19639 46734 19645
rect 47384 19715 47478 19721
rect 47384 19645 47396 19715
rect 47466 19645 47478 19715
rect 47384 19639 47478 19645
rect 48128 19715 48222 19721
rect 48128 19645 48140 19715
rect 48210 19645 48222 19715
rect 48128 19639 48222 19645
rect 48872 19715 48966 19721
rect 48872 19645 48884 19715
rect 48954 19645 48966 19715
rect 48872 19639 48966 19645
rect 49534 19719 49678 19725
rect 49534 19649 49546 19719
rect 49616 19649 49678 19719
rect 49534 19643 49678 19649
rect 40824 19607 41390 19619
rect 40824 19561 40836 19607
rect 40825 19556 40836 19561
rect 40826 19551 40836 19556
rect 41006 19561 41208 19607
rect 41006 19556 41017 19561
rect 41006 19551 41016 19556
rect 41072 19524 41142 19561
rect 41197 19556 41208 19561
rect 41198 19551 41208 19556
rect 41378 19561 41390 19607
rect 41378 19556 41389 19561
rect 41378 19551 41388 19556
rect 41450 19525 41508 19639
rect 41570 19602 41580 19607
rect 41569 19556 41580 19602
rect 41750 19602 41760 19607
rect 41942 19602 41952 19607
rect 41570 19551 41580 19556
rect 41750 19556 41761 19602
rect 41941 19556 41952 19602
rect 42122 19602 42132 19607
rect 41750 19551 41760 19556
rect 41942 19551 41952 19556
rect 42122 19556 42133 19602
rect 42122 19551 42132 19556
rect 42194 19525 42252 19639
rect 42314 19602 42324 19607
rect 42313 19556 42324 19602
rect 42494 19602 42504 19607
rect 42686 19602 42696 19607
rect 42314 19551 42324 19556
rect 42494 19556 42505 19602
rect 42685 19556 42696 19602
rect 42866 19602 42876 19607
rect 42494 19551 42504 19556
rect 42686 19551 42696 19556
rect 42866 19556 42877 19602
rect 42866 19551 42876 19556
rect 42938 19525 42996 19639
rect 43056 19607 43622 19619
rect 43056 19561 43068 19607
rect 43057 19556 43068 19561
rect 43058 19551 43068 19556
rect 43238 19561 43440 19607
rect 43238 19556 43249 19561
rect 43238 19551 43248 19556
rect 41444 19524 41514 19525
rect 41816 19524 41886 19525
rect 42188 19524 42258 19525
rect 42560 19524 42630 19525
rect 42932 19524 43002 19525
rect 43304 19524 43374 19561
rect 43429 19556 43440 19561
rect 43430 19551 43440 19556
rect 43610 19561 43622 19607
rect 43610 19556 43621 19561
rect 43610 19551 43620 19556
rect 43682 19525 43740 19639
rect 43802 19602 43812 19607
rect 43801 19556 43812 19602
rect 43982 19602 43992 19607
rect 44174 19602 44184 19607
rect 43802 19551 43812 19556
rect 43982 19556 43993 19602
rect 44173 19556 44184 19602
rect 44354 19602 44364 19607
rect 43982 19551 43992 19556
rect 44174 19551 44184 19556
rect 44354 19556 44365 19602
rect 44354 19551 44364 19556
rect 44426 19525 44484 19639
rect 44546 19602 44556 19607
rect 44545 19556 44556 19602
rect 44726 19602 44736 19607
rect 44918 19602 44928 19607
rect 44546 19551 44556 19556
rect 44726 19556 44737 19602
rect 44917 19556 44928 19602
rect 45098 19602 45108 19607
rect 44726 19551 44736 19556
rect 44918 19551 44928 19556
rect 45098 19556 45109 19602
rect 45098 19551 45108 19556
rect 45170 19525 45228 19639
rect 45290 19602 45300 19607
rect 45289 19556 45300 19602
rect 45470 19602 45480 19607
rect 45662 19602 45672 19607
rect 45290 19551 45300 19556
rect 45470 19556 45481 19602
rect 45661 19556 45672 19602
rect 45842 19602 45852 19607
rect 45470 19551 45480 19556
rect 45662 19551 45672 19556
rect 45842 19556 45853 19602
rect 45842 19551 45852 19556
rect 45914 19525 45972 19639
rect 46034 19602 46044 19607
rect 46033 19556 46044 19602
rect 46214 19602 46224 19607
rect 46406 19602 46416 19607
rect 46034 19551 46044 19556
rect 46214 19556 46225 19602
rect 46405 19556 46416 19602
rect 46586 19602 46596 19607
rect 46214 19551 46224 19556
rect 46406 19551 46416 19556
rect 46586 19556 46597 19602
rect 46586 19551 46596 19556
rect 46658 19525 46716 19639
rect 46778 19602 46788 19607
rect 46777 19556 46788 19602
rect 46958 19602 46968 19607
rect 47150 19602 47160 19607
rect 46778 19551 46788 19556
rect 46958 19556 46969 19602
rect 47149 19556 47160 19602
rect 47330 19602 47340 19607
rect 46958 19551 46968 19556
rect 47150 19551 47160 19556
rect 47330 19556 47341 19602
rect 47330 19551 47340 19556
rect 47402 19525 47460 19639
rect 47522 19602 47532 19607
rect 47521 19556 47532 19602
rect 47702 19602 47712 19607
rect 47894 19602 47904 19607
rect 47522 19551 47532 19556
rect 47702 19556 47713 19602
rect 47893 19556 47904 19602
rect 48074 19602 48084 19607
rect 47702 19551 47712 19556
rect 47894 19551 47904 19556
rect 48074 19556 48085 19602
rect 48074 19551 48084 19556
rect 48146 19525 48204 19639
rect 48266 19602 48276 19607
rect 48265 19556 48276 19602
rect 48446 19602 48456 19607
rect 48638 19602 48648 19607
rect 48266 19551 48276 19556
rect 48446 19556 48457 19602
rect 48637 19556 48648 19602
rect 48818 19602 48828 19607
rect 48446 19551 48456 19556
rect 48638 19551 48648 19556
rect 48818 19556 48829 19602
rect 48818 19551 48828 19556
rect 48890 19525 48948 19639
rect 49010 19602 49020 19607
rect 49009 19556 49020 19602
rect 49190 19602 49200 19607
rect 49382 19602 49392 19607
rect 49010 19551 49020 19556
rect 49190 19556 49201 19602
rect 49381 19556 49392 19602
rect 49562 19602 49572 19607
rect 49190 19551 49200 19556
rect 49382 19551 49392 19556
rect 49562 19556 49573 19602
rect 49562 19551 49572 19556
rect 43676 19524 43746 19525
rect 44048 19524 44118 19525
rect 44420 19524 44490 19525
rect 44792 19524 44862 19525
rect 45164 19524 45234 19525
rect 45536 19524 45606 19525
rect 45908 19524 45978 19525
rect 46280 19524 46350 19525
rect 46652 19524 46722 19525
rect 47024 19524 47094 19525
rect 47396 19524 47466 19525
rect 47768 19524 47838 19525
rect 48140 19524 48210 19525
rect 48512 19524 48582 19525
rect 48884 19524 48954 19525
rect 49256 19524 49326 19525
rect 49604 19524 49678 19643
rect 40720 19512 40815 19524
rect 40720 19336 40775 19512
rect 40809 19336 40815 19512
rect 40720 19324 40815 19336
rect 41027 19512 41187 19524
rect 41027 19336 41033 19512
rect 41067 19336 41147 19512
rect 41181 19336 41187 19512
rect 41027 19324 41187 19336
rect 41399 19512 41559 19524
rect 41399 19336 41405 19512
rect 41439 19336 41519 19512
rect 41553 19336 41559 19512
rect 41399 19324 41559 19336
rect 41771 19512 41931 19524
rect 41771 19336 41777 19512
rect 41811 19336 41891 19512
rect 41925 19336 41931 19512
rect 41771 19324 41931 19336
rect 42143 19512 42303 19524
rect 42143 19336 42149 19512
rect 42183 19336 42263 19512
rect 42297 19336 42303 19512
rect 42143 19324 42303 19336
rect 42515 19512 42675 19524
rect 42515 19336 42521 19512
rect 42555 19336 42635 19512
rect 42669 19336 42675 19512
rect 42515 19324 42675 19336
rect 42887 19512 43047 19524
rect 42887 19336 42893 19512
rect 42927 19336 43007 19512
rect 43041 19336 43047 19512
rect 42887 19324 43047 19336
rect 43259 19512 43419 19524
rect 43259 19336 43265 19512
rect 43299 19336 43379 19512
rect 43413 19336 43419 19512
rect 43259 19324 43419 19336
rect 43631 19512 43791 19524
rect 43631 19336 43637 19512
rect 43671 19336 43751 19512
rect 43785 19336 43791 19512
rect 43631 19324 43791 19336
rect 44003 19512 44163 19524
rect 44003 19336 44009 19512
rect 44043 19336 44123 19512
rect 44157 19336 44163 19512
rect 44003 19324 44163 19336
rect 44375 19512 44535 19524
rect 44375 19336 44381 19512
rect 44415 19336 44495 19512
rect 44529 19336 44535 19512
rect 44375 19324 44535 19336
rect 44747 19512 44907 19524
rect 44747 19336 44753 19512
rect 44787 19336 44867 19512
rect 44901 19336 44907 19512
rect 44747 19324 44907 19336
rect 45119 19512 45279 19524
rect 45119 19336 45125 19512
rect 45159 19336 45239 19512
rect 45273 19336 45279 19512
rect 45119 19324 45279 19336
rect 45491 19512 45651 19524
rect 45491 19336 45497 19512
rect 45531 19336 45611 19512
rect 45645 19336 45651 19512
rect 45491 19324 45651 19336
rect 45863 19512 46023 19524
rect 45863 19336 45869 19512
rect 45903 19336 45983 19512
rect 46017 19336 46023 19512
rect 45863 19324 46023 19336
rect 46235 19512 46395 19524
rect 46235 19336 46241 19512
rect 46275 19336 46355 19512
rect 46389 19336 46395 19512
rect 46235 19324 46395 19336
rect 46607 19512 46767 19524
rect 46607 19336 46613 19512
rect 46647 19336 46727 19512
rect 46761 19336 46767 19512
rect 46607 19324 46767 19336
rect 46979 19512 47139 19524
rect 46979 19336 46985 19512
rect 47019 19336 47099 19512
rect 47133 19336 47139 19512
rect 46979 19324 47139 19336
rect 47351 19512 47511 19524
rect 47351 19336 47357 19512
rect 47391 19336 47471 19512
rect 47505 19336 47511 19512
rect 47351 19324 47511 19336
rect 47723 19512 47883 19524
rect 47723 19336 47729 19512
rect 47763 19336 47843 19512
rect 47877 19336 47883 19512
rect 47723 19324 47883 19336
rect 48095 19512 48255 19524
rect 48095 19336 48101 19512
rect 48135 19336 48215 19512
rect 48249 19336 48255 19512
rect 48095 19324 48255 19336
rect 48467 19512 48627 19524
rect 48467 19336 48473 19512
rect 48507 19336 48587 19512
rect 48621 19336 48627 19512
rect 48467 19324 48627 19336
rect 48839 19512 48999 19524
rect 48839 19336 48845 19512
rect 48879 19336 48959 19512
rect 48993 19336 48999 19512
rect 48839 19324 48999 19336
rect 49211 19512 49371 19524
rect 49211 19336 49217 19512
rect 49251 19336 49331 19512
rect 49365 19336 49371 19512
rect 49211 19324 49371 19336
rect 49583 19512 49678 19524
rect 49583 19336 49589 19512
rect 49623 19336 49678 19512
rect 49583 19324 49678 19336
rect 40720 19106 40794 19324
rect 41072 19293 41142 19324
rect 40824 19287 41390 19293
rect 40824 19143 40836 19287
rect 41006 19143 41208 19287
rect 41378 19143 41390 19287
rect 40824 19137 41390 19143
rect 41072 19106 41142 19137
rect 41444 19106 41514 19324
rect 41569 19287 41761 19292
rect 41569 19246 41580 19287
rect 41570 19184 41580 19246
rect 41569 19143 41580 19184
rect 41750 19246 41761 19287
rect 41750 19184 41760 19246
rect 41750 19143 41761 19184
rect 41569 19138 41761 19143
rect 41816 19106 41886 19324
rect 41941 19287 42133 19292
rect 41941 19246 41952 19287
rect 41942 19184 41952 19246
rect 41941 19143 41952 19184
rect 42122 19246 42133 19287
rect 42122 19184 42132 19246
rect 42122 19143 42133 19184
rect 41941 19138 42133 19143
rect 42188 19106 42258 19324
rect 42313 19287 42505 19292
rect 42313 19246 42324 19287
rect 42314 19184 42324 19246
rect 42313 19143 42324 19184
rect 42494 19246 42505 19287
rect 42494 19184 42504 19246
rect 42494 19143 42505 19184
rect 42313 19138 42505 19143
rect 42560 19106 42630 19324
rect 42685 19287 42877 19292
rect 42685 19246 42696 19287
rect 42686 19184 42696 19246
rect 42685 19143 42696 19184
rect 42866 19246 42877 19287
rect 42866 19184 42876 19246
rect 42866 19143 42877 19184
rect 42685 19138 42877 19143
rect 42932 19106 43002 19324
rect 43304 19293 43374 19324
rect 43056 19287 43622 19293
rect 43056 19143 43068 19287
rect 43238 19143 43440 19287
rect 43610 19143 43622 19287
rect 43056 19137 43622 19143
rect 43304 19106 43374 19137
rect 43676 19106 43746 19324
rect 43801 19287 43993 19292
rect 43801 19246 43812 19287
rect 43802 19184 43812 19246
rect 43801 19143 43812 19184
rect 43982 19246 43993 19287
rect 43982 19184 43992 19246
rect 43982 19143 43993 19184
rect 43801 19138 43993 19143
rect 44048 19106 44118 19324
rect 44173 19287 44365 19292
rect 44173 19246 44184 19287
rect 44174 19184 44184 19246
rect 44173 19143 44184 19184
rect 44354 19246 44365 19287
rect 44354 19184 44364 19246
rect 44354 19143 44365 19184
rect 44173 19138 44365 19143
rect 44420 19106 44490 19324
rect 44545 19287 44737 19292
rect 44545 19246 44556 19287
rect 44546 19184 44556 19246
rect 44545 19143 44556 19184
rect 44726 19246 44737 19287
rect 44726 19184 44736 19246
rect 44726 19143 44737 19184
rect 44545 19138 44737 19143
rect 44792 19106 44862 19324
rect 44917 19287 45109 19292
rect 44917 19246 44928 19287
rect 44918 19184 44928 19246
rect 44917 19143 44928 19184
rect 45098 19246 45109 19287
rect 45098 19184 45108 19246
rect 45098 19143 45109 19184
rect 44917 19138 45109 19143
rect 45164 19106 45234 19324
rect 45289 19287 45481 19292
rect 45289 19246 45300 19287
rect 45290 19184 45300 19246
rect 45289 19143 45300 19184
rect 45470 19246 45481 19287
rect 45470 19184 45480 19246
rect 45470 19143 45481 19184
rect 45289 19138 45481 19143
rect 45536 19106 45606 19324
rect 45661 19287 45853 19292
rect 45661 19246 45672 19287
rect 45662 19184 45672 19246
rect 45661 19143 45672 19184
rect 45842 19246 45853 19287
rect 45842 19184 45852 19246
rect 45842 19143 45853 19184
rect 45661 19138 45853 19143
rect 45908 19106 45978 19324
rect 46033 19287 46225 19292
rect 46033 19246 46044 19287
rect 46034 19184 46044 19246
rect 46033 19143 46044 19184
rect 46214 19246 46225 19287
rect 46214 19184 46224 19246
rect 46214 19143 46225 19184
rect 46033 19138 46225 19143
rect 46280 19106 46350 19324
rect 46405 19287 46597 19292
rect 46405 19246 46416 19287
rect 46406 19184 46416 19246
rect 46405 19143 46416 19184
rect 46586 19246 46597 19287
rect 46586 19184 46596 19246
rect 46586 19143 46597 19184
rect 46405 19138 46597 19143
rect 46652 19106 46722 19324
rect 46777 19287 46969 19292
rect 46777 19246 46788 19287
rect 46778 19184 46788 19246
rect 46777 19143 46788 19184
rect 46958 19246 46969 19287
rect 46958 19184 46968 19246
rect 46958 19143 46969 19184
rect 46777 19138 46969 19143
rect 47024 19106 47094 19324
rect 47149 19287 47341 19292
rect 47149 19246 47160 19287
rect 47150 19184 47160 19246
rect 47149 19143 47160 19184
rect 47330 19246 47341 19287
rect 47330 19184 47340 19246
rect 47330 19143 47341 19184
rect 47149 19138 47341 19143
rect 47396 19106 47466 19324
rect 47521 19287 47713 19292
rect 47521 19246 47532 19287
rect 47522 19184 47532 19246
rect 47521 19143 47532 19184
rect 47702 19246 47713 19287
rect 47702 19184 47712 19246
rect 47702 19143 47713 19184
rect 47521 19138 47713 19143
rect 47768 19106 47838 19324
rect 47893 19287 48085 19292
rect 47893 19246 47904 19287
rect 47894 19184 47904 19246
rect 47893 19143 47904 19184
rect 48074 19246 48085 19287
rect 48074 19184 48084 19246
rect 48074 19143 48085 19184
rect 47893 19138 48085 19143
rect 48140 19106 48210 19324
rect 48265 19287 48457 19292
rect 48265 19246 48276 19287
rect 48266 19184 48276 19246
rect 48265 19143 48276 19184
rect 48446 19246 48457 19287
rect 48446 19184 48456 19246
rect 48446 19143 48457 19184
rect 48265 19138 48457 19143
rect 48512 19106 48582 19324
rect 48637 19287 48829 19292
rect 48637 19246 48648 19287
rect 48638 19184 48648 19246
rect 48637 19143 48648 19184
rect 48818 19246 48829 19287
rect 48818 19184 48828 19246
rect 48818 19143 48829 19184
rect 48637 19138 48829 19143
rect 48884 19106 48954 19324
rect 49009 19287 49201 19292
rect 49009 19246 49020 19287
rect 49010 19184 49020 19246
rect 49009 19143 49020 19184
rect 49190 19246 49201 19287
rect 49190 19184 49200 19246
rect 49190 19143 49201 19184
rect 49009 19138 49201 19143
rect 49256 19106 49326 19324
rect 49381 19287 49573 19292
rect 49381 19246 49392 19287
rect 49382 19184 49392 19246
rect 49381 19143 49392 19184
rect 49562 19246 49573 19287
rect 49562 19184 49572 19246
rect 49562 19143 49573 19184
rect 49381 19138 49573 19143
rect 49604 19106 49678 19324
rect 40720 19094 40815 19106
rect 40720 18918 40775 19094
rect 40809 18918 40815 19094
rect 40720 18906 40815 18918
rect 41027 19094 41187 19106
rect 41027 18918 41033 19094
rect 41067 18918 41147 19094
rect 41181 18918 41187 19094
rect 41027 18906 41187 18918
rect 41399 19094 41559 19106
rect 41399 18918 41405 19094
rect 41439 18918 41519 19094
rect 41553 18918 41559 19094
rect 41399 18906 41559 18918
rect 41771 19094 41931 19106
rect 41771 18918 41777 19094
rect 41811 18918 41891 19094
rect 41925 18918 41931 19094
rect 41771 18906 41931 18918
rect 42143 19094 42303 19106
rect 42143 18918 42149 19094
rect 42183 18918 42263 19094
rect 42297 18918 42303 19094
rect 42143 18906 42303 18918
rect 42515 19094 42675 19106
rect 42515 18918 42521 19094
rect 42555 18918 42635 19094
rect 42669 18918 42675 19094
rect 42515 18906 42675 18918
rect 42887 19094 43047 19106
rect 42887 18918 42893 19094
rect 42927 18918 43007 19094
rect 43041 18918 43047 19094
rect 42887 18906 43047 18918
rect 43259 19094 43419 19106
rect 43259 18918 43265 19094
rect 43299 18918 43379 19094
rect 43413 18918 43419 19094
rect 43259 18906 43419 18918
rect 43631 19094 43791 19106
rect 43631 18918 43637 19094
rect 43671 18918 43751 19094
rect 43785 18918 43791 19094
rect 43631 18906 43791 18918
rect 44003 19094 44163 19106
rect 44003 18918 44009 19094
rect 44043 18918 44123 19094
rect 44157 18918 44163 19094
rect 44003 18906 44163 18918
rect 44375 19094 44535 19106
rect 44375 18918 44381 19094
rect 44415 18918 44495 19094
rect 44529 18918 44535 19094
rect 44375 18906 44535 18918
rect 44747 19094 44907 19106
rect 44747 18918 44753 19094
rect 44787 18918 44867 19094
rect 44901 18918 44907 19094
rect 44747 18906 44907 18918
rect 45119 19094 45279 19106
rect 45119 18918 45125 19094
rect 45159 18918 45239 19094
rect 45273 18918 45279 19094
rect 45119 18906 45279 18918
rect 45491 19094 45651 19106
rect 45491 18918 45497 19094
rect 45531 18918 45611 19094
rect 45645 18918 45651 19094
rect 45491 18906 45651 18918
rect 45863 19094 46023 19106
rect 45863 18918 45869 19094
rect 45903 18918 45983 19094
rect 46017 18918 46023 19094
rect 45863 18906 46023 18918
rect 46235 19094 46395 19106
rect 46235 18918 46241 19094
rect 46275 18918 46355 19094
rect 46389 18918 46395 19094
rect 46235 18906 46395 18918
rect 46607 19094 46767 19106
rect 46607 18918 46613 19094
rect 46647 18918 46727 19094
rect 46761 18918 46767 19094
rect 46607 18906 46767 18918
rect 46979 19094 47139 19106
rect 46979 18918 46985 19094
rect 47019 18918 47099 19094
rect 47133 18918 47139 19094
rect 46979 18906 47139 18918
rect 47351 19094 47511 19106
rect 47351 18918 47357 19094
rect 47391 18918 47471 19094
rect 47505 18918 47511 19094
rect 47351 18906 47511 18918
rect 47723 19094 47883 19106
rect 47723 18918 47729 19094
rect 47763 18918 47843 19094
rect 47877 18918 47883 19094
rect 47723 18906 47883 18918
rect 48095 19094 48255 19106
rect 48095 18918 48101 19094
rect 48135 18918 48215 19094
rect 48249 18918 48255 19094
rect 48095 18906 48255 18918
rect 48467 19094 48627 19106
rect 48467 18918 48473 19094
rect 48507 18918 48587 19094
rect 48621 18918 48627 19094
rect 48467 18906 48627 18918
rect 48839 19094 48999 19106
rect 48839 18918 48845 19094
rect 48879 18918 48959 19094
rect 48993 18918 48999 19094
rect 48839 18906 48999 18918
rect 49211 19094 49371 19106
rect 49211 18918 49217 19094
rect 49251 18918 49331 19094
rect 49365 18918 49371 19094
rect 49211 18906 49371 18918
rect 49583 19094 49678 19106
rect 49583 18918 49589 19094
rect 49623 18918 49678 19094
rect 49583 18906 49678 18918
rect 40720 18688 40794 18906
rect 41072 18875 41142 18906
rect 40824 18869 41390 18875
rect 40824 18725 40836 18869
rect 41006 18725 41208 18869
rect 41378 18725 41390 18869
rect 40824 18719 41390 18725
rect 41072 18688 41142 18719
rect 41444 18688 41514 18906
rect 41569 18869 41761 18874
rect 41569 18828 41580 18869
rect 41570 18766 41580 18828
rect 41569 18725 41580 18766
rect 41750 18828 41761 18869
rect 41750 18766 41760 18828
rect 41750 18725 41761 18766
rect 41569 18720 41761 18725
rect 41816 18688 41886 18906
rect 41941 18869 42133 18874
rect 41941 18828 41952 18869
rect 41942 18766 41952 18828
rect 41941 18725 41952 18766
rect 42122 18828 42133 18869
rect 42122 18766 42132 18828
rect 42122 18725 42133 18766
rect 41941 18720 42133 18725
rect 42188 18688 42258 18906
rect 42313 18869 42505 18874
rect 42313 18828 42324 18869
rect 42314 18766 42324 18828
rect 42313 18725 42324 18766
rect 42494 18828 42505 18869
rect 42494 18766 42504 18828
rect 42494 18725 42505 18766
rect 42313 18720 42505 18725
rect 42560 18688 42630 18906
rect 42685 18869 42877 18874
rect 42685 18828 42696 18869
rect 42686 18766 42696 18828
rect 42685 18725 42696 18766
rect 42866 18828 42877 18869
rect 42866 18766 42876 18828
rect 42866 18725 42877 18766
rect 42685 18720 42877 18725
rect 42932 18688 43002 18906
rect 43304 18875 43374 18906
rect 43056 18869 43622 18875
rect 43056 18725 43068 18869
rect 43238 18725 43440 18869
rect 43610 18725 43622 18869
rect 43056 18719 43622 18725
rect 43304 18688 43374 18719
rect 43676 18688 43746 18906
rect 43801 18869 43993 18874
rect 43801 18828 43812 18869
rect 43802 18766 43812 18828
rect 43801 18725 43812 18766
rect 43982 18828 43993 18869
rect 43982 18766 43992 18828
rect 43982 18725 43993 18766
rect 43801 18720 43993 18725
rect 44048 18688 44118 18906
rect 44173 18869 44365 18874
rect 44173 18828 44184 18869
rect 44174 18766 44184 18828
rect 44173 18725 44184 18766
rect 44354 18828 44365 18869
rect 44354 18766 44364 18828
rect 44354 18725 44365 18766
rect 44173 18720 44365 18725
rect 44420 18688 44490 18906
rect 44545 18869 44737 18874
rect 44545 18828 44556 18869
rect 44546 18766 44556 18828
rect 44545 18725 44556 18766
rect 44726 18828 44737 18869
rect 44726 18766 44736 18828
rect 44726 18725 44737 18766
rect 44545 18720 44737 18725
rect 44792 18688 44862 18906
rect 44917 18869 45109 18874
rect 44917 18828 44928 18869
rect 44918 18766 44928 18828
rect 44917 18725 44928 18766
rect 45098 18828 45109 18869
rect 45098 18766 45108 18828
rect 45098 18725 45109 18766
rect 44917 18720 45109 18725
rect 45164 18688 45234 18906
rect 45289 18869 45481 18874
rect 45289 18828 45300 18869
rect 45290 18766 45300 18828
rect 45289 18725 45300 18766
rect 45470 18828 45481 18869
rect 45470 18766 45480 18828
rect 45470 18725 45481 18766
rect 45289 18720 45481 18725
rect 45536 18688 45606 18906
rect 45661 18869 45853 18874
rect 45661 18828 45672 18869
rect 45662 18766 45672 18828
rect 45661 18725 45672 18766
rect 45842 18828 45853 18869
rect 45842 18766 45852 18828
rect 45842 18725 45853 18766
rect 45661 18720 45853 18725
rect 45908 18688 45978 18906
rect 46033 18869 46225 18874
rect 46033 18828 46044 18869
rect 46034 18766 46044 18828
rect 46033 18725 46044 18766
rect 46214 18828 46225 18869
rect 46214 18766 46224 18828
rect 46214 18725 46225 18766
rect 46033 18720 46225 18725
rect 46280 18688 46350 18906
rect 46405 18869 46597 18874
rect 46405 18828 46416 18869
rect 46406 18766 46416 18828
rect 46405 18725 46416 18766
rect 46586 18828 46597 18869
rect 46586 18766 46596 18828
rect 46586 18725 46597 18766
rect 46405 18720 46597 18725
rect 46652 18688 46722 18906
rect 46777 18869 46969 18874
rect 46777 18828 46788 18869
rect 46778 18766 46788 18828
rect 46777 18725 46788 18766
rect 46958 18828 46969 18869
rect 46958 18766 46968 18828
rect 46958 18725 46969 18766
rect 46777 18720 46969 18725
rect 47024 18688 47094 18906
rect 47149 18869 47341 18874
rect 47149 18828 47160 18869
rect 47150 18766 47160 18828
rect 47149 18725 47160 18766
rect 47330 18828 47341 18869
rect 47330 18766 47340 18828
rect 47330 18725 47341 18766
rect 47149 18720 47341 18725
rect 47396 18688 47466 18906
rect 47521 18869 47713 18874
rect 47521 18828 47532 18869
rect 47522 18766 47532 18828
rect 47521 18725 47532 18766
rect 47702 18828 47713 18869
rect 47702 18766 47712 18828
rect 47702 18725 47713 18766
rect 47521 18720 47713 18725
rect 47768 18688 47838 18906
rect 47893 18869 48085 18874
rect 47893 18828 47904 18869
rect 47894 18766 47904 18828
rect 47893 18725 47904 18766
rect 48074 18828 48085 18869
rect 48074 18766 48084 18828
rect 48074 18725 48085 18766
rect 47893 18720 48085 18725
rect 48140 18688 48210 18906
rect 48265 18869 48457 18874
rect 48265 18828 48276 18869
rect 48266 18766 48276 18828
rect 48265 18725 48276 18766
rect 48446 18828 48457 18869
rect 48446 18766 48456 18828
rect 48446 18725 48457 18766
rect 48265 18720 48457 18725
rect 48512 18688 48582 18906
rect 48637 18869 48829 18874
rect 48637 18828 48648 18869
rect 48638 18766 48648 18828
rect 48637 18725 48648 18766
rect 48818 18828 48829 18869
rect 48818 18766 48828 18828
rect 48818 18725 48829 18766
rect 48637 18720 48829 18725
rect 48884 18688 48954 18906
rect 49009 18869 49201 18874
rect 49009 18828 49020 18869
rect 49010 18766 49020 18828
rect 49009 18725 49020 18766
rect 49190 18828 49201 18869
rect 49190 18766 49200 18828
rect 49190 18725 49201 18766
rect 49009 18720 49201 18725
rect 49256 18688 49326 18906
rect 49381 18869 49573 18874
rect 49381 18828 49392 18869
rect 49382 18766 49392 18828
rect 49381 18725 49392 18766
rect 49562 18828 49573 18869
rect 49562 18766 49572 18828
rect 49562 18725 49573 18766
rect 49381 18720 49573 18725
rect 49604 18688 49678 18906
rect 40720 18676 40815 18688
rect 40720 18500 40775 18676
rect 40809 18500 40815 18676
rect 40720 18488 40815 18500
rect 41027 18676 41187 18688
rect 41027 18500 41033 18676
rect 41067 18500 41147 18676
rect 41181 18500 41187 18676
rect 41027 18488 41187 18500
rect 41399 18676 41559 18688
rect 41399 18500 41405 18676
rect 41439 18500 41519 18676
rect 41553 18500 41559 18676
rect 41399 18488 41559 18500
rect 41771 18676 41931 18688
rect 41771 18500 41777 18676
rect 41811 18500 41891 18676
rect 41925 18500 41931 18676
rect 41771 18488 41931 18500
rect 42143 18676 42303 18688
rect 42143 18500 42149 18676
rect 42183 18500 42263 18676
rect 42297 18500 42303 18676
rect 42143 18488 42303 18500
rect 42515 18676 42675 18688
rect 42515 18500 42521 18676
rect 42555 18500 42635 18676
rect 42669 18500 42675 18676
rect 42515 18488 42675 18500
rect 42887 18676 43047 18688
rect 42887 18500 42893 18676
rect 42927 18500 43007 18676
rect 43041 18500 43047 18676
rect 42887 18488 43047 18500
rect 43259 18676 43419 18688
rect 43259 18500 43265 18676
rect 43299 18500 43379 18676
rect 43413 18500 43419 18676
rect 43259 18488 43419 18500
rect 43631 18676 43791 18688
rect 43631 18500 43637 18676
rect 43671 18500 43751 18676
rect 43785 18500 43791 18676
rect 43631 18488 43791 18500
rect 44003 18676 44163 18688
rect 44003 18500 44009 18676
rect 44043 18500 44123 18676
rect 44157 18500 44163 18676
rect 44003 18488 44163 18500
rect 44375 18676 44535 18688
rect 44375 18500 44381 18676
rect 44415 18500 44495 18676
rect 44529 18500 44535 18676
rect 44375 18488 44535 18500
rect 44747 18676 44907 18688
rect 44747 18500 44753 18676
rect 44787 18500 44867 18676
rect 44901 18500 44907 18676
rect 44747 18488 44907 18500
rect 45119 18676 45279 18688
rect 45119 18500 45125 18676
rect 45159 18500 45239 18676
rect 45273 18500 45279 18676
rect 45119 18488 45279 18500
rect 45491 18676 45651 18688
rect 45491 18500 45497 18676
rect 45531 18500 45611 18676
rect 45645 18500 45651 18676
rect 45491 18488 45651 18500
rect 45863 18676 46023 18688
rect 45863 18500 45869 18676
rect 45903 18500 45983 18676
rect 46017 18500 46023 18676
rect 45863 18488 46023 18500
rect 46235 18676 46395 18688
rect 46235 18500 46241 18676
rect 46275 18500 46355 18676
rect 46389 18500 46395 18676
rect 46235 18488 46395 18500
rect 46607 18676 46767 18688
rect 46607 18500 46613 18676
rect 46647 18500 46727 18676
rect 46761 18500 46767 18676
rect 46607 18488 46767 18500
rect 46979 18676 47139 18688
rect 46979 18500 46985 18676
rect 47019 18500 47099 18676
rect 47133 18500 47139 18676
rect 46979 18488 47139 18500
rect 47351 18676 47511 18688
rect 47351 18500 47357 18676
rect 47391 18500 47471 18676
rect 47505 18500 47511 18676
rect 47351 18488 47511 18500
rect 47723 18676 47883 18688
rect 47723 18500 47729 18676
rect 47763 18500 47843 18676
rect 47877 18500 47883 18676
rect 47723 18488 47883 18500
rect 48095 18676 48255 18688
rect 48095 18500 48101 18676
rect 48135 18500 48215 18676
rect 48249 18500 48255 18676
rect 48095 18488 48255 18500
rect 48467 18676 48627 18688
rect 48467 18500 48473 18676
rect 48507 18500 48587 18676
rect 48621 18500 48627 18676
rect 48467 18488 48627 18500
rect 48839 18676 48999 18688
rect 48839 18500 48845 18676
rect 48879 18500 48959 18676
rect 48993 18500 48999 18676
rect 48839 18488 48999 18500
rect 49211 18676 49371 18688
rect 49211 18500 49217 18676
rect 49251 18500 49331 18676
rect 49365 18500 49371 18676
rect 49211 18488 49371 18500
rect 49583 18676 49678 18688
rect 49583 18500 49589 18676
rect 49623 18500 49678 18676
rect 49583 18488 49678 18500
rect 40720 18270 40794 18488
rect 41072 18457 41142 18488
rect 40824 18451 41390 18457
rect 40824 18307 40836 18451
rect 41006 18307 41208 18451
rect 41378 18307 41390 18451
rect 40824 18301 41390 18307
rect 41072 18270 41142 18301
rect 41444 18270 41514 18488
rect 41569 18451 41761 18456
rect 41569 18410 41580 18451
rect 41570 18348 41580 18410
rect 41569 18307 41580 18348
rect 41750 18410 41761 18451
rect 41750 18348 41760 18410
rect 41750 18307 41761 18348
rect 41569 18302 41761 18307
rect 41816 18270 41886 18488
rect 41941 18451 42133 18456
rect 41941 18410 41952 18451
rect 41942 18348 41952 18410
rect 41941 18307 41952 18348
rect 42122 18410 42133 18451
rect 42122 18348 42132 18410
rect 42122 18307 42133 18348
rect 41941 18302 42133 18307
rect 42188 18270 42258 18488
rect 42313 18451 42505 18456
rect 42313 18410 42324 18451
rect 42314 18348 42324 18410
rect 42313 18307 42324 18348
rect 42494 18410 42505 18451
rect 42494 18348 42504 18410
rect 42494 18307 42505 18348
rect 42313 18302 42505 18307
rect 42560 18270 42630 18488
rect 42685 18451 42877 18456
rect 42685 18410 42696 18451
rect 42686 18348 42696 18410
rect 42685 18307 42696 18348
rect 42866 18410 42877 18451
rect 42866 18348 42876 18410
rect 42866 18307 42877 18348
rect 42685 18302 42877 18307
rect 42932 18270 43002 18488
rect 43304 18457 43374 18488
rect 43056 18451 43622 18457
rect 43056 18307 43068 18451
rect 43238 18307 43440 18451
rect 43610 18307 43622 18451
rect 43056 18301 43622 18307
rect 43304 18270 43374 18301
rect 43676 18270 43746 18488
rect 43801 18451 43993 18456
rect 43801 18410 43812 18451
rect 43802 18348 43812 18410
rect 43801 18307 43812 18348
rect 43982 18410 43993 18451
rect 43982 18348 43992 18410
rect 43982 18307 43993 18348
rect 43801 18302 43993 18307
rect 44048 18270 44118 18488
rect 44173 18451 44365 18456
rect 44173 18410 44184 18451
rect 44174 18348 44184 18410
rect 44173 18307 44184 18348
rect 44354 18410 44365 18451
rect 44354 18348 44364 18410
rect 44354 18307 44365 18348
rect 44173 18302 44365 18307
rect 44420 18270 44490 18488
rect 44545 18451 44737 18456
rect 44545 18410 44556 18451
rect 44546 18348 44556 18410
rect 44545 18307 44556 18348
rect 44726 18410 44737 18451
rect 44726 18348 44736 18410
rect 44726 18307 44737 18348
rect 44545 18302 44737 18307
rect 44792 18270 44862 18488
rect 44917 18451 45109 18456
rect 44917 18410 44928 18451
rect 44918 18348 44928 18410
rect 44917 18307 44928 18348
rect 45098 18410 45109 18451
rect 45098 18348 45108 18410
rect 45098 18307 45109 18348
rect 44917 18302 45109 18307
rect 45164 18270 45234 18488
rect 45289 18451 45481 18456
rect 45289 18410 45300 18451
rect 45290 18348 45300 18410
rect 45289 18307 45300 18348
rect 45470 18410 45481 18451
rect 45470 18348 45480 18410
rect 45470 18307 45481 18348
rect 45289 18302 45481 18307
rect 45536 18270 45606 18488
rect 45661 18451 45853 18456
rect 45661 18410 45672 18451
rect 45662 18348 45672 18410
rect 45661 18307 45672 18348
rect 45842 18410 45853 18451
rect 45842 18348 45852 18410
rect 45842 18307 45853 18348
rect 45661 18302 45853 18307
rect 45908 18270 45978 18488
rect 46033 18451 46225 18456
rect 46033 18410 46044 18451
rect 46034 18348 46044 18410
rect 46033 18307 46044 18348
rect 46214 18410 46225 18451
rect 46214 18348 46224 18410
rect 46214 18307 46225 18348
rect 46033 18302 46225 18307
rect 46280 18270 46350 18488
rect 46405 18451 46597 18456
rect 46405 18410 46416 18451
rect 46406 18348 46416 18410
rect 46405 18307 46416 18348
rect 46586 18410 46597 18451
rect 46586 18348 46596 18410
rect 46586 18307 46597 18348
rect 46405 18302 46597 18307
rect 46652 18270 46722 18488
rect 46777 18451 46969 18456
rect 46777 18410 46788 18451
rect 46778 18348 46788 18410
rect 46777 18307 46788 18348
rect 46958 18410 46969 18451
rect 46958 18348 46968 18410
rect 46958 18307 46969 18348
rect 46777 18302 46969 18307
rect 47024 18270 47094 18488
rect 47149 18451 47341 18456
rect 47149 18410 47160 18451
rect 47150 18348 47160 18410
rect 47149 18307 47160 18348
rect 47330 18410 47341 18451
rect 47330 18348 47340 18410
rect 47330 18307 47341 18348
rect 47149 18302 47341 18307
rect 47396 18270 47466 18488
rect 47521 18451 47713 18456
rect 47521 18410 47532 18451
rect 47522 18348 47532 18410
rect 47521 18307 47532 18348
rect 47702 18410 47713 18451
rect 47702 18348 47712 18410
rect 47702 18307 47713 18348
rect 47521 18302 47713 18307
rect 47768 18270 47838 18488
rect 47893 18451 48085 18456
rect 47893 18410 47904 18451
rect 47894 18348 47904 18410
rect 47893 18307 47904 18348
rect 48074 18410 48085 18451
rect 48074 18348 48084 18410
rect 48074 18307 48085 18348
rect 47893 18302 48085 18307
rect 48140 18270 48210 18488
rect 48265 18451 48457 18456
rect 48265 18410 48276 18451
rect 48266 18348 48276 18410
rect 48265 18307 48276 18348
rect 48446 18410 48457 18451
rect 48446 18348 48456 18410
rect 48446 18307 48457 18348
rect 48265 18302 48457 18307
rect 48512 18270 48582 18488
rect 48637 18451 48829 18456
rect 48637 18410 48648 18451
rect 48638 18348 48648 18410
rect 48637 18307 48648 18348
rect 48818 18410 48829 18451
rect 48818 18348 48828 18410
rect 48818 18307 48829 18348
rect 48637 18302 48829 18307
rect 48884 18270 48954 18488
rect 49009 18451 49201 18456
rect 49009 18410 49020 18451
rect 49010 18348 49020 18410
rect 49009 18307 49020 18348
rect 49190 18410 49201 18451
rect 49190 18348 49200 18410
rect 49190 18307 49201 18348
rect 49009 18302 49201 18307
rect 49256 18270 49326 18488
rect 49381 18451 49573 18456
rect 49381 18410 49392 18451
rect 49382 18348 49392 18410
rect 49381 18307 49392 18348
rect 49562 18410 49573 18451
rect 49562 18348 49572 18410
rect 49562 18307 49573 18348
rect 49381 18302 49573 18307
rect 49604 18270 49678 18488
rect 40720 18258 40815 18270
rect 40720 18082 40775 18258
rect 40809 18082 40815 18258
rect 40720 18070 40815 18082
rect 41027 18258 41187 18270
rect 41027 18082 41033 18258
rect 41067 18082 41147 18258
rect 41181 18082 41187 18258
rect 41027 18070 41187 18082
rect 41399 18258 41559 18270
rect 41399 18082 41405 18258
rect 41439 18082 41519 18258
rect 41553 18082 41559 18258
rect 41399 18070 41559 18082
rect 41771 18258 41931 18270
rect 41771 18082 41777 18258
rect 41811 18082 41891 18258
rect 41925 18082 41931 18258
rect 41771 18070 41931 18082
rect 42143 18258 42303 18270
rect 42143 18082 42149 18258
rect 42183 18082 42263 18258
rect 42297 18082 42303 18258
rect 42143 18070 42303 18082
rect 42515 18258 42675 18270
rect 42515 18082 42521 18258
rect 42555 18082 42635 18258
rect 42669 18082 42675 18258
rect 42515 18070 42675 18082
rect 42887 18258 43047 18270
rect 42887 18082 42893 18258
rect 42927 18082 43007 18258
rect 43041 18082 43047 18258
rect 42887 18070 43047 18082
rect 43259 18258 43419 18270
rect 43259 18082 43265 18258
rect 43299 18082 43379 18258
rect 43413 18082 43419 18258
rect 43259 18070 43419 18082
rect 43631 18258 43791 18270
rect 43631 18082 43637 18258
rect 43671 18082 43751 18258
rect 43785 18082 43791 18258
rect 43631 18070 43791 18082
rect 44003 18258 44163 18270
rect 44003 18082 44009 18258
rect 44043 18082 44123 18258
rect 44157 18082 44163 18258
rect 44003 18070 44163 18082
rect 44375 18258 44535 18270
rect 44375 18082 44381 18258
rect 44415 18082 44495 18258
rect 44529 18082 44535 18258
rect 44375 18070 44535 18082
rect 44747 18258 44907 18270
rect 44747 18082 44753 18258
rect 44787 18082 44867 18258
rect 44901 18082 44907 18258
rect 44747 18070 44907 18082
rect 45119 18258 45279 18270
rect 45119 18082 45125 18258
rect 45159 18082 45239 18258
rect 45273 18082 45279 18258
rect 45119 18070 45279 18082
rect 45491 18258 45651 18270
rect 45491 18082 45497 18258
rect 45531 18082 45611 18258
rect 45645 18082 45651 18258
rect 45491 18070 45651 18082
rect 45863 18258 46023 18270
rect 45863 18082 45869 18258
rect 45903 18082 45983 18258
rect 46017 18082 46023 18258
rect 45863 18070 46023 18082
rect 46235 18258 46395 18270
rect 46235 18082 46241 18258
rect 46275 18082 46355 18258
rect 46389 18082 46395 18258
rect 46235 18070 46395 18082
rect 46607 18258 46767 18270
rect 46607 18082 46613 18258
rect 46647 18082 46727 18258
rect 46761 18082 46767 18258
rect 46607 18070 46767 18082
rect 46979 18258 47139 18270
rect 46979 18082 46985 18258
rect 47019 18082 47099 18258
rect 47133 18082 47139 18258
rect 46979 18070 47139 18082
rect 47351 18258 47511 18270
rect 47351 18082 47357 18258
rect 47391 18082 47471 18258
rect 47505 18082 47511 18258
rect 47351 18070 47511 18082
rect 47723 18258 47883 18270
rect 47723 18082 47729 18258
rect 47763 18082 47843 18258
rect 47877 18082 47883 18258
rect 47723 18070 47883 18082
rect 48095 18258 48255 18270
rect 48095 18082 48101 18258
rect 48135 18082 48215 18258
rect 48249 18082 48255 18258
rect 48095 18070 48255 18082
rect 48467 18258 48627 18270
rect 48467 18082 48473 18258
rect 48507 18082 48587 18258
rect 48621 18082 48627 18258
rect 48467 18070 48627 18082
rect 48839 18258 48999 18270
rect 48839 18082 48845 18258
rect 48879 18082 48959 18258
rect 48993 18082 48999 18258
rect 48839 18070 48999 18082
rect 49211 18258 49371 18270
rect 49211 18082 49217 18258
rect 49251 18082 49331 18258
rect 49365 18082 49371 18258
rect 49211 18070 49371 18082
rect 49583 18258 49678 18270
rect 49583 18082 49589 18258
rect 49623 18082 49678 18258
rect 49583 18070 49678 18082
rect 40720 18069 40794 18070
rect 40826 18038 40836 18043
rect 40825 18033 40836 18038
rect 40824 17987 40836 18033
rect 41006 18038 41016 18043
rect 41006 18033 41017 18038
rect 41072 18033 41142 18070
rect 41444 18069 41514 18070
rect 41198 18038 41208 18043
rect 41197 18033 41208 18038
rect 41006 17987 41208 18033
rect 41378 18038 41388 18043
rect 41570 18038 41580 18043
rect 41378 18033 41389 18038
rect 41378 17987 41390 18033
rect 41569 17992 41580 18038
rect 41750 18038 41760 18043
rect 41570 17987 41580 17992
rect 41750 17992 41761 18038
rect 41750 17987 41760 17992
rect 40824 17977 41390 17987
rect 38304 17108 38314 17616
rect 38800 17108 38810 17616
rect 40826 17380 40836 17383
rect 40825 17334 40836 17380
rect 41006 17380 41016 17383
rect 40826 17329 40836 17334
rect 41006 17334 41017 17380
rect 41006 17329 41016 17334
rect 41072 17293 41142 17977
rect 41816 17849 41886 18070
rect 42188 18069 42258 18070
rect 41942 18038 41952 18043
rect 41941 17992 41952 18038
rect 42122 18038 42132 18043
rect 42314 18038 42324 18043
rect 41942 17987 41952 17992
rect 42122 17992 42133 18038
rect 42313 17992 42324 18038
rect 42494 18038 42504 18043
rect 42122 17987 42132 17992
rect 42314 17987 42324 17992
rect 42494 17992 42505 18038
rect 42494 17987 42504 17992
rect 42560 17849 42630 18070
rect 42932 18069 43002 18070
rect 42686 18038 42696 18043
rect 42685 17992 42696 18038
rect 42866 18038 42876 18043
rect 43058 18038 43068 18043
rect 42686 17987 42696 17992
rect 42866 17992 42877 18038
rect 43057 18033 43068 18038
rect 42866 17987 42876 17992
rect 43056 17987 43068 18033
rect 43238 18038 43248 18043
rect 43238 18033 43249 18038
rect 43304 18033 43374 18070
rect 43676 18069 43746 18070
rect 43430 18038 43440 18043
rect 43429 18033 43440 18038
rect 43238 17987 43440 18033
rect 43610 18038 43620 18043
rect 43802 18038 43812 18043
rect 43610 18033 43621 18038
rect 43610 17987 43622 18033
rect 43801 17992 43812 18038
rect 43982 18038 43992 18043
rect 43802 17987 43812 17992
rect 43982 17992 43993 18038
rect 43982 17987 43992 17992
rect 43056 17977 43622 17987
rect 41806 17669 41816 17849
rect 42630 17669 42640 17849
rect 41198 17380 41208 17383
rect 41197 17334 41208 17380
rect 41378 17380 41388 17383
rect 41570 17380 41580 17383
rect 41198 17329 41208 17334
rect 41378 17334 41389 17380
rect 41569 17334 41580 17380
rect 41750 17380 41760 17383
rect 41378 17329 41388 17334
rect 41570 17329 41580 17334
rect 41750 17334 41761 17380
rect 41750 17329 41760 17334
rect 41816 17293 41886 17669
rect 41942 17380 41952 17383
rect 41941 17334 41952 17380
rect 42122 17380 42132 17383
rect 42314 17380 42324 17383
rect 41942 17329 41952 17334
rect 42122 17334 42133 17380
rect 42313 17334 42324 17380
rect 42494 17380 42504 17383
rect 42122 17329 42132 17334
rect 42314 17329 42324 17334
rect 42494 17334 42505 17380
rect 42494 17329 42504 17334
rect 42560 17293 42630 17669
rect 42686 17380 42696 17383
rect 42685 17334 42696 17380
rect 42866 17380 42876 17383
rect 43058 17380 43068 17383
rect 42686 17329 42696 17334
rect 42866 17334 42877 17380
rect 43057 17334 43068 17380
rect 43238 17380 43248 17383
rect 42866 17329 42876 17334
rect 43058 17329 43068 17334
rect 43238 17334 43249 17380
rect 43238 17329 43248 17334
rect 43304 17293 43374 17977
rect 44048 17525 44118 18070
rect 44420 18069 44490 18070
rect 44174 18038 44184 18043
rect 44173 17992 44184 18038
rect 44354 18038 44364 18043
rect 44546 18038 44556 18043
rect 44174 17987 44184 17992
rect 44354 17992 44365 18038
rect 44545 17992 44556 18038
rect 44726 18038 44736 18043
rect 44354 17987 44364 17992
rect 44546 17987 44556 17992
rect 44726 17992 44737 18038
rect 44726 17987 44736 17992
rect 44792 17525 44862 18070
rect 45164 18069 45234 18070
rect 44918 18038 44928 18043
rect 44917 17992 44928 18038
rect 45098 18038 45108 18043
rect 45290 18038 45300 18043
rect 44918 17987 44928 17992
rect 45098 17992 45109 18038
rect 45289 17992 45300 18038
rect 45470 18038 45480 18043
rect 45098 17987 45108 17992
rect 45290 17987 45300 17992
rect 45470 17992 45481 18038
rect 45470 17987 45480 17992
rect 45536 17525 45606 18070
rect 45908 18069 45978 18070
rect 45662 18038 45672 18043
rect 45661 17992 45672 18038
rect 45842 18038 45852 18043
rect 46034 18038 46044 18043
rect 45662 17987 45672 17992
rect 45842 17992 45853 18038
rect 46033 17992 46044 18038
rect 46214 18038 46224 18043
rect 45842 17987 45852 17992
rect 46034 17987 46044 17992
rect 46214 17992 46225 18038
rect 46214 17987 46224 17992
rect 45816 17541 45826 17815
rect 46104 17541 46114 17815
rect 45912 17529 46026 17541
rect 43430 17380 43440 17383
rect 43429 17334 43440 17380
rect 43610 17380 43620 17383
rect 43430 17329 43440 17334
rect 43610 17334 43621 17380
rect 43610 17329 43620 17334
rect 40722 17281 40815 17293
rect 38390 6698 38728 17108
rect 40722 16505 40775 17281
rect 40809 16505 40815 17281
rect 40722 16493 40815 16505
rect 41027 17281 41187 17293
rect 41027 16505 41033 17281
rect 41067 16505 41147 17281
rect 41181 16505 41187 17281
rect 41027 16493 41187 16505
rect 41399 17281 41559 17293
rect 41399 16505 41405 17281
rect 41439 16505 41519 17281
rect 41553 16505 41559 17281
rect 41399 16493 41559 16505
rect 41771 17281 41931 17293
rect 41771 16505 41777 17281
rect 41811 16505 41891 17281
rect 41925 16505 41931 17281
rect 41771 16493 41931 16505
rect 42143 17281 42303 17293
rect 42143 16505 42149 17281
rect 42183 16505 42263 17281
rect 42297 16505 42303 17281
rect 42143 16493 42303 16505
rect 42515 17281 42675 17293
rect 42515 16505 42521 17281
rect 42555 16505 42635 17281
rect 42669 16505 42675 17281
rect 42515 16493 42675 16505
rect 42887 17281 43047 17293
rect 42887 16505 42893 17281
rect 42927 16505 43007 17281
rect 43041 16505 43047 17281
rect 42887 16493 43047 16505
rect 43259 17281 43419 17293
rect 43259 16505 43265 17281
rect 43299 16505 43379 17281
rect 43413 16505 43419 17281
rect 43259 16493 43419 16505
rect 43631 17281 43724 17293
rect 43631 16505 43637 17281
rect 43671 16505 43724 17281
rect 43932 17253 43942 17525
rect 44224 17253 44234 17525
rect 44676 17253 44686 17525
rect 44968 17253 44978 17525
rect 45420 17253 45430 17525
rect 45712 17253 45722 17525
rect 45952 17481 46026 17529
rect 46280 17525 46350 18070
rect 46652 18069 46722 18070
rect 46406 18038 46416 18043
rect 46405 17992 46416 18038
rect 46586 18038 46596 18043
rect 46778 18038 46788 18043
rect 46406 17987 46416 17992
rect 46586 17992 46597 18038
rect 46777 17992 46788 18038
rect 46958 18038 46968 18043
rect 46586 17987 46596 17992
rect 46778 17987 46788 17992
rect 46958 17992 46969 18038
rect 46958 17987 46968 17992
rect 47024 17525 47094 18070
rect 47396 18069 47466 18070
rect 47150 18038 47160 18043
rect 47149 17992 47160 18038
rect 47330 18038 47340 18043
rect 47522 18038 47532 18043
rect 47150 17987 47160 17992
rect 47330 17992 47341 18038
rect 47521 17992 47532 18038
rect 47702 18038 47712 18043
rect 47330 17987 47340 17992
rect 47522 17987 47532 17992
rect 47702 17992 47713 18038
rect 47702 17987 47712 17992
rect 47768 17525 47838 18070
rect 48140 18069 48210 18070
rect 47894 18038 47904 18043
rect 47893 17992 47904 18038
rect 48074 18038 48084 18043
rect 48266 18038 48276 18043
rect 47894 17987 47904 17992
rect 48074 17992 48085 18038
rect 48265 17992 48276 18038
rect 48446 18038 48456 18043
rect 48074 17987 48084 17992
rect 48266 17987 48276 17992
rect 48446 17992 48457 18038
rect 48446 17987 48456 17992
rect 48512 17525 48582 18070
rect 48884 18069 48954 18070
rect 48638 18038 48648 18043
rect 48637 17992 48648 18038
rect 48818 18038 48828 18043
rect 49010 18038 49020 18043
rect 48638 17987 48648 17992
rect 48818 17992 48829 18038
rect 49009 17992 49020 18038
rect 49190 18038 49200 18043
rect 48818 17987 48828 17992
rect 49010 17987 49020 17992
rect 49190 17992 49201 18038
rect 49190 17987 49200 17992
rect 49256 17525 49326 18070
rect 49604 18057 49678 18070
rect 49382 18038 49392 18043
rect 49381 17992 49392 18038
rect 49562 18038 49572 18043
rect 49382 17987 49392 17992
rect 49562 17992 49573 18038
rect 49562 17987 49572 17992
rect 43631 16493 43724 16505
rect 40722 16257 40770 16493
rect 40825 16447 41017 16452
rect 40825 16406 40836 16447
rect 40826 16344 40836 16406
rect 40825 16303 40836 16344
rect 41006 16406 41017 16447
rect 41006 16344 41016 16406
rect 41006 16303 41017 16344
rect 40825 16298 41017 16303
rect 41072 16257 41142 16493
rect 41197 16447 41389 16452
rect 41197 16406 41208 16447
rect 41198 16344 41208 16406
rect 41197 16303 41208 16344
rect 41378 16406 41389 16447
rect 41378 16344 41388 16406
rect 41378 16303 41389 16344
rect 41197 16298 41389 16303
rect 41444 16257 41514 16493
rect 41569 16447 41761 16452
rect 41569 16406 41580 16447
rect 41570 16344 41580 16406
rect 41569 16303 41580 16344
rect 41750 16406 41761 16447
rect 41750 16344 41760 16406
rect 41750 16303 41761 16344
rect 41569 16298 41761 16303
rect 41816 16257 41886 16493
rect 41941 16447 42133 16452
rect 41941 16406 41952 16447
rect 41942 16344 41952 16406
rect 41941 16303 41952 16344
rect 42122 16406 42133 16447
rect 42122 16344 42132 16406
rect 42122 16303 42133 16344
rect 41941 16298 42133 16303
rect 42188 16257 42258 16493
rect 42313 16447 42505 16452
rect 42313 16406 42324 16447
rect 42314 16344 42324 16406
rect 42313 16303 42324 16344
rect 42494 16406 42505 16447
rect 42494 16344 42504 16406
rect 42494 16303 42505 16344
rect 42313 16298 42505 16303
rect 42560 16257 42630 16493
rect 42685 16447 42877 16452
rect 42685 16406 42696 16447
rect 42686 16344 42696 16406
rect 42685 16303 42696 16344
rect 42866 16406 42877 16447
rect 42866 16344 42876 16406
rect 42866 16303 42877 16344
rect 42685 16298 42877 16303
rect 42932 16257 43002 16493
rect 43057 16447 43249 16452
rect 43057 16406 43068 16447
rect 43058 16344 43068 16406
rect 43057 16303 43068 16344
rect 43238 16406 43249 16447
rect 43238 16344 43248 16406
rect 43238 16303 43249 16344
rect 43057 16298 43249 16303
rect 43304 16257 43374 16493
rect 43429 16447 43621 16452
rect 43429 16406 43440 16447
rect 43430 16344 43440 16406
rect 43429 16303 43440 16344
rect 43610 16406 43621 16447
rect 43610 16344 43620 16406
rect 43610 16303 43621 16344
rect 43429 16298 43621 16303
rect 43670 16257 43724 16493
rect 45556 16304 45566 16470
rect 45734 16420 45744 16470
rect 45954 16434 46026 17481
rect 46164 17253 46174 17525
rect 46456 17253 46466 17525
rect 46908 17253 46918 17525
rect 47200 17253 47210 17525
rect 47652 17253 47662 17525
rect 47944 17253 47954 17525
rect 48396 17253 48406 17525
rect 48688 17253 48698 17525
rect 49140 17253 49150 17525
rect 49432 17253 49442 17525
rect 45734 16419 45864 16420
rect 45734 16413 45879 16419
rect 45734 16365 45813 16413
rect 45867 16365 45879 16413
rect 45734 16359 45879 16365
rect 45734 16358 45864 16359
rect 45734 16304 45744 16358
rect 40722 16245 40815 16257
rect 40722 15469 40775 16245
rect 40809 15469 40815 16245
rect 40722 15457 40815 15469
rect 41027 16245 41187 16257
rect 41027 15469 41033 16245
rect 41067 15469 41147 16245
rect 41181 15469 41187 16245
rect 41027 15457 41187 15469
rect 41399 16245 41559 16257
rect 41399 15469 41405 16245
rect 41439 15469 41519 16245
rect 41553 15469 41559 16245
rect 41399 15457 41559 15469
rect 41771 16245 41931 16257
rect 41771 15469 41777 16245
rect 41811 15469 41891 16245
rect 41925 15469 41931 16245
rect 41771 15457 41931 15469
rect 42143 16245 42303 16257
rect 42143 15469 42149 16245
rect 42183 15469 42263 16245
rect 42297 15469 42303 16245
rect 42143 15457 42303 15469
rect 42515 16245 42675 16257
rect 42515 15469 42521 16245
rect 42555 15469 42635 16245
rect 42669 15469 42675 16245
rect 42515 15457 42675 15469
rect 42887 16245 43047 16257
rect 42887 15469 42893 16245
rect 42927 15469 43007 16245
rect 43041 15469 43047 16245
rect 42887 15457 43047 15469
rect 43259 16245 43419 16257
rect 43259 15469 43265 16245
rect 43299 15469 43379 16245
rect 43413 15469 43419 16245
rect 43259 15457 43419 15469
rect 43631 16245 43724 16257
rect 43631 15469 43637 16245
rect 43671 15469 43724 16245
rect 45556 15904 45566 16070
rect 45734 16020 45744 16070
rect 45954 16037 45971 16434
rect 46009 16037 46026 16434
rect 45734 16019 45864 16020
rect 45954 16019 46026 16037
rect 45734 16013 45879 16019
rect 45734 15965 45813 16013
rect 45867 15965 45879 16013
rect 45734 15959 45879 15965
rect 45734 15958 45864 15959
rect 45734 15904 45744 15958
rect 45954 15903 46026 15921
rect 45556 15504 45566 15670
rect 45734 15620 45744 15670
rect 45734 15619 45864 15620
rect 45734 15613 45879 15619
rect 45734 15565 45813 15613
rect 45867 15565 45879 15613
rect 45734 15559 45879 15565
rect 45734 15558 45864 15559
rect 45734 15504 45744 15558
rect 45954 15506 45971 15903
rect 46009 15506 46026 15903
rect 43631 15457 43724 15469
rect 40722 15221 40770 15457
rect 40825 15411 41017 15416
rect 40825 15370 40836 15411
rect 40826 15308 40836 15370
rect 40825 15267 40836 15308
rect 41006 15370 41017 15411
rect 41006 15308 41016 15370
rect 41006 15267 41017 15308
rect 40825 15262 41017 15267
rect 41072 15221 41142 15457
rect 41197 15411 41389 15416
rect 41197 15370 41208 15411
rect 41198 15308 41208 15370
rect 41197 15267 41208 15308
rect 41378 15370 41389 15411
rect 41378 15308 41388 15370
rect 41378 15267 41389 15308
rect 41197 15262 41389 15267
rect 41444 15221 41514 15457
rect 41569 15411 41761 15416
rect 41569 15370 41580 15411
rect 41570 15308 41580 15370
rect 41569 15267 41580 15308
rect 41750 15370 41761 15411
rect 41750 15308 41760 15370
rect 41750 15267 41761 15308
rect 41569 15262 41761 15267
rect 41816 15221 41886 15457
rect 41941 15411 42133 15416
rect 41941 15370 41952 15411
rect 41942 15308 41952 15370
rect 41941 15267 41952 15308
rect 42122 15370 42133 15411
rect 42122 15308 42132 15370
rect 42122 15267 42133 15308
rect 41941 15262 42133 15267
rect 42188 15221 42258 15457
rect 42313 15411 42505 15416
rect 42313 15370 42324 15411
rect 42314 15308 42324 15370
rect 42313 15267 42324 15308
rect 42494 15370 42505 15411
rect 42494 15308 42504 15370
rect 42494 15267 42505 15308
rect 42313 15262 42505 15267
rect 42560 15221 42630 15457
rect 42685 15411 42877 15416
rect 42685 15370 42696 15411
rect 42686 15308 42696 15370
rect 42685 15267 42696 15308
rect 42866 15370 42877 15411
rect 42866 15308 42876 15370
rect 42866 15267 42877 15308
rect 42685 15262 42877 15267
rect 42932 15221 43002 15457
rect 43057 15411 43249 15416
rect 43057 15370 43068 15411
rect 43058 15308 43068 15370
rect 43057 15267 43068 15308
rect 43238 15370 43249 15411
rect 43238 15308 43248 15370
rect 43238 15267 43249 15308
rect 43057 15262 43249 15267
rect 43304 15221 43374 15457
rect 43429 15411 43621 15416
rect 43429 15370 43440 15411
rect 43430 15308 43440 15370
rect 43429 15267 43440 15308
rect 43610 15370 43621 15411
rect 43610 15308 43620 15370
rect 43610 15267 43621 15308
rect 43429 15262 43621 15267
rect 43670 15221 43724 15457
rect 40722 15209 40815 15221
rect 40722 14433 40775 15209
rect 40809 14433 40815 15209
rect 40722 14421 40815 14433
rect 41027 15209 41187 15221
rect 41027 14433 41033 15209
rect 41067 14433 41147 15209
rect 41181 14433 41187 15209
rect 41027 14421 41187 14433
rect 41399 15209 41559 15221
rect 41399 14433 41405 15209
rect 41439 14433 41519 15209
rect 41553 14433 41559 15209
rect 41399 14421 41559 14433
rect 41771 15209 41931 15221
rect 41771 14433 41777 15209
rect 41811 14433 41891 15209
rect 41925 14433 41931 15209
rect 41771 14421 41931 14433
rect 42143 15209 42303 15221
rect 42143 14433 42149 15209
rect 42183 14433 42263 15209
rect 42297 14433 42303 15209
rect 42143 14421 42303 14433
rect 42515 15209 42675 15221
rect 42515 14433 42521 15209
rect 42555 14433 42635 15209
rect 42669 14433 42675 15209
rect 42515 14421 42675 14433
rect 42887 15209 43047 15221
rect 42887 14433 42893 15209
rect 42927 14433 43007 15209
rect 43041 14433 43047 15209
rect 42887 14421 43047 14433
rect 43259 15209 43419 15221
rect 43259 14433 43265 15209
rect 43299 14433 43379 15209
rect 43413 14433 43419 15209
rect 43259 14421 43419 14433
rect 43631 15209 43724 15221
rect 43631 14433 43637 15209
rect 43671 14433 43724 15209
rect 45954 15117 46026 15506
rect 45842 14845 45852 15117
rect 46134 14845 46144 15117
rect 43631 14421 43724 14433
rect 40722 14185 40770 14421
rect 40825 14375 41017 14380
rect 40825 14334 40836 14375
rect 40826 14272 40836 14334
rect 40825 14231 40836 14272
rect 41006 14334 41017 14375
rect 41006 14272 41016 14334
rect 41006 14231 41017 14272
rect 40825 14226 41017 14231
rect 41072 14185 41142 14421
rect 41197 14375 41389 14380
rect 41197 14334 41208 14375
rect 41198 14272 41208 14334
rect 41197 14231 41208 14272
rect 41378 14334 41389 14375
rect 41378 14272 41388 14334
rect 41378 14231 41389 14272
rect 41197 14226 41389 14231
rect 41444 14185 41514 14421
rect 41569 14375 41761 14380
rect 41569 14334 41580 14375
rect 41570 14272 41580 14334
rect 41569 14231 41580 14272
rect 41750 14334 41761 14375
rect 41750 14272 41760 14334
rect 41750 14231 41761 14272
rect 41569 14226 41761 14231
rect 41816 14185 41886 14421
rect 41941 14375 42133 14380
rect 41941 14334 41952 14375
rect 41942 14272 41952 14334
rect 41941 14231 41952 14272
rect 42122 14334 42133 14375
rect 42122 14272 42132 14334
rect 42122 14231 42133 14272
rect 41941 14226 42133 14231
rect 42188 14185 42258 14421
rect 42313 14375 42505 14380
rect 42313 14334 42324 14375
rect 42314 14272 42324 14334
rect 42313 14231 42324 14272
rect 42494 14334 42505 14375
rect 42494 14272 42504 14334
rect 42494 14231 42505 14272
rect 42313 14226 42505 14231
rect 42560 14185 42630 14421
rect 42685 14375 42877 14380
rect 42685 14334 42696 14375
rect 42686 14272 42696 14334
rect 42685 14231 42696 14272
rect 42866 14334 42877 14375
rect 42866 14272 42876 14334
rect 42866 14231 42877 14272
rect 42685 14226 42877 14231
rect 42932 14185 43002 14421
rect 43057 14375 43249 14380
rect 43057 14334 43068 14375
rect 43058 14272 43068 14334
rect 43057 14231 43068 14272
rect 43238 14334 43249 14375
rect 43238 14272 43248 14334
rect 43238 14231 43249 14272
rect 43057 14226 43249 14231
rect 43304 14185 43374 14421
rect 43429 14375 43621 14380
rect 43429 14334 43440 14375
rect 43430 14272 43440 14334
rect 43429 14231 43440 14272
rect 43610 14334 43621 14375
rect 43610 14272 43620 14334
rect 43610 14231 43621 14272
rect 43429 14226 43621 14231
rect 43670 14185 43724 14421
rect 40722 14173 40815 14185
rect 40722 13397 40775 14173
rect 40809 13397 40815 14173
rect 40722 13385 40815 13397
rect 41027 14173 41187 14185
rect 41027 13397 41033 14173
rect 41067 13397 41147 14173
rect 41181 13397 41187 14173
rect 41027 13385 41187 13397
rect 41399 14173 41559 14185
rect 41399 13397 41405 14173
rect 41439 13397 41519 14173
rect 41553 13397 41559 14173
rect 41399 13385 41559 13397
rect 41771 14173 41931 14185
rect 41771 13397 41777 14173
rect 41811 13397 41891 14173
rect 41925 13397 41931 14173
rect 41771 13385 41931 13397
rect 42143 14173 42303 14185
rect 42143 13397 42149 14173
rect 42183 13397 42263 14173
rect 42297 13397 42303 14173
rect 42143 13385 42303 13397
rect 42515 14173 42675 14185
rect 42515 13397 42521 14173
rect 42555 13397 42635 14173
rect 42669 13397 42675 14173
rect 42515 13385 42675 13397
rect 42887 14173 43047 14185
rect 42887 13397 42893 14173
rect 42927 13397 43007 14173
rect 43041 13397 43047 14173
rect 42887 13385 43047 13397
rect 43259 14173 43419 14185
rect 43259 13397 43265 14173
rect 43299 13397 43379 14173
rect 43413 13397 43419 14173
rect 43259 13385 43419 13397
rect 43631 14173 43724 14185
rect 43631 13397 43637 14173
rect 43671 13397 43724 14173
rect 43631 13385 43724 13397
rect 40722 13261 40776 13385
rect 40826 13344 40836 13353
rect 40825 13298 40836 13344
rect 41006 13344 41016 13353
rect 41198 13344 41208 13353
rect 40826 13289 40836 13298
rect 41006 13298 41017 13344
rect 41197 13298 41208 13344
rect 41378 13344 41388 13353
rect 41006 13289 41016 13298
rect 41198 13289 41208 13298
rect 41378 13298 41389 13344
rect 41378 13289 41388 13298
rect 41450 13261 41508 13385
rect 41570 13344 41580 13353
rect 41569 13298 41580 13344
rect 41750 13344 41760 13353
rect 41942 13344 41952 13353
rect 41570 13289 41580 13298
rect 41750 13298 41761 13344
rect 41941 13298 41952 13344
rect 42122 13344 42132 13353
rect 41750 13289 41760 13298
rect 41942 13289 41952 13298
rect 42122 13298 42133 13344
rect 42122 13289 42132 13298
rect 42194 13261 42252 13385
rect 42314 13344 42324 13353
rect 42313 13298 42324 13344
rect 42494 13344 42504 13353
rect 42686 13344 42696 13353
rect 42314 13289 42324 13298
rect 42494 13298 42505 13344
rect 42685 13298 42696 13344
rect 42866 13344 42876 13353
rect 42494 13289 42504 13298
rect 42686 13289 42696 13298
rect 42866 13298 42877 13344
rect 42866 13289 42876 13298
rect 42938 13261 42996 13385
rect 43058 13344 43068 13353
rect 43057 13298 43068 13344
rect 43238 13344 43248 13353
rect 43430 13344 43440 13353
rect 43058 13289 43068 13298
rect 43238 13298 43249 13344
rect 43429 13298 43440 13344
rect 43610 13344 43620 13353
rect 43238 13289 43248 13298
rect 43430 13289 43440 13298
rect 43610 13298 43621 13344
rect 43610 13289 43620 13298
rect 43670 13261 43724 13385
rect 40722 13255 40828 13261
rect 40722 13185 40746 13255
rect 40816 13185 40828 13255
rect 40722 13179 40828 13185
rect 41106 13255 41200 13261
rect 41106 13185 41118 13255
rect 41188 13185 41200 13255
rect 41106 13179 41200 13185
rect 41450 13255 41572 13261
rect 41450 13185 41490 13255
rect 41560 13185 41572 13255
rect 41450 13179 41572 13185
rect 41850 13255 41944 13261
rect 41850 13185 41862 13255
rect 41932 13185 41944 13255
rect 41850 13179 41944 13185
rect 42194 13255 42316 13261
rect 42194 13185 42234 13255
rect 42304 13185 42316 13255
rect 42194 13179 42316 13185
rect 42594 13255 42688 13261
rect 42594 13185 42606 13255
rect 42676 13185 42688 13255
rect 42594 13179 42688 13185
rect 42938 13255 43060 13261
rect 42938 13185 42978 13255
rect 43048 13185 43060 13255
rect 42938 13179 43060 13185
rect 43338 13255 43432 13261
rect 43338 13185 43350 13255
rect 43420 13185 43432 13255
rect 43338 13179 43432 13185
rect 43600 13255 43724 13261
rect 43600 13185 43612 13255
rect 43682 13185 43724 13255
rect 43600 13179 43724 13185
rect 40722 13075 40776 13179
rect 41118 13075 41188 13179
rect 41450 13075 41508 13179
rect 41862 13075 41932 13179
rect 42194 13075 42252 13179
rect 42606 13075 42676 13179
rect 42938 13075 42996 13179
rect 43350 13075 43420 13179
rect 43670 13075 43724 13179
rect 39962 13011 44484 13075
rect 45422 13071 45432 13343
rect 45714 13071 45724 13343
rect 46166 13071 46176 13343
rect 46458 13071 46468 13343
rect 46910 13071 46920 13343
rect 47202 13071 47212 13343
rect 47654 13071 47664 13343
rect 47946 13071 47956 13343
rect 48398 13071 48408 13343
rect 48690 13071 48700 13343
rect 49142 13071 49152 13343
rect 49434 13071 49444 13343
rect 49886 13071 49896 13343
rect 50178 13071 50188 13343
rect 50630 13071 50640 13343
rect 50922 13071 50932 13343
rect 39280 12703 39348 12763
rect 39518 12756 39528 12763
rect 39710 12756 39720 12763
rect 39518 12710 39529 12756
rect 39709 12710 39720 12756
rect 39890 12756 39900 12763
rect 39518 12703 39528 12710
rect 39710 12703 39720 12710
rect 39890 12710 39901 12756
rect 39890 12703 39900 12710
rect 39280 12657 39328 12703
rect 39962 12669 40020 13011
rect 40580 12763 40910 12765
rect 40082 12756 40092 12763
rect 40081 12710 40092 12756
rect 40262 12756 40272 12763
rect 40454 12756 40464 12763
rect 40082 12703 40092 12710
rect 40262 12710 40273 12756
rect 40453 12710 40464 12756
rect 40262 12703 40272 12710
rect 40454 12703 40464 12710
rect 40634 12703 40836 12763
rect 41006 12756 41016 12763
rect 41198 12756 41208 12763
rect 41006 12710 41017 12756
rect 41197 12710 41208 12756
rect 41378 12756 41388 12763
rect 41006 12703 41016 12710
rect 41198 12703 41208 12710
rect 41378 12710 41389 12756
rect 41378 12703 41388 12710
rect 40706 12669 40764 12703
rect 41450 12669 41508 13011
rect 41570 12756 41580 12763
rect 41569 12710 41580 12756
rect 41750 12756 41760 12763
rect 41942 12756 41952 12763
rect 41570 12703 41580 12710
rect 41750 12710 41761 12756
rect 41941 12710 41952 12756
rect 41750 12703 41760 12710
rect 41942 12703 41952 12710
rect 42122 12703 42324 12763
rect 42494 12756 42504 12763
rect 42686 12756 42696 12763
rect 42494 12710 42505 12756
rect 42685 12710 42696 12756
rect 42866 12756 42876 12763
rect 42494 12703 42504 12710
rect 42686 12703 42696 12710
rect 42866 12710 42877 12756
rect 42866 12703 42876 12710
rect 42194 12669 42252 12703
rect 42938 12669 42996 13011
rect 43058 12756 43068 12763
rect 43057 12710 43068 12756
rect 43238 12756 43248 12763
rect 43430 12756 43440 12763
rect 43058 12703 43068 12710
rect 43238 12710 43249 12756
rect 43429 12710 43440 12756
rect 43238 12703 43248 12710
rect 43430 12703 43440 12710
rect 43610 12703 43812 12763
rect 43982 12756 43992 12763
rect 44174 12756 44184 12763
rect 43982 12710 43993 12756
rect 44173 12710 44184 12756
rect 44354 12756 44364 12763
rect 43982 12703 43992 12710
rect 44174 12703 44184 12710
rect 44354 12710 44365 12756
rect 44354 12703 44364 12710
rect 43682 12669 43740 12703
rect 44426 12669 44484 13011
rect 44546 12756 44556 12763
rect 44545 12710 44556 12756
rect 44726 12756 44736 12763
rect 44918 12756 44928 12763
rect 44546 12703 44556 12710
rect 44726 12710 44737 12756
rect 44917 12710 44928 12756
rect 44726 12703 44736 12710
rect 44918 12703 44928 12710
rect 45098 12703 45170 12763
rect 45286 12703 45300 12763
rect 45470 12756 45480 12763
rect 45470 12710 45481 12756
rect 45470 12703 45480 12710
rect 39280 12281 39287 12657
rect 39321 12281 39328 12657
rect 39280 12233 39328 12281
rect 39539 12657 39699 12669
rect 39539 12281 39545 12657
rect 39579 12281 39659 12657
rect 39693 12281 39699 12657
rect 39539 12269 39699 12281
rect 39911 12657 40071 12669
rect 39911 12281 39917 12657
rect 39951 12281 40031 12657
rect 40065 12281 40071 12657
rect 39911 12269 40071 12281
rect 40283 12657 40443 12669
rect 40283 12281 40289 12657
rect 40323 12281 40403 12657
rect 40437 12281 40443 12657
rect 40283 12269 40443 12281
rect 40655 12657 40815 12669
rect 40655 12281 40661 12657
rect 40695 12281 40775 12657
rect 40809 12281 40815 12657
rect 40655 12269 40815 12281
rect 41027 12657 41187 12669
rect 41027 12281 41033 12657
rect 41067 12281 41147 12657
rect 41181 12281 41187 12657
rect 41027 12269 41187 12281
rect 41399 12657 41559 12669
rect 41399 12281 41405 12657
rect 41439 12281 41519 12657
rect 41553 12281 41559 12657
rect 41399 12269 41559 12281
rect 41771 12657 41931 12669
rect 41771 12281 41777 12657
rect 41811 12281 41891 12657
rect 41925 12281 41931 12657
rect 41771 12269 41931 12281
rect 42143 12657 42303 12669
rect 42143 12281 42149 12657
rect 42183 12281 42263 12657
rect 42297 12281 42303 12657
rect 42143 12269 42303 12281
rect 42515 12657 42675 12669
rect 42515 12281 42521 12657
rect 42555 12281 42635 12657
rect 42669 12281 42675 12657
rect 42515 12269 42675 12281
rect 42887 12657 43047 12669
rect 42887 12281 42893 12657
rect 42927 12281 43007 12657
rect 43041 12281 43047 12657
rect 42887 12269 43047 12281
rect 43259 12657 43419 12669
rect 43259 12281 43265 12657
rect 43299 12281 43379 12657
rect 43413 12281 43419 12657
rect 43259 12269 43419 12281
rect 43631 12657 43791 12669
rect 43631 12281 43637 12657
rect 43671 12281 43751 12657
rect 43785 12281 43791 12657
rect 43631 12269 43791 12281
rect 44003 12657 44163 12669
rect 44003 12281 44009 12657
rect 44043 12281 44123 12657
rect 44157 12281 44163 12657
rect 44003 12269 44163 12281
rect 44375 12657 44535 12669
rect 44375 12281 44381 12657
rect 44415 12281 44495 12657
rect 44529 12281 44535 12657
rect 44375 12269 44535 12281
rect 44747 12657 44907 12669
rect 44747 12281 44753 12657
rect 44787 12281 44867 12657
rect 44901 12281 44907 12657
rect 44747 12269 44907 12281
rect 45118 12657 45170 12703
rect 45536 12669 45606 13071
rect 45662 12756 45672 12763
rect 45661 12710 45672 12756
rect 45842 12756 45852 12763
rect 46034 12756 46044 12763
rect 45662 12703 45672 12710
rect 45842 12710 45853 12756
rect 46033 12710 46044 12756
rect 46214 12756 46224 12763
rect 45842 12703 45852 12710
rect 46034 12703 46044 12710
rect 46214 12710 46225 12756
rect 46214 12703 46224 12710
rect 46280 12669 46350 13071
rect 46406 12756 46416 12763
rect 46405 12710 46416 12756
rect 46586 12756 46596 12763
rect 46778 12756 46788 12763
rect 46406 12703 46416 12710
rect 46586 12710 46597 12756
rect 46777 12710 46788 12756
rect 46958 12756 46968 12763
rect 46586 12703 46596 12710
rect 46778 12703 46788 12710
rect 46958 12710 46969 12756
rect 46958 12703 46968 12710
rect 47024 12669 47094 13071
rect 47150 12756 47160 12763
rect 47149 12710 47160 12756
rect 47330 12756 47340 12763
rect 47522 12756 47532 12763
rect 47150 12703 47160 12710
rect 47330 12710 47341 12756
rect 47521 12710 47532 12756
rect 47702 12756 47712 12763
rect 47330 12703 47340 12710
rect 47522 12703 47532 12710
rect 47702 12710 47713 12756
rect 47702 12703 47712 12710
rect 47768 12669 47838 13071
rect 47894 12756 47904 12763
rect 47893 12710 47904 12756
rect 48074 12756 48084 12763
rect 48266 12756 48276 12763
rect 47894 12703 47904 12710
rect 48074 12710 48085 12756
rect 48265 12710 48276 12756
rect 48446 12756 48456 12763
rect 48074 12703 48084 12710
rect 48266 12703 48276 12710
rect 48446 12710 48457 12756
rect 48446 12703 48456 12710
rect 48512 12669 48582 13071
rect 48638 12756 48648 12763
rect 48637 12710 48648 12756
rect 48818 12756 48828 12763
rect 49010 12756 49020 12763
rect 48638 12703 48648 12710
rect 48818 12710 48829 12756
rect 49009 12710 49020 12756
rect 49190 12756 49200 12763
rect 48818 12703 48828 12710
rect 49010 12703 49020 12710
rect 49190 12710 49201 12756
rect 49190 12703 49200 12710
rect 49256 12669 49326 13071
rect 49382 12756 49392 12763
rect 49381 12710 49392 12756
rect 49562 12756 49572 12763
rect 49754 12756 49764 12763
rect 49382 12703 49392 12710
rect 49562 12710 49573 12756
rect 49753 12710 49764 12756
rect 49934 12756 49944 12763
rect 49562 12703 49572 12710
rect 49754 12703 49764 12710
rect 49934 12710 49945 12756
rect 49934 12703 49944 12710
rect 50000 12669 50070 13071
rect 50126 12756 50136 12763
rect 50125 12710 50136 12756
rect 50306 12756 50316 12763
rect 50498 12756 50508 12763
rect 50126 12703 50136 12710
rect 50306 12710 50317 12756
rect 50497 12710 50508 12756
rect 50678 12756 50688 12763
rect 50306 12703 50316 12710
rect 50498 12703 50508 12710
rect 50678 12710 50689 12756
rect 50678 12703 50688 12710
rect 50744 12669 50814 13071
rect 50870 12756 50880 12763
rect 50869 12710 50880 12756
rect 51050 12756 51060 12763
rect 50870 12703 50880 12710
rect 51050 12710 51061 12756
rect 51050 12703 51060 12710
rect 45118 12281 45125 12657
rect 45159 12281 45170 12657
rect 39280 12228 39370 12233
rect 39280 12223 39529 12228
rect 39280 12079 39348 12223
rect 39518 12182 39529 12223
rect 39518 12120 39528 12182
rect 39518 12079 39529 12120
rect 39280 12074 39529 12079
rect 39280 12073 39370 12074
rect 39280 12021 39328 12073
rect 39584 12033 39654 12269
rect 39709 12223 39901 12228
rect 39709 12182 39720 12223
rect 39710 12120 39720 12182
rect 39709 12079 39720 12120
rect 39890 12182 39901 12223
rect 39890 12120 39900 12182
rect 39890 12079 39901 12120
rect 39709 12074 39901 12079
rect 39956 12033 40026 12269
rect 40081 12223 40273 12228
rect 40081 12182 40092 12223
rect 40082 12120 40092 12182
rect 40081 12079 40092 12120
rect 40262 12182 40273 12223
rect 40262 12120 40272 12182
rect 40262 12079 40273 12120
rect 40081 12074 40273 12079
rect 40328 12033 40398 12269
rect 40700 12229 40770 12269
rect 40494 12228 40970 12229
rect 40453 12223 41017 12228
rect 40453 12182 40464 12223
rect 40454 12120 40464 12182
rect 40453 12079 40464 12120
rect 40634 12079 40836 12223
rect 41006 12182 41017 12223
rect 41006 12120 41016 12182
rect 41006 12079 41017 12120
rect 40453 12077 41017 12079
rect 40453 12074 40645 12077
rect 40700 12033 40770 12077
rect 40825 12074 41017 12077
rect 41072 12033 41142 12269
rect 41197 12223 41389 12228
rect 41197 12182 41208 12223
rect 41198 12120 41208 12182
rect 41197 12079 41208 12120
rect 41378 12182 41389 12223
rect 41378 12120 41388 12182
rect 41378 12079 41389 12120
rect 41197 12074 41389 12079
rect 41444 12033 41514 12269
rect 41569 12223 41761 12228
rect 41569 12182 41580 12223
rect 41570 12120 41580 12182
rect 41569 12079 41580 12120
rect 41750 12182 41761 12223
rect 41750 12120 41760 12182
rect 41750 12079 41761 12120
rect 41569 12074 41761 12079
rect 41816 12033 41886 12269
rect 42188 12229 42258 12269
rect 42016 12228 42434 12229
rect 41941 12223 42505 12228
rect 41941 12182 41952 12223
rect 41942 12120 41952 12182
rect 41941 12079 41952 12120
rect 42122 12079 42324 12223
rect 42494 12182 42505 12223
rect 42494 12120 42504 12182
rect 42494 12079 42505 12120
rect 41941 12074 42505 12079
rect 42016 12073 42434 12074
rect 42188 12033 42258 12073
rect 42560 12033 42630 12269
rect 42685 12223 42877 12228
rect 42685 12182 42696 12223
rect 42686 12120 42696 12182
rect 42685 12079 42696 12120
rect 42866 12182 42877 12223
rect 42866 12120 42876 12182
rect 42866 12079 42877 12120
rect 42685 12074 42877 12079
rect 42932 12033 43002 12269
rect 43057 12223 43249 12228
rect 43057 12182 43068 12223
rect 43058 12120 43068 12182
rect 43057 12079 43068 12120
rect 43238 12182 43249 12223
rect 43238 12120 43248 12182
rect 43238 12079 43249 12120
rect 43057 12074 43249 12079
rect 43304 12033 43374 12269
rect 43676 12229 43746 12269
rect 43512 12228 43888 12229
rect 43429 12223 43993 12228
rect 43429 12182 43440 12223
rect 43430 12120 43440 12182
rect 43429 12079 43440 12120
rect 43610 12079 43812 12223
rect 43982 12182 43993 12223
rect 43982 12120 43992 12182
rect 43982 12079 43993 12120
rect 43429 12074 43993 12079
rect 43512 12073 43888 12074
rect 43676 12033 43746 12073
rect 44048 12033 44118 12269
rect 44173 12223 44365 12228
rect 44173 12182 44184 12223
rect 44174 12120 44184 12182
rect 44173 12079 44184 12120
rect 44354 12182 44365 12223
rect 44354 12120 44364 12182
rect 44354 12079 44365 12120
rect 44173 12074 44365 12079
rect 44420 12033 44490 12269
rect 44545 12223 44737 12228
rect 44545 12182 44556 12223
rect 44546 12120 44556 12182
rect 44545 12079 44556 12120
rect 44726 12182 44737 12223
rect 44726 12120 44736 12182
rect 44726 12079 44737 12120
rect 44545 12074 44737 12079
rect 44792 12033 44862 12269
rect 45118 12229 45170 12281
rect 45028 12228 45170 12229
rect 44917 12223 45170 12228
rect 44917 12182 44928 12223
rect 44918 12120 44928 12182
rect 44917 12079 44928 12120
rect 45098 12079 45170 12223
rect 44917 12074 45170 12079
rect 45028 12073 45170 12074
rect 39280 11645 39287 12021
rect 39321 11645 39328 12021
rect 39280 11593 39328 11645
rect 39539 12021 39699 12033
rect 39539 11645 39545 12021
rect 39579 11645 39659 12021
rect 39693 11645 39699 12021
rect 39539 11633 39699 11645
rect 39911 12021 40071 12033
rect 39911 11645 39917 12021
rect 39951 11645 40031 12021
rect 40065 11645 40071 12021
rect 39911 11633 40071 11645
rect 40283 12021 40443 12033
rect 40283 11645 40289 12021
rect 40323 11645 40403 12021
rect 40437 11645 40443 12021
rect 40283 11633 40443 11645
rect 40655 12021 40815 12033
rect 40655 11645 40661 12021
rect 40695 11645 40775 12021
rect 40809 11645 40815 12021
rect 40655 11633 40815 11645
rect 41027 12021 41187 12033
rect 41027 11645 41033 12021
rect 41067 11645 41147 12021
rect 41181 11645 41187 12021
rect 41027 11633 41187 11645
rect 41399 12021 41559 12033
rect 41399 11645 41405 12021
rect 41439 11645 41519 12021
rect 41553 11645 41559 12021
rect 41399 11633 41559 11645
rect 41771 12021 41931 12033
rect 41771 11645 41777 12021
rect 41811 11645 41891 12021
rect 41925 11645 41931 12021
rect 41771 11633 41931 11645
rect 42143 12021 42303 12033
rect 42143 11645 42149 12021
rect 42183 11645 42263 12021
rect 42297 11645 42303 12021
rect 42143 11633 42303 11645
rect 42515 12021 42675 12033
rect 42515 11645 42521 12021
rect 42555 11645 42635 12021
rect 42669 11645 42675 12021
rect 42515 11633 42675 11645
rect 42887 12021 43047 12033
rect 42887 11645 42893 12021
rect 42927 11645 43007 12021
rect 43041 11645 43047 12021
rect 42887 11633 43047 11645
rect 43259 12021 43419 12033
rect 43259 11645 43265 12021
rect 43299 11645 43379 12021
rect 43413 11645 43419 12021
rect 43259 11633 43419 11645
rect 43631 12021 43791 12033
rect 43631 11645 43637 12021
rect 43671 11645 43751 12021
rect 43785 11645 43791 12021
rect 43631 11633 43791 11645
rect 44003 12021 44163 12033
rect 44003 11645 44009 12021
rect 44043 11645 44123 12021
rect 44157 11645 44163 12021
rect 44003 11633 44163 11645
rect 44375 12021 44535 12033
rect 44375 11645 44381 12021
rect 44415 11645 44495 12021
rect 44529 11645 44535 12021
rect 44375 11633 44535 11645
rect 44747 12021 44907 12033
rect 44747 11645 44753 12021
rect 44787 11645 44867 12021
rect 44901 11645 44907 12021
rect 44747 11633 44907 11645
rect 45118 12021 45170 12073
rect 45118 11645 45125 12021
rect 45159 11645 45170 12021
rect 39280 11592 39366 11593
rect 39280 11587 39529 11592
rect 39280 11443 39348 11587
rect 39518 11546 39529 11587
rect 39518 11484 39528 11546
rect 39518 11443 39529 11484
rect 39280 11438 39529 11443
rect 39280 11437 39368 11438
rect 39280 11385 39328 11437
rect 39584 11397 39654 11633
rect 39709 11587 39901 11592
rect 39709 11546 39720 11587
rect 39710 11484 39720 11546
rect 39709 11443 39720 11484
rect 39890 11546 39901 11587
rect 39890 11484 39900 11546
rect 39890 11443 39901 11484
rect 39709 11438 39901 11443
rect 39956 11397 40026 11633
rect 40081 11587 40273 11592
rect 40081 11546 40092 11587
rect 40082 11484 40092 11546
rect 40081 11443 40092 11484
rect 40262 11546 40273 11587
rect 40262 11484 40272 11546
rect 40262 11443 40273 11484
rect 40081 11438 40273 11443
rect 40328 11397 40398 11633
rect 40453 11591 40645 11592
rect 40700 11591 40770 11633
rect 40825 11591 41017 11592
rect 40453 11587 41017 11591
rect 40453 11546 40464 11587
rect 40454 11484 40464 11546
rect 40453 11443 40464 11484
rect 40634 11443 40836 11587
rect 41006 11546 41017 11587
rect 41006 11484 41016 11546
rect 41006 11443 41017 11484
rect 40453 11439 41017 11443
rect 40453 11438 40645 11439
rect 40700 11397 40770 11439
rect 40825 11438 41017 11439
rect 41072 11397 41142 11633
rect 41197 11587 41389 11592
rect 41197 11546 41208 11587
rect 41198 11484 41208 11546
rect 41197 11443 41208 11484
rect 41378 11546 41389 11587
rect 41378 11484 41388 11546
rect 41378 11443 41389 11484
rect 41197 11438 41389 11443
rect 41444 11397 41514 11633
rect 41569 11587 41761 11592
rect 41569 11546 41580 11587
rect 41570 11484 41580 11546
rect 41569 11443 41580 11484
rect 41750 11546 41761 11587
rect 41750 11484 41760 11546
rect 41750 11443 41761 11484
rect 41569 11438 41761 11443
rect 41816 11397 41886 11633
rect 42188 11593 42258 11633
rect 41996 11592 42414 11593
rect 41941 11587 42505 11592
rect 41941 11546 41952 11587
rect 41942 11484 41952 11546
rect 41941 11443 41952 11484
rect 42122 11443 42324 11587
rect 42494 11546 42505 11587
rect 42494 11484 42504 11546
rect 42494 11443 42505 11484
rect 41941 11438 42505 11443
rect 41996 11437 42414 11438
rect 42188 11397 42258 11437
rect 42560 11397 42630 11633
rect 42685 11587 42877 11592
rect 42685 11546 42696 11587
rect 42686 11484 42696 11546
rect 42685 11443 42696 11484
rect 42866 11546 42877 11587
rect 42866 11484 42876 11546
rect 42866 11443 42877 11484
rect 42685 11438 42877 11443
rect 42932 11397 43002 11633
rect 43057 11587 43249 11592
rect 43057 11546 43068 11587
rect 43058 11484 43068 11546
rect 43057 11443 43068 11484
rect 43238 11546 43249 11587
rect 43238 11484 43248 11546
rect 43238 11443 43249 11484
rect 43057 11438 43249 11443
rect 43304 11397 43374 11633
rect 43676 11593 43746 11633
rect 43524 11592 43900 11593
rect 43429 11587 43993 11592
rect 43429 11546 43440 11587
rect 43430 11484 43440 11546
rect 43429 11443 43440 11484
rect 43610 11443 43812 11587
rect 43982 11546 43993 11587
rect 43982 11484 43992 11546
rect 43982 11443 43993 11484
rect 43429 11438 43993 11443
rect 43524 11437 43900 11438
rect 43676 11397 43746 11437
rect 44048 11397 44118 11633
rect 44173 11587 44365 11592
rect 44173 11546 44184 11587
rect 44174 11484 44184 11546
rect 44173 11443 44184 11484
rect 44354 11546 44365 11587
rect 44354 11484 44364 11546
rect 44354 11443 44365 11484
rect 44173 11438 44365 11443
rect 44420 11397 44490 11633
rect 44545 11587 44737 11592
rect 44545 11546 44556 11587
rect 44546 11484 44556 11546
rect 44545 11443 44556 11484
rect 44726 11546 44737 11587
rect 44726 11484 44736 11546
rect 44726 11443 44737 11484
rect 44545 11438 44737 11443
rect 44792 11397 44862 11633
rect 45118 11593 45170 11645
rect 45012 11592 45170 11593
rect 44917 11587 45170 11592
rect 44917 11546 44928 11587
rect 44918 11484 44928 11546
rect 44917 11443 44928 11484
rect 45098 11443 45170 11587
rect 44917 11438 45170 11443
rect 45012 11437 45170 11438
rect 39280 11009 39287 11385
rect 39321 11009 39328 11385
rect 39280 10963 39328 11009
rect 39539 11385 39699 11397
rect 39539 11009 39545 11385
rect 39579 11009 39659 11385
rect 39693 11009 39699 11385
rect 39539 10997 39699 11009
rect 39911 11385 40071 11397
rect 39911 11009 39917 11385
rect 39951 11009 40031 11385
rect 40065 11009 40071 11385
rect 39911 10997 40071 11009
rect 40283 11385 40443 11397
rect 40283 11009 40289 11385
rect 40323 11009 40403 11385
rect 40437 11009 40443 11385
rect 40283 10997 40443 11009
rect 40655 11385 40815 11397
rect 40655 11009 40661 11385
rect 40695 11009 40775 11385
rect 40809 11009 40815 11385
rect 40655 10997 40815 11009
rect 41027 11385 41187 11397
rect 41027 11009 41033 11385
rect 41067 11009 41147 11385
rect 41181 11009 41187 11385
rect 41027 10997 41187 11009
rect 41399 11385 41559 11397
rect 41399 11009 41405 11385
rect 41439 11009 41519 11385
rect 41553 11009 41559 11385
rect 41399 10997 41559 11009
rect 41771 11385 41931 11397
rect 41771 11009 41777 11385
rect 41811 11009 41891 11385
rect 41925 11009 41931 11385
rect 41771 10997 41931 11009
rect 42143 11385 42303 11397
rect 42143 11009 42149 11385
rect 42183 11009 42263 11385
rect 42297 11009 42303 11385
rect 42143 10997 42303 11009
rect 42515 11385 42675 11397
rect 42515 11009 42521 11385
rect 42555 11009 42635 11385
rect 42669 11009 42675 11385
rect 42515 10997 42675 11009
rect 42887 11385 43047 11397
rect 42887 11009 42893 11385
rect 42927 11009 43007 11385
rect 43041 11009 43047 11385
rect 42887 10997 43047 11009
rect 43259 11385 43419 11397
rect 43259 11009 43265 11385
rect 43299 11009 43379 11385
rect 43413 11009 43419 11385
rect 43259 10997 43419 11009
rect 43631 11385 43791 11397
rect 43631 11009 43637 11385
rect 43671 11009 43751 11385
rect 43785 11009 43791 11385
rect 43631 10997 43791 11009
rect 44003 11385 44163 11397
rect 44003 11009 44009 11385
rect 44043 11009 44123 11385
rect 44157 11009 44163 11385
rect 44003 10997 44163 11009
rect 44375 11385 44535 11397
rect 44375 11009 44381 11385
rect 44415 11009 44495 11385
rect 44529 11009 44535 11385
rect 44375 10997 44535 11009
rect 44747 11385 44907 11397
rect 44747 11009 44753 11385
rect 44787 11009 44867 11385
rect 44901 11009 44907 11385
rect 44747 10997 44907 11009
rect 45118 11385 45170 11437
rect 45118 11009 45125 11385
rect 45159 11009 45170 11385
rect 39280 10903 39348 10963
rect 39518 10956 39528 10963
rect 39518 10910 39529 10956
rect 39518 10903 39528 10910
rect 39590 10873 39648 10997
rect 39710 10956 39720 10963
rect 39709 10910 39720 10956
rect 39890 10956 39900 10963
rect 40082 10956 40092 10963
rect 39710 10903 39720 10910
rect 39890 10910 39901 10956
rect 40081 10910 40092 10956
rect 40262 10956 40272 10963
rect 39890 10903 39900 10910
rect 40082 10903 40092 10910
rect 40262 10910 40273 10956
rect 40262 10903 40272 10910
rect 40334 10873 40392 10997
rect 40706 10963 40764 10997
rect 40454 10956 40464 10963
rect 40453 10910 40464 10956
rect 40454 10903 40464 10910
rect 40634 10903 40836 10963
rect 41006 10956 41016 10963
rect 41006 10910 41017 10956
rect 41006 10903 41016 10910
rect 41078 10873 41136 10997
rect 41198 10956 41208 10963
rect 41197 10910 41208 10956
rect 41378 10956 41388 10963
rect 41570 10956 41580 10963
rect 41198 10903 41208 10910
rect 41378 10910 41389 10956
rect 41569 10910 41580 10956
rect 41750 10956 41760 10963
rect 41378 10903 41388 10910
rect 41570 10903 41580 10910
rect 41750 10910 41761 10956
rect 41750 10903 41760 10910
rect 41822 10873 41880 10997
rect 42194 10963 42252 10997
rect 41942 10956 41952 10963
rect 41941 10910 41952 10956
rect 41942 10903 41952 10910
rect 42122 10903 42324 10963
rect 42494 10956 42504 10963
rect 42494 10910 42505 10956
rect 42494 10903 42504 10910
rect 42566 10873 42624 10997
rect 42686 10956 42696 10963
rect 42685 10910 42696 10956
rect 42866 10956 42876 10963
rect 43058 10956 43068 10963
rect 42686 10903 42696 10910
rect 42866 10910 42877 10956
rect 43057 10910 43068 10956
rect 43238 10956 43248 10963
rect 42866 10903 42876 10910
rect 43058 10903 43068 10910
rect 43238 10910 43249 10956
rect 43238 10903 43248 10910
rect 43310 10873 43368 10997
rect 43682 10963 43740 10997
rect 43430 10956 43440 10963
rect 43429 10910 43440 10956
rect 43430 10903 43440 10910
rect 43610 10903 43812 10963
rect 43982 10956 43992 10963
rect 43982 10910 43993 10956
rect 43982 10903 43992 10910
rect 44054 10873 44112 10997
rect 44174 10956 44184 10963
rect 44173 10910 44184 10956
rect 44354 10956 44364 10963
rect 44546 10956 44556 10963
rect 44174 10903 44184 10910
rect 44354 10910 44365 10956
rect 44545 10910 44556 10956
rect 44726 10956 44736 10963
rect 44354 10903 44364 10910
rect 44546 10903 44556 10910
rect 44726 10910 44737 10956
rect 44726 10903 44736 10910
rect 44798 10873 44856 10997
rect 45118 10963 45170 11009
rect 44918 10956 44928 10963
rect 44917 10910 44928 10956
rect 44918 10903 44928 10910
rect 45098 10903 45170 10963
rect 45208 12657 45279 12669
rect 45208 12281 45239 12657
rect 45273 12281 45279 12657
rect 45208 12269 45279 12281
rect 45491 12657 45651 12669
rect 45491 12281 45497 12657
rect 45531 12281 45611 12657
rect 45645 12281 45651 12657
rect 45491 12269 45651 12281
rect 45863 12657 46023 12669
rect 45863 12281 45869 12657
rect 45903 12281 45983 12657
rect 46017 12281 46023 12657
rect 45863 12269 46023 12281
rect 46235 12657 46395 12669
rect 46235 12281 46241 12657
rect 46275 12281 46355 12657
rect 46389 12281 46395 12657
rect 46235 12269 46395 12281
rect 46607 12657 46767 12669
rect 46607 12281 46613 12657
rect 46647 12281 46727 12657
rect 46761 12281 46767 12657
rect 46607 12269 46767 12281
rect 46979 12657 47139 12669
rect 46979 12281 46985 12657
rect 47019 12281 47099 12657
rect 47133 12281 47139 12657
rect 46979 12269 47139 12281
rect 47351 12657 47511 12669
rect 47351 12281 47357 12657
rect 47391 12281 47471 12657
rect 47505 12281 47511 12657
rect 47351 12269 47511 12281
rect 47723 12657 47883 12669
rect 47723 12281 47729 12657
rect 47763 12281 47843 12657
rect 47877 12281 47883 12657
rect 47723 12269 47883 12281
rect 48095 12657 48255 12669
rect 48095 12281 48101 12657
rect 48135 12281 48215 12657
rect 48249 12281 48255 12657
rect 48095 12269 48255 12281
rect 48467 12657 48627 12669
rect 48467 12281 48473 12657
rect 48507 12281 48587 12657
rect 48621 12281 48627 12657
rect 48467 12269 48627 12281
rect 48839 12657 48999 12669
rect 48839 12281 48845 12657
rect 48879 12281 48959 12657
rect 48993 12281 48999 12657
rect 48839 12269 48999 12281
rect 49211 12657 49371 12669
rect 49211 12281 49217 12657
rect 49251 12281 49331 12657
rect 49365 12281 49371 12657
rect 49211 12269 49371 12281
rect 49583 12657 49743 12669
rect 49583 12281 49589 12657
rect 49623 12281 49703 12657
rect 49737 12281 49743 12657
rect 49583 12269 49743 12281
rect 49955 12657 50115 12669
rect 49955 12281 49961 12657
rect 49995 12281 50075 12657
rect 50109 12281 50115 12657
rect 49955 12269 50115 12281
rect 50327 12657 50487 12669
rect 50327 12281 50333 12657
rect 50367 12281 50447 12657
rect 50481 12281 50487 12657
rect 50327 12269 50487 12281
rect 50699 12657 50859 12669
rect 50699 12281 50705 12657
rect 50739 12281 50819 12657
rect 50853 12281 50859 12657
rect 50699 12269 50859 12281
rect 51071 12657 51162 12669
rect 51071 12281 51077 12657
rect 51111 12281 51162 12657
rect 51071 12269 51162 12281
rect 45208 12033 45260 12269
rect 45288 12228 45430 12229
rect 45288 12223 45481 12228
rect 45288 12079 45300 12223
rect 45470 12182 45481 12223
rect 45470 12120 45480 12182
rect 45470 12079 45481 12120
rect 45288 12074 45481 12079
rect 45288 12073 45430 12074
rect 45536 12033 45606 12269
rect 45661 12223 45853 12228
rect 45661 12182 45672 12223
rect 45662 12120 45672 12182
rect 45661 12079 45672 12120
rect 45842 12182 45853 12223
rect 45842 12120 45852 12182
rect 45842 12079 45853 12120
rect 45661 12074 45853 12079
rect 45908 12033 45978 12269
rect 46033 12223 46225 12228
rect 46033 12182 46044 12223
rect 46034 12120 46044 12182
rect 46033 12079 46044 12120
rect 46214 12182 46225 12223
rect 46214 12120 46224 12182
rect 46214 12079 46225 12120
rect 46033 12074 46225 12079
rect 46280 12033 46350 12269
rect 46405 12223 46597 12228
rect 46405 12182 46416 12223
rect 46406 12120 46416 12182
rect 46405 12079 46416 12120
rect 46586 12182 46597 12223
rect 46586 12120 46596 12182
rect 46586 12079 46597 12120
rect 46405 12074 46597 12079
rect 46652 12033 46722 12269
rect 46777 12223 46969 12228
rect 46777 12182 46788 12223
rect 46778 12120 46788 12182
rect 46777 12079 46788 12120
rect 46958 12182 46969 12223
rect 46958 12120 46968 12182
rect 46958 12079 46969 12120
rect 46777 12074 46969 12079
rect 47024 12033 47094 12269
rect 47149 12223 47341 12228
rect 47149 12182 47160 12223
rect 47150 12120 47160 12182
rect 47149 12079 47160 12120
rect 47330 12182 47341 12223
rect 47330 12120 47340 12182
rect 47330 12079 47341 12120
rect 47149 12074 47341 12079
rect 47396 12033 47466 12269
rect 47521 12223 47713 12228
rect 47521 12182 47532 12223
rect 47522 12120 47532 12182
rect 47521 12079 47532 12120
rect 47702 12182 47713 12223
rect 47702 12120 47712 12182
rect 47702 12079 47713 12120
rect 47521 12074 47713 12079
rect 47768 12033 47838 12269
rect 47893 12223 48085 12228
rect 47893 12182 47904 12223
rect 47894 12120 47904 12182
rect 47893 12079 47904 12120
rect 48074 12182 48085 12223
rect 48074 12120 48084 12182
rect 48074 12079 48085 12120
rect 47893 12074 48085 12079
rect 48140 12033 48210 12269
rect 48265 12223 48457 12228
rect 48265 12182 48276 12223
rect 48266 12120 48276 12182
rect 48265 12079 48276 12120
rect 48446 12182 48457 12223
rect 48446 12120 48456 12182
rect 48446 12079 48457 12120
rect 48265 12074 48457 12079
rect 48512 12033 48582 12269
rect 48637 12223 48829 12228
rect 48637 12182 48648 12223
rect 48638 12120 48648 12182
rect 48637 12079 48648 12120
rect 48818 12182 48829 12223
rect 48818 12120 48828 12182
rect 48818 12079 48829 12120
rect 48637 12074 48829 12079
rect 48884 12033 48954 12269
rect 49009 12223 49201 12228
rect 49009 12182 49020 12223
rect 49010 12120 49020 12182
rect 49009 12079 49020 12120
rect 49190 12182 49201 12223
rect 49190 12120 49200 12182
rect 49190 12079 49201 12120
rect 49009 12074 49201 12079
rect 49256 12033 49326 12269
rect 49381 12223 49573 12228
rect 49381 12182 49392 12223
rect 49382 12120 49392 12182
rect 49381 12079 49392 12120
rect 49562 12182 49573 12223
rect 49562 12120 49572 12182
rect 49562 12079 49573 12120
rect 49381 12074 49573 12079
rect 49628 12033 49698 12269
rect 49753 12223 49945 12228
rect 49753 12182 49764 12223
rect 49754 12120 49764 12182
rect 49753 12079 49764 12120
rect 49934 12182 49945 12223
rect 49934 12120 49944 12182
rect 49934 12079 49945 12120
rect 49753 12074 49945 12079
rect 50000 12033 50070 12269
rect 50125 12223 50317 12228
rect 50125 12182 50136 12223
rect 50126 12120 50136 12182
rect 50125 12079 50136 12120
rect 50306 12182 50317 12223
rect 50306 12120 50316 12182
rect 50306 12079 50317 12120
rect 50125 12074 50317 12079
rect 50372 12033 50442 12269
rect 50497 12223 50689 12228
rect 50497 12182 50508 12223
rect 50498 12120 50508 12182
rect 50497 12079 50508 12120
rect 50678 12182 50689 12223
rect 50678 12120 50688 12182
rect 50678 12079 50689 12120
rect 50497 12074 50689 12079
rect 50744 12033 50814 12269
rect 50869 12223 51061 12228
rect 50869 12182 50880 12223
rect 50870 12120 50880 12182
rect 50869 12079 50880 12120
rect 51050 12182 51061 12223
rect 51050 12120 51060 12182
rect 51050 12079 51061 12120
rect 50869 12074 51061 12079
rect 51104 12033 51162 12269
rect 45208 12021 45279 12033
rect 45208 11645 45239 12021
rect 45273 11645 45279 12021
rect 45208 11633 45279 11645
rect 45491 12021 45651 12033
rect 45491 11645 45497 12021
rect 45531 11645 45611 12021
rect 45645 11645 45651 12021
rect 45491 11633 45651 11645
rect 45863 12021 46023 12033
rect 45863 11645 45869 12021
rect 45903 11645 45983 12021
rect 46017 11645 46023 12021
rect 45863 11633 46023 11645
rect 46235 12021 46395 12033
rect 46235 11645 46241 12021
rect 46275 11645 46355 12021
rect 46389 11645 46395 12021
rect 46235 11633 46395 11645
rect 46607 12021 46767 12033
rect 46607 11645 46613 12021
rect 46647 11645 46727 12021
rect 46761 11645 46767 12021
rect 46607 11633 46767 11645
rect 46979 12021 47139 12033
rect 46979 11645 46985 12021
rect 47019 11645 47099 12021
rect 47133 11645 47139 12021
rect 46979 11633 47139 11645
rect 47351 12021 47511 12033
rect 47351 11645 47357 12021
rect 47391 11645 47471 12021
rect 47505 11645 47511 12021
rect 47351 11633 47511 11645
rect 47723 12021 47883 12033
rect 47723 11645 47729 12021
rect 47763 11645 47843 12021
rect 47877 11645 47883 12021
rect 47723 11633 47883 11645
rect 48095 12021 48255 12033
rect 48095 11645 48101 12021
rect 48135 11645 48215 12021
rect 48249 11645 48255 12021
rect 48095 11633 48255 11645
rect 48467 12021 48627 12033
rect 48467 11645 48473 12021
rect 48507 11645 48587 12021
rect 48621 11645 48627 12021
rect 48467 11633 48627 11645
rect 48839 12021 48999 12033
rect 48839 11645 48845 12021
rect 48879 11645 48959 12021
rect 48993 11645 48999 12021
rect 48839 11633 48999 11645
rect 49211 12021 49371 12033
rect 49211 11645 49217 12021
rect 49251 11645 49331 12021
rect 49365 11645 49371 12021
rect 49211 11633 49371 11645
rect 49583 12021 49743 12033
rect 49583 11645 49589 12021
rect 49623 11645 49703 12021
rect 49737 11645 49743 12021
rect 49583 11633 49743 11645
rect 49955 12021 50115 12033
rect 49955 11645 49961 12021
rect 49995 11645 50075 12021
rect 50109 11645 50115 12021
rect 49955 11633 50115 11645
rect 50327 12021 50487 12033
rect 50327 11645 50333 12021
rect 50367 11645 50447 12021
rect 50481 11645 50487 12021
rect 50327 11633 50487 11645
rect 50699 12021 50859 12033
rect 50699 11645 50705 12021
rect 50739 11645 50819 12021
rect 50853 11645 50859 12021
rect 50699 11633 50859 11645
rect 51071 12021 51162 12033
rect 51071 11645 51077 12021
rect 51111 11645 51162 12021
rect 51071 11633 51162 11645
rect 45208 11397 45260 11633
rect 45288 11592 45414 11593
rect 45288 11587 45481 11592
rect 45288 11443 45300 11587
rect 45470 11546 45481 11587
rect 45470 11484 45480 11546
rect 45470 11443 45481 11484
rect 45288 11438 45481 11443
rect 45288 11437 45414 11438
rect 45536 11397 45606 11633
rect 45661 11587 45853 11592
rect 45661 11546 45672 11587
rect 45662 11484 45672 11546
rect 45661 11443 45672 11484
rect 45842 11546 45853 11587
rect 45842 11484 45852 11546
rect 45842 11443 45853 11484
rect 45661 11438 45853 11443
rect 45908 11397 45978 11633
rect 46033 11587 46225 11592
rect 46033 11546 46044 11587
rect 46034 11484 46044 11546
rect 46033 11443 46044 11484
rect 46214 11546 46225 11587
rect 46214 11484 46224 11546
rect 46214 11443 46225 11484
rect 46033 11438 46225 11443
rect 46280 11397 46350 11633
rect 46405 11587 46597 11592
rect 46405 11546 46416 11587
rect 46406 11484 46416 11546
rect 46405 11443 46416 11484
rect 46586 11546 46597 11587
rect 46586 11484 46596 11546
rect 46586 11443 46597 11484
rect 46405 11438 46597 11443
rect 46652 11397 46722 11633
rect 46777 11587 46969 11592
rect 46777 11546 46788 11587
rect 46778 11484 46788 11546
rect 46777 11443 46788 11484
rect 46958 11546 46969 11587
rect 46958 11484 46968 11546
rect 46958 11443 46969 11484
rect 46777 11438 46969 11443
rect 47024 11397 47094 11633
rect 47149 11587 47341 11592
rect 47149 11546 47160 11587
rect 47150 11484 47160 11546
rect 47149 11443 47160 11484
rect 47330 11546 47341 11587
rect 47330 11484 47340 11546
rect 47330 11443 47341 11484
rect 47149 11438 47341 11443
rect 47396 11397 47466 11633
rect 47521 11587 47713 11592
rect 47521 11546 47532 11587
rect 47522 11484 47532 11546
rect 47521 11443 47532 11484
rect 47702 11546 47713 11587
rect 47702 11484 47712 11546
rect 47702 11443 47713 11484
rect 47521 11438 47713 11443
rect 47768 11397 47838 11633
rect 47893 11587 48085 11592
rect 47893 11546 47904 11587
rect 47894 11484 47904 11546
rect 47893 11443 47904 11484
rect 48074 11546 48085 11587
rect 48074 11484 48084 11546
rect 48074 11443 48085 11484
rect 47893 11438 48085 11443
rect 48140 11397 48210 11633
rect 48265 11587 48457 11592
rect 48265 11546 48276 11587
rect 48266 11484 48276 11546
rect 48265 11443 48276 11484
rect 48446 11546 48457 11587
rect 48446 11484 48456 11546
rect 48446 11443 48457 11484
rect 48265 11438 48457 11443
rect 48512 11397 48582 11633
rect 48637 11587 48829 11592
rect 48637 11546 48648 11587
rect 48638 11484 48648 11546
rect 48637 11443 48648 11484
rect 48818 11546 48829 11587
rect 48818 11484 48828 11546
rect 48818 11443 48829 11484
rect 48637 11438 48829 11443
rect 48884 11397 48954 11633
rect 49009 11587 49201 11592
rect 49009 11546 49020 11587
rect 49010 11484 49020 11546
rect 49009 11443 49020 11484
rect 49190 11546 49201 11587
rect 49190 11484 49200 11546
rect 49190 11443 49201 11484
rect 49009 11438 49201 11443
rect 49256 11397 49326 11633
rect 49381 11587 49573 11592
rect 49381 11546 49392 11587
rect 49382 11484 49392 11546
rect 49381 11443 49392 11484
rect 49562 11546 49573 11587
rect 49562 11484 49572 11546
rect 49562 11443 49573 11484
rect 49381 11438 49573 11443
rect 49628 11397 49698 11633
rect 49753 11587 49945 11592
rect 49753 11546 49764 11587
rect 49754 11484 49764 11546
rect 49753 11443 49764 11484
rect 49934 11546 49945 11587
rect 49934 11484 49944 11546
rect 49934 11443 49945 11484
rect 49753 11438 49945 11443
rect 50000 11397 50070 11633
rect 50125 11587 50317 11592
rect 50125 11546 50136 11587
rect 50126 11484 50136 11546
rect 50125 11443 50136 11484
rect 50306 11546 50317 11587
rect 50306 11484 50316 11546
rect 50306 11443 50317 11484
rect 50125 11438 50317 11443
rect 50372 11397 50442 11633
rect 50497 11587 50689 11592
rect 50497 11546 50508 11587
rect 50498 11484 50508 11546
rect 50497 11443 50508 11484
rect 50678 11546 50689 11587
rect 50678 11484 50688 11546
rect 50678 11443 50689 11484
rect 50497 11438 50689 11443
rect 50744 11397 50814 11633
rect 50869 11587 51061 11592
rect 50869 11546 50880 11587
rect 50870 11484 50880 11546
rect 50869 11443 50880 11484
rect 51050 11546 51061 11587
rect 51050 11484 51060 11546
rect 51050 11443 51061 11484
rect 50869 11438 51061 11443
rect 51104 11397 51162 11633
rect 45208 11385 45279 11397
rect 45208 11009 45239 11385
rect 45273 11009 45279 11385
rect 45208 10997 45279 11009
rect 45491 11385 45651 11397
rect 45491 11009 45497 11385
rect 45531 11009 45611 11385
rect 45645 11009 45651 11385
rect 45491 10997 45651 11009
rect 45863 11385 46023 11397
rect 45863 11009 45869 11385
rect 45903 11009 45983 11385
rect 46017 11009 46023 11385
rect 45863 10997 46023 11009
rect 46235 11385 46395 11397
rect 46235 11009 46241 11385
rect 46275 11009 46355 11385
rect 46389 11009 46395 11385
rect 46235 10997 46395 11009
rect 46607 11385 46767 11397
rect 46607 11009 46613 11385
rect 46647 11009 46727 11385
rect 46761 11009 46767 11385
rect 46607 10997 46767 11009
rect 46979 11385 47139 11397
rect 46979 11009 46985 11385
rect 47019 11009 47099 11385
rect 47133 11009 47139 11385
rect 46979 10997 47139 11009
rect 47351 11385 47511 11397
rect 47351 11009 47357 11385
rect 47391 11009 47471 11385
rect 47505 11009 47511 11385
rect 47351 10997 47511 11009
rect 47723 11385 47883 11397
rect 47723 11009 47729 11385
rect 47763 11009 47843 11385
rect 47877 11009 47883 11385
rect 47723 10997 47883 11009
rect 48095 11385 48255 11397
rect 48095 11009 48101 11385
rect 48135 11009 48215 11385
rect 48249 11009 48255 11385
rect 48095 10997 48255 11009
rect 48467 11385 48627 11397
rect 48467 11009 48473 11385
rect 48507 11009 48587 11385
rect 48621 11009 48627 11385
rect 48467 10997 48627 11009
rect 48839 11385 48999 11397
rect 48839 11009 48845 11385
rect 48879 11009 48959 11385
rect 48993 11009 48999 11385
rect 48839 10997 48999 11009
rect 49211 11385 49371 11397
rect 49211 11009 49217 11385
rect 49251 11009 49331 11385
rect 49365 11009 49371 11385
rect 49211 10997 49371 11009
rect 49583 11385 49743 11397
rect 49583 11009 49589 11385
rect 49623 11009 49703 11385
rect 49737 11009 49743 11385
rect 49583 10997 49743 11009
rect 49955 11385 50115 11397
rect 49955 11009 49961 11385
rect 49995 11009 50075 11385
rect 50109 11009 50115 11385
rect 49955 10997 50115 11009
rect 50327 11385 50487 11397
rect 50327 11009 50333 11385
rect 50367 11009 50447 11385
rect 50481 11009 50487 11385
rect 50327 10997 50487 11009
rect 50699 11385 50859 11397
rect 50699 11009 50705 11385
rect 50739 11009 50819 11385
rect 50853 11009 50859 11385
rect 50699 10997 50859 11009
rect 51071 11385 51162 11397
rect 51071 11009 51077 11385
rect 51111 11009 51162 11385
rect 51071 10997 51162 11009
rect 45208 10873 45260 10997
rect 45294 10903 45300 10963
rect 45470 10956 45480 10963
rect 45662 10956 45672 10963
rect 45470 10910 45481 10956
rect 45661 10910 45672 10956
rect 45842 10956 45852 10963
rect 45470 10903 45480 10910
rect 45662 10903 45672 10910
rect 45842 10910 45853 10956
rect 45842 10903 45852 10910
rect 45914 10873 45972 10997
rect 46034 10956 46044 10963
rect 46033 10910 46044 10956
rect 46214 10956 46224 10963
rect 46406 10956 46416 10963
rect 46034 10903 46044 10910
rect 46214 10910 46225 10956
rect 46405 10910 46416 10956
rect 46586 10956 46596 10963
rect 46214 10903 46224 10910
rect 46406 10903 46416 10910
rect 46586 10910 46597 10956
rect 46586 10903 46596 10910
rect 46658 10873 46716 10997
rect 46778 10956 46788 10963
rect 46777 10910 46788 10956
rect 46958 10956 46968 10963
rect 47150 10956 47160 10963
rect 46778 10903 46788 10910
rect 46958 10910 46969 10956
rect 47149 10910 47160 10956
rect 47330 10956 47340 10963
rect 46958 10903 46968 10910
rect 47150 10903 47160 10910
rect 47330 10910 47341 10956
rect 47330 10903 47340 10910
rect 47402 10873 47460 10997
rect 47522 10956 47532 10963
rect 47521 10910 47532 10956
rect 47702 10956 47712 10963
rect 47894 10956 47904 10963
rect 47522 10903 47532 10910
rect 47702 10910 47713 10956
rect 47893 10910 47904 10956
rect 48074 10956 48084 10963
rect 47702 10903 47712 10910
rect 47894 10903 47904 10910
rect 48074 10910 48085 10956
rect 48074 10903 48084 10910
rect 48146 10873 48204 10997
rect 48266 10956 48276 10963
rect 48265 10910 48276 10956
rect 48446 10956 48456 10963
rect 48638 10956 48648 10963
rect 48266 10903 48276 10910
rect 48446 10910 48457 10956
rect 48637 10910 48648 10956
rect 48818 10956 48828 10963
rect 48446 10903 48456 10910
rect 48638 10903 48648 10910
rect 48818 10910 48829 10956
rect 48818 10903 48828 10910
rect 48890 10873 48948 10997
rect 49010 10956 49020 10963
rect 49009 10910 49020 10956
rect 49190 10956 49200 10963
rect 49382 10956 49392 10963
rect 49010 10903 49020 10910
rect 49190 10910 49201 10956
rect 49381 10910 49392 10956
rect 49562 10956 49572 10963
rect 49190 10903 49200 10910
rect 49382 10903 49392 10910
rect 49562 10910 49573 10956
rect 49562 10903 49572 10910
rect 49634 10873 49692 10997
rect 49754 10956 49764 10963
rect 49753 10910 49764 10956
rect 49934 10956 49944 10963
rect 50126 10956 50136 10963
rect 49754 10903 49764 10910
rect 49934 10910 49945 10956
rect 50125 10910 50136 10956
rect 50306 10956 50316 10963
rect 49934 10903 49944 10910
rect 50126 10903 50136 10910
rect 50306 10910 50317 10956
rect 50306 10903 50316 10910
rect 50378 10873 50436 10997
rect 50498 10956 50508 10963
rect 50497 10910 50508 10956
rect 50678 10956 50688 10963
rect 50870 10956 50880 10963
rect 50498 10903 50508 10910
rect 50678 10910 50689 10956
rect 50869 10910 50880 10956
rect 51050 10956 51060 10963
rect 50678 10903 50688 10910
rect 50870 10903 50880 10910
rect 51050 10910 51061 10956
rect 51050 10903 51060 10910
rect 51104 10873 51162 10997
rect 39572 10867 39666 10873
rect 39572 10797 39584 10867
rect 39654 10797 39666 10867
rect 39572 10791 39666 10797
rect 40316 10867 40410 10873
rect 40316 10797 40328 10867
rect 40398 10797 40410 10867
rect 40316 10791 40410 10797
rect 41060 10867 41154 10873
rect 41060 10797 41072 10867
rect 41142 10797 41154 10867
rect 41060 10791 41154 10797
rect 41804 10867 41898 10873
rect 41804 10797 41816 10867
rect 41886 10797 41898 10867
rect 41804 10791 41898 10797
rect 42548 10867 42642 10873
rect 42548 10797 42560 10867
rect 42630 10797 42642 10867
rect 42548 10791 42642 10797
rect 43292 10867 43386 10873
rect 43292 10797 43304 10867
rect 43374 10797 43386 10867
rect 43292 10791 43386 10797
rect 44036 10867 44130 10873
rect 44036 10797 44048 10867
rect 44118 10797 44130 10867
rect 44036 10791 44130 10797
rect 44780 10867 44874 10873
rect 44780 10797 44792 10867
rect 44862 10797 44874 10867
rect 44780 10791 44874 10797
rect 45152 10867 45260 10873
rect 45152 10797 45164 10867
rect 45234 10797 45260 10867
rect 45152 10791 45260 10797
rect 45896 10867 45990 10873
rect 45896 10797 45908 10867
rect 45978 10797 45990 10867
rect 45896 10791 45990 10797
rect 46640 10867 46734 10873
rect 46640 10797 46652 10867
rect 46722 10797 46734 10867
rect 46640 10791 46734 10797
rect 47384 10867 47478 10873
rect 47384 10797 47396 10867
rect 47466 10797 47478 10867
rect 47384 10791 47478 10797
rect 48128 10867 48222 10873
rect 48128 10797 48140 10867
rect 48210 10797 48222 10867
rect 48128 10791 48222 10797
rect 48872 10867 48966 10873
rect 48872 10797 48884 10867
rect 48954 10797 48966 10867
rect 48872 10791 48966 10797
rect 49616 10867 49710 10873
rect 49616 10797 49628 10867
rect 49698 10797 49710 10867
rect 49616 10791 49710 10797
rect 50360 10867 50454 10873
rect 50360 10797 50372 10867
rect 50442 10797 50454 10867
rect 50360 10791 50454 10797
rect 51050 10867 51162 10873
rect 51050 10797 51062 10867
rect 51132 10797 51162 10867
rect 51050 10791 51162 10797
rect 39590 10715 39648 10791
rect 40334 10715 40392 10791
rect 41078 10715 41136 10791
rect 41822 10715 41880 10791
rect 42566 10715 42624 10791
rect 43310 10715 43368 10791
rect 44054 10715 44112 10791
rect 44798 10725 44856 10791
rect 44778 10715 44856 10725
rect 45208 10715 45260 10791
rect 45914 10715 45972 10791
rect 46658 10715 46716 10791
rect 47402 10715 47460 10791
rect 48146 10715 48204 10791
rect 48890 10715 48948 10791
rect 49634 10715 49692 10791
rect 50378 10715 50436 10791
rect 51104 10731 51162 10791
rect 51104 10715 51180 10731
rect 39508 10515 39518 10715
rect 39718 10515 39728 10715
rect 40252 10515 40262 10715
rect 40462 10515 40472 10715
rect 40996 10515 41006 10715
rect 41206 10515 41216 10715
rect 41740 10515 41750 10715
rect 41950 10515 41960 10715
rect 42484 10515 42494 10715
rect 42694 10515 42704 10715
rect 43228 10515 43238 10715
rect 43438 10515 43448 10715
rect 43972 10515 43982 10715
rect 44182 10515 44192 10715
rect 44716 10515 44726 10715
rect 44926 10515 44936 10715
rect 45088 10515 45098 10715
rect 45298 10515 45308 10715
rect 45832 10515 45842 10715
rect 46042 10515 46052 10715
rect 46576 10515 46586 10715
rect 46786 10515 46796 10715
rect 47320 10515 47330 10715
rect 47530 10515 47540 10715
rect 48064 10515 48074 10715
rect 48274 10515 48284 10715
rect 48808 10515 48818 10715
rect 49018 10515 49028 10715
rect 49552 10515 49562 10715
rect 49762 10515 49772 10715
rect 50296 10515 50306 10715
rect 50506 10515 50516 10715
rect 51040 10515 51050 10715
rect 51250 10515 51260 10715
rect 39508 9150 39518 9350
rect 39718 9150 39728 9350
rect 40252 9150 40262 9350
rect 40462 9150 40472 9350
rect 40996 9150 41006 9350
rect 41206 9150 41216 9350
rect 41740 9150 41750 9350
rect 41950 9150 41960 9350
rect 42484 9150 42494 9350
rect 42694 9150 42704 9350
rect 43228 9150 43238 9350
rect 43438 9150 43448 9350
rect 43972 9150 43982 9350
rect 44182 9150 44192 9350
rect 44716 9150 44726 9350
rect 44926 9150 44936 9350
rect 45088 9150 45098 9350
rect 45298 9150 45308 9350
rect 45832 9150 45842 9350
rect 46042 9150 46052 9350
rect 46576 9150 46586 9350
rect 46786 9150 46796 9350
rect 47320 9150 47330 9350
rect 47530 9150 47540 9350
rect 48064 9150 48074 9350
rect 48274 9150 48284 9350
rect 48808 9150 48818 9350
rect 49018 9150 49028 9350
rect 49552 9150 49562 9350
rect 49762 9150 49772 9350
rect 50296 9150 50306 9350
rect 50506 9150 50516 9350
rect 51040 9150 51050 9350
rect 51250 9150 51260 9350
rect 39590 9074 39648 9150
rect 40334 9074 40392 9150
rect 41078 9074 41136 9150
rect 41822 9074 41880 9150
rect 42566 9074 42624 9150
rect 43310 9074 43368 9150
rect 44054 9074 44112 9150
rect 44778 9140 44856 9150
rect 44798 9074 44856 9140
rect 45208 9074 45260 9150
rect 45914 9074 45972 9150
rect 46658 9074 46716 9150
rect 47402 9074 47460 9150
rect 48146 9074 48204 9150
rect 48890 9074 48948 9150
rect 49634 9074 49692 9150
rect 50378 9074 50436 9150
rect 51104 9134 51180 9150
rect 51104 9074 51162 9134
rect 39572 9068 39666 9074
rect 39572 8998 39584 9068
rect 39654 8998 39666 9068
rect 39572 8992 39666 8998
rect 40316 9068 40410 9074
rect 40316 8998 40328 9068
rect 40398 8998 40410 9068
rect 40316 8992 40410 8998
rect 41060 9068 41154 9074
rect 41060 8998 41072 9068
rect 41142 8998 41154 9068
rect 41060 8992 41154 8998
rect 41804 9068 41898 9074
rect 41804 8998 41816 9068
rect 41886 8998 41898 9068
rect 41804 8992 41898 8998
rect 42548 9068 42642 9074
rect 42548 8998 42560 9068
rect 42630 8998 42642 9068
rect 42548 8992 42642 8998
rect 43292 9068 43386 9074
rect 43292 8998 43304 9068
rect 43374 8998 43386 9068
rect 43292 8992 43386 8998
rect 44036 9068 44130 9074
rect 44036 8998 44048 9068
rect 44118 8998 44130 9068
rect 44036 8992 44130 8998
rect 44780 9068 44874 9074
rect 44780 8998 44792 9068
rect 44862 8998 44874 9068
rect 44780 8992 44874 8998
rect 45152 9068 45260 9074
rect 45152 8998 45164 9068
rect 45234 8998 45260 9068
rect 45152 8992 45260 8998
rect 45896 9068 45990 9074
rect 45896 8998 45908 9068
rect 45978 8998 45990 9068
rect 45896 8992 45990 8998
rect 46640 9068 46734 9074
rect 46640 8998 46652 9068
rect 46722 8998 46734 9068
rect 46640 8992 46734 8998
rect 47384 9068 47478 9074
rect 47384 8998 47396 9068
rect 47466 8998 47478 9068
rect 47384 8992 47478 8998
rect 48128 9068 48222 9074
rect 48128 8998 48140 9068
rect 48210 8998 48222 9068
rect 48128 8992 48222 8998
rect 48872 9068 48966 9074
rect 48872 8998 48884 9068
rect 48954 8998 48966 9068
rect 48872 8992 48966 8998
rect 49616 9068 49710 9074
rect 49616 8998 49628 9068
rect 49698 8998 49710 9068
rect 49616 8992 49710 8998
rect 50360 9068 50454 9074
rect 50360 8998 50372 9068
rect 50442 8998 50454 9068
rect 50360 8992 50454 8998
rect 51050 9068 51162 9074
rect 51050 8998 51062 9068
rect 51132 8998 51162 9068
rect 51050 8992 51162 8998
rect 39280 8902 39348 8962
rect 39518 8955 39528 8962
rect 39518 8909 39529 8955
rect 39518 8902 39528 8909
rect 39280 8856 39328 8902
rect 39590 8868 39648 8992
rect 39710 8955 39720 8962
rect 39709 8909 39720 8955
rect 39890 8955 39900 8962
rect 40082 8955 40092 8962
rect 39710 8902 39720 8909
rect 39890 8909 39901 8955
rect 40081 8909 40092 8955
rect 40262 8955 40272 8962
rect 39890 8902 39900 8909
rect 40082 8902 40092 8909
rect 40262 8909 40273 8955
rect 40262 8902 40272 8909
rect 40334 8868 40392 8992
rect 40454 8955 40464 8962
rect 40453 8909 40464 8955
rect 40454 8902 40464 8909
rect 40634 8902 40836 8962
rect 41006 8955 41016 8962
rect 41006 8909 41017 8955
rect 41006 8902 41016 8909
rect 40706 8868 40764 8902
rect 41078 8868 41136 8992
rect 41198 8955 41208 8962
rect 41197 8909 41208 8955
rect 41378 8955 41388 8962
rect 41570 8955 41580 8962
rect 41198 8902 41208 8909
rect 41378 8909 41389 8955
rect 41569 8909 41580 8955
rect 41750 8955 41760 8962
rect 41378 8902 41388 8909
rect 41570 8902 41580 8909
rect 41750 8909 41761 8955
rect 41750 8902 41760 8909
rect 41822 8868 41880 8992
rect 41942 8955 41952 8962
rect 41941 8909 41952 8955
rect 41942 8902 41952 8909
rect 42122 8902 42324 8962
rect 42494 8955 42504 8962
rect 42494 8909 42505 8955
rect 42494 8902 42504 8909
rect 42194 8868 42252 8902
rect 42566 8868 42624 8992
rect 42686 8955 42696 8962
rect 42685 8909 42696 8955
rect 42866 8955 42876 8962
rect 43058 8955 43068 8962
rect 42686 8902 42696 8909
rect 42866 8909 42877 8955
rect 43057 8909 43068 8955
rect 43238 8955 43248 8962
rect 42866 8902 42876 8909
rect 43058 8902 43068 8909
rect 43238 8909 43249 8955
rect 43238 8902 43248 8909
rect 43310 8868 43368 8992
rect 43430 8955 43440 8962
rect 43429 8909 43440 8955
rect 43430 8902 43440 8909
rect 43610 8902 43812 8962
rect 43982 8955 43992 8962
rect 43982 8909 43993 8955
rect 43982 8902 43992 8909
rect 43682 8868 43740 8902
rect 44054 8868 44112 8992
rect 44174 8955 44184 8962
rect 44173 8909 44184 8955
rect 44354 8955 44364 8962
rect 44546 8955 44556 8962
rect 44174 8902 44184 8909
rect 44354 8909 44365 8955
rect 44545 8909 44556 8955
rect 44726 8955 44736 8962
rect 44354 8902 44364 8909
rect 44546 8902 44556 8909
rect 44726 8909 44737 8955
rect 44726 8902 44736 8909
rect 44798 8868 44856 8992
rect 44918 8955 44928 8962
rect 44917 8909 44928 8955
rect 44918 8902 44928 8909
rect 45098 8902 45170 8962
rect 39280 8480 39287 8856
rect 39321 8480 39328 8856
rect 39280 8428 39328 8480
rect 39539 8856 39699 8868
rect 39539 8480 39545 8856
rect 39579 8480 39659 8856
rect 39693 8480 39699 8856
rect 39539 8468 39699 8480
rect 39911 8856 40071 8868
rect 39911 8480 39917 8856
rect 39951 8480 40031 8856
rect 40065 8480 40071 8856
rect 39911 8468 40071 8480
rect 40283 8856 40443 8868
rect 40283 8480 40289 8856
rect 40323 8480 40403 8856
rect 40437 8480 40443 8856
rect 40283 8468 40443 8480
rect 40655 8856 40815 8868
rect 40655 8480 40661 8856
rect 40695 8480 40775 8856
rect 40809 8480 40815 8856
rect 40655 8468 40815 8480
rect 41027 8856 41187 8868
rect 41027 8480 41033 8856
rect 41067 8480 41147 8856
rect 41181 8480 41187 8856
rect 41027 8468 41187 8480
rect 41399 8856 41559 8868
rect 41399 8480 41405 8856
rect 41439 8480 41519 8856
rect 41553 8480 41559 8856
rect 41399 8468 41559 8480
rect 41771 8856 41931 8868
rect 41771 8480 41777 8856
rect 41811 8480 41891 8856
rect 41925 8480 41931 8856
rect 41771 8468 41931 8480
rect 42143 8856 42303 8868
rect 42143 8480 42149 8856
rect 42183 8480 42263 8856
rect 42297 8480 42303 8856
rect 42143 8468 42303 8480
rect 42515 8856 42675 8868
rect 42515 8480 42521 8856
rect 42555 8480 42635 8856
rect 42669 8480 42675 8856
rect 42515 8468 42675 8480
rect 42887 8856 43047 8868
rect 42887 8480 42893 8856
rect 42927 8480 43007 8856
rect 43041 8480 43047 8856
rect 42887 8468 43047 8480
rect 43259 8856 43419 8868
rect 43259 8480 43265 8856
rect 43299 8480 43379 8856
rect 43413 8480 43419 8856
rect 43259 8468 43419 8480
rect 43631 8856 43791 8868
rect 43631 8480 43637 8856
rect 43671 8480 43751 8856
rect 43785 8480 43791 8856
rect 43631 8468 43791 8480
rect 44003 8856 44163 8868
rect 44003 8480 44009 8856
rect 44043 8480 44123 8856
rect 44157 8480 44163 8856
rect 44003 8468 44163 8480
rect 44375 8856 44535 8868
rect 44375 8480 44381 8856
rect 44415 8480 44495 8856
rect 44529 8480 44535 8856
rect 44375 8468 44535 8480
rect 44747 8856 44907 8868
rect 44747 8480 44753 8856
rect 44787 8480 44867 8856
rect 44901 8480 44907 8856
rect 44747 8468 44907 8480
rect 45118 8856 45170 8902
rect 45118 8480 45125 8856
rect 45159 8480 45170 8856
rect 39280 8427 39368 8428
rect 39280 8422 39529 8427
rect 39280 8278 39348 8422
rect 39518 8381 39529 8422
rect 39518 8319 39528 8381
rect 39518 8278 39529 8319
rect 39280 8273 39529 8278
rect 39280 8272 39366 8273
rect 39280 8220 39328 8272
rect 39584 8232 39654 8468
rect 39709 8422 39901 8427
rect 39709 8381 39720 8422
rect 39710 8319 39720 8381
rect 39709 8278 39720 8319
rect 39890 8381 39901 8422
rect 39890 8319 39900 8381
rect 39890 8278 39901 8319
rect 39709 8273 39901 8278
rect 39956 8232 40026 8468
rect 40081 8422 40273 8427
rect 40081 8381 40092 8422
rect 40082 8319 40092 8381
rect 40081 8278 40092 8319
rect 40262 8381 40273 8422
rect 40262 8319 40272 8381
rect 40262 8278 40273 8319
rect 40081 8273 40273 8278
rect 40328 8232 40398 8468
rect 40453 8426 40645 8427
rect 40700 8426 40770 8468
rect 40825 8426 41017 8427
rect 40453 8422 41017 8426
rect 40453 8381 40464 8422
rect 40454 8319 40464 8381
rect 40453 8278 40464 8319
rect 40634 8278 40836 8422
rect 41006 8381 41017 8422
rect 41006 8319 41016 8381
rect 41006 8278 41017 8319
rect 40453 8274 41017 8278
rect 40453 8273 40645 8274
rect 40700 8232 40770 8274
rect 40825 8273 41017 8274
rect 41072 8232 41142 8468
rect 41197 8422 41389 8427
rect 41197 8381 41208 8422
rect 41198 8319 41208 8381
rect 41197 8278 41208 8319
rect 41378 8381 41389 8422
rect 41378 8319 41388 8381
rect 41378 8278 41389 8319
rect 41197 8273 41389 8278
rect 41444 8232 41514 8468
rect 41569 8422 41761 8427
rect 41569 8381 41580 8422
rect 41570 8319 41580 8381
rect 41569 8278 41580 8319
rect 41750 8381 41761 8422
rect 41750 8319 41760 8381
rect 41750 8278 41761 8319
rect 41569 8273 41761 8278
rect 41816 8232 41886 8468
rect 42188 8428 42258 8468
rect 41996 8427 42414 8428
rect 41941 8422 42505 8427
rect 41941 8381 41952 8422
rect 41942 8319 41952 8381
rect 41941 8278 41952 8319
rect 42122 8278 42324 8422
rect 42494 8381 42505 8422
rect 42494 8319 42504 8381
rect 42494 8278 42505 8319
rect 41941 8273 42505 8278
rect 41996 8272 42414 8273
rect 42188 8232 42258 8272
rect 42560 8232 42630 8468
rect 42685 8422 42877 8427
rect 42685 8381 42696 8422
rect 42686 8319 42696 8381
rect 42685 8278 42696 8319
rect 42866 8381 42877 8422
rect 42866 8319 42876 8381
rect 42866 8278 42877 8319
rect 42685 8273 42877 8278
rect 42932 8232 43002 8468
rect 43057 8422 43249 8427
rect 43057 8381 43068 8422
rect 43058 8319 43068 8381
rect 43057 8278 43068 8319
rect 43238 8381 43249 8422
rect 43238 8319 43248 8381
rect 43238 8278 43249 8319
rect 43057 8273 43249 8278
rect 43304 8232 43374 8468
rect 43676 8428 43746 8468
rect 43524 8427 43900 8428
rect 43429 8422 43993 8427
rect 43429 8381 43440 8422
rect 43430 8319 43440 8381
rect 43429 8278 43440 8319
rect 43610 8278 43812 8422
rect 43982 8381 43993 8422
rect 43982 8319 43992 8381
rect 43982 8278 43993 8319
rect 43429 8273 43993 8278
rect 43524 8272 43900 8273
rect 43676 8232 43746 8272
rect 44048 8232 44118 8468
rect 44173 8422 44365 8427
rect 44173 8381 44184 8422
rect 44174 8319 44184 8381
rect 44173 8278 44184 8319
rect 44354 8381 44365 8422
rect 44354 8319 44364 8381
rect 44354 8278 44365 8319
rect 44173 8273 44365 8278
rect 44420 8232 44490 8468
rect 44545 8422 44737 8427
rect 44545 8381 44556 8422
rect 44546 8319 44556 8381
rect 44545 8278 44556 8319
rect 44726 8381 44737 8422
rect 44726 8319 44736 8381
rect 44726 8278 44737 8319
rect 44545 8273 44737 8278
rect 44792 8232 44862 8468
rect 45118 8428 45170 8480
rect 45012 8427 45170 8428
rect 44917 8422 45170 8427
rect 44917 8381 44928 8422
rect 44918 8319 44928 8381
rect 44917 8278 44928 8319
rect 45098 8278 45170 8422
rect 44917 8273 45170 8278
rect 45012 8272 45170 8273
rect 39280 7844 39287 8220
rect 39321 7844 39328 8220
rect 39280 7792 39328 7844
rect 39539 8220 39699 8232
rect 39539 7844 39545 8220
rect 39579 7844 39659 8220
rect 39693 7844 39699 8220
rect 39539 7832 39699 7844
rect 39911 8220 40071 8232
rect 39911 7844 39917 8220
rect 39951 7844 40031 8220
rect 40065 7844 40071 8220
rect 39911 7832 40071 7844
rect 40283 8220 40443 8232
rect 40283 7844 40289 8220
rect 40323 7844 40403 8220
rect 40437 7844 40443 8220
rect 40283 7832 40443 7844
rect 40655 8220 40815 8232
rect 40655 7844 40661 8220
rect 40695 7844 40775 8220
rect 40809 7844 40815 8220
rect 40655 7832 40815 7844
rect 41027 8220 41187 8232
rect 41027 7844 41033 8220
rect 41067 7844 41147 8220
rect 41181 7844 41187 8220
rect 41027 7832 41187 7844
rect 41399 8220 41559 8232
rect 41399 7844 41405 8220
rect 41439 7844 41519 8220
rect 41553 7844 41559 8220
rect 41399 7832 41559 7844
rect 41771 8220 41931 8232
rect 41771 7844 41777 8220
rect 41811 7844 41891 8220
rect 41925 7844 41931 8220
rect 41771 7832 41931 7844
rect 42143 8220 42303 8232
rect 42143 7844 42149 8220
rect 42183 7844 42263 8220
rect 42297 7844 42303 8220
rect 42143 7832 42303 7844
rect 42515 8220 42675 8232
rect 42515 7844 42521 8220
rect 42555 7844 42635 8220
rect 42669 7844 42675 8220
rect 42515 7832 42675 7844
rect 42887 8220 43047 8232
rect 42887 7844 42893 8220
rect 42927 7844 43007 8220
rect 43041 7844 43047 8220
rect 42887 7832 43047 7844
rect 43259 8220 43419 8232
rect 43259 7844 43265 8220
rect 43299 7844 43379 8220
rect 43413 7844 43419 8220
rect 43259 7832 43419 7844
rect 43631 8220 43791 8232
rect 43631 7844 43637 8220
rect 43671 7844 43751 8220
rect 43785 7844 43791 8220
rect 43631 7832 43791 7844
rect 44003 8220 44163 8232
rect 44003 7844 44009 8220
rect 44043 7844 44123 8220
rect 44157 7844 44163 8220
rect 44003 7832 44163 7844
rect 44375 8220 44535 8232
rect 44375 7844 44381 8220
rect 44415 7844 44495 8220
rect 44529 7844 44535 8220
rect 44375 7832 44535 7844
rect 44747 8220 44907 8232
rect 44747 7844 44753 8220
rect 44787 7844 44867 8220
rect 44901 7844 44907 8220
rect 44747 7832 44907 7844
rect 45118 8220 45170 8272
rect 45118 7844 45125 8220
rect 45159 7844 45170 8220
rect 39280 7791 39370 7792
rect 39280 7786 39529 7791
rect 39280 7642 39348 7786
rect 39518 7745 39529 7786
rect 39518 7683 39528 7745
rect 39518 7642 39529 7683
rect 39280 7637 39529 7642
rect 39280 7632 39370 7637
rect 39280 7584 39328 7632
rect 39584 7596 39654 7832
rect 39709 7786 39901 7791
rect 39709 7745 39720 7786
rect 39710 7683 39720 7745
rect 39709 7642 39720 7683
rect 39890 7745 39901 7786
rect 39890 7683 39900 7745
rect 39890 7642 39901 7683
rect 39709 7637 39901 7642
rect 39956 7596 40026 7832
rect 40081 7786 40273 7791
rect 40081 7745 40092 7786
rect 40082 7683 40092 7745
rect 40081 7642 40092 7683
rect 40262 7745 40273 7786
rect 40262 7683 40272 7745
rect 40262 7642 40273 7683
rect 40081 7637 40273 7642
rect 40328 7596 40398 7832
rect 40453 7788 40645 7791
rect 40700 7788 40770 7832
rect 40825 7788 41017 7791
rect 40453 7786 41017 7788
rect 40453 7745 40464 7786
rect 40454 7683 40464 7745
rect 40453 7642 40464 7683
rect 40634 7642 40836 7786
rect 41006 7745 41017 7786
rect 41006 7683 41016 7745
rect 41006 7642 41017 7683
rect 40453 7637 41017 7642
rect 40494 7636 40970 7637
rect 40700 7596 40770 7636
rect 41072 7596 41142 7832
rect 41197 7786 41389 7791
rect 41197 7745 41208 7786
rect 41198 7683 41208 7745
rect 41197 7642 41208 7683
rect 41378 7745 41389 7786
rect 41378 7683 41388 7745
rect 41378 7642 41389 7683
rect 41197 7637 41389 7642
rect 41444 7596 41514 7832
rect 41569 7786 41761 7791
rect 41569 7745 41580 7786
rect 41570 7683 41580 7745
rect 41569 7642 41580 7683
rect 41750 7745 41761 7786
rect 41750 7683 41760 7745
rect 41750 7642 41761 7683
rect 41569 7637 41761 7642
rect 41816 7596 41886 7832
rect 42188 7792 42258 7832
rect 42016 7791 42434 7792
rect 41941 7786 42505 7791
rect 41941 7745 41952 7786
rect 41942 7683 41952 7745
rect 41941 7642 41952 7683
rect 42122 7642 42324 7786
rect 42494 7745 42505 7786
rect 42494 7683 42504 7745
rect 42494 7642 42505 7683
rect 41941 7637 42505 7642
rect 42016 7636 42434 7637
rect 42188 7596 42258 7636
rect 42560 7596 42630 7832
rect 42685 7786 42877 7791
rect 42685 7745 42696 7786
rect 42686 7683 42696 7745
rect 42685 7642 42696 7683
rect 42866 7745 42877 7786
rect 42866 7683 42876 7745
rect 42866 7642 42877 7683
rect 42685 7637 42877 7642
rect 42932 7596 43002 7832
rect 43057 7786 43249 7791
rect 43057 7745 43068 7786
rect 43058 7683 43068 7745
rect 43057 7642 43068 7683
rect 43238 7745 43249 7786
rect 43238 7683 43248 7745
rect 43238 7642 43249 7683
rect 43057 7637 43249 7642
rect 43304 7596 43374 7832
rect 43676 7792 43746 7832
rect 43512 7791 43888 7792
rect 43429 7786 43993 7791
rect 43429 7745 43440 7786
rect 43430 7683 43440 7745
rect 43429 7642 43440 7683
rect 43610 7642 43812 7786
rect 43982 7745 43993 7786
rect 43982 7683 43992 7745
rect 43982 7642 43993 7683
rect 43429 7637 43993 7642
rect 43512 7636 43888 7637
rect 43676 7596 43746 7636
rect 44048 7596 44118 7832
rect 44173 7786 44365 7791
rect 44173 7745 44184 7786
rect 44174 7683 44184 7745
rect 44173 7642 44184 7683
rect 44354 7745 44365 7786
rect 44354 7683 44364 7745
rect 44354 7642 44365 7683
rect 44173 7637 44365 7642
rect 44420 7596 44490 7832
rect 44545 7786 44737 7791
rect 44545 7745 44556 7786
rect 44546 7683 44556 7745
rect 44545 7642 44556 7683
rect 44726 7745 44737 7786
rect 44726 7683 44736 7745
rect 44726 7642 44737 7683
rect 44545 7637 44737 7642
rect 44792 7596 44862 7832
rect 45118 7792 45170 7844
rect 45028 7791 45170 7792
rect 44917 7786 45170 7791
rect 44917 7745 44928 7786
rect 44918 7683 44928 7745
rect 44917 7642 44928 7683
rect 45098 7642 45170 7786
rect 44917 7637 45170 7642
rect 45028 7636 45170 7637
rect 39280 7208 39287 7584
rect 39321 7208 39328 7584
rect 39280 7162 39328 7208
rect 39539 7584 39699 7596
rect 39539 7208 39545 7584
rect 39579 7208 39659 7584
rect 39693 7208 39699 7584
rect 39539 7196 39699 7208
rect 39911 7584 40071 7596
rect 39911 7208 39917 7584
rect 39951 7208 40031 7584
rect 40065 7208 40071 7584
rect 39911 7196 40071 7208
rect 40283 7584 40443 7596
rect 40283 7208 40289 7584
rect 40323 7208 40403 7584
rect 40437 7208 40443 7584
rect 40283 7196 40443 7208
rect 40655 7584 40815 7596
rect 40655 7208 40661 7584
rect 40695 7208 40775 7584
rect 40809 7208 40815 7584
rect 40655 7196 40815 7208
rect 41027 7584 41187 7596
rect 41027 7208 41033 7584
rect 41067 7208 41147 7584
rect 41181 7208 41187 7584
rect 41027 7196 41187 7208
rect 41399 7584 41559 7596
rect 41399 7208 41405 7584
rect 41439 7208 41519 7584
rect 41553 7208 41559 7584
rect 41399 7196 41559 7208
rect 41771 7584 41931 7596
rect 41771 7208 41777 7584
rect 41811 7208 41891 7584
rect 41925 7208 41931 7584
rect 41771 7196 41931 7208
rect 42143 7584 42303 7596
rect 42143 7208 42149 7584
rect 42183 7208 42263 7584
rect 42297 7208 42303 7584
rect 42143 7196 42303 7208
rect 42515 7584 42675 7596
rect 42515 7208 42521 7584
rect 42555 7208 42635 7584
rect 42669 7208 42675 7584
rect 42515 7196 42675 7208
rect 42887 7584 43047 7596
rect 42887 7208 42893 7584
rect 42927 7208 43007 7584
rect 43041 7208 43047 7584
rect 42887 7196 43047 7208
rect 43259 7584 43419 7596
rect 43259 7208 43265 7584
rect 43299 7208 43379 7584
rect 43413 7208 43419 7584
rect 43259 7196 43419 7208
rect 43631 7584 43791 7596
rect 43631 7208 43637 7584
rect 43671 7208 43751 7584
rect 43785 7208 43791 7584
rect 43631 7196 43791 7208
rect 44003 7584 44163 7596
rect 44003 7208 44009 7584
rect 44043 7208 44123 7584
rect 44157 7208 44163 7584
rect 44003 7196 44163 7208
rect 44375 7584 44535 7596
rect 44375 7208 44381 7584
rect 44415 7208 44495 7584
rect 44529 7208 44535 7584
rect 44375 7196 44535 7208
rect 44747 7584 44907 7596
rect 44747 7208 44753 7584
rect 44787 7208 44867 7584
rect 44901 7208 44907 7584
rect 44747 7196 44907 7208
rect 45118 7584 45170 7636
rect 45118 7208 45125 7584
rect 45159 7208 45170 7584
rect 39280 7102 39348 7162
rect 39518 7155 39528 7162
rect 39710 7155 39720 7162
rect 39518 7109 39529 7155
rect 39709 7109 39720 7155
rect 39890 7155 39900 7162
rect 39518 7102 39528 7109
rect 39710 7102 39720 7109
rect 39890 7109 39901 7155
rect 39890 7102 39900 7109
rect 39962 6854 40020 7196
rect 40706 7162 40764 7196
rect 40082 7155 40092 7162
rect 40081 7109 40092 7155
rect 40262 7155 40272 7162
rect 40454 7155 40464 7162
rect 40082 7102 40092 7109
rect 40262 7109 40273 7155
rect 40453 7109 40464 7155
rect 40262 7102 40272 7109
rect 40454 7102 40464 7109
rect 40634 7102 40836 7162
rect 41006 7155 41016 7162
rect 41198 7155 41208 7162
rect 41006 7109 41017 7155
rect 41197 7109 41208 7155
rect 41378 7155 41388 7162
rect 41006 7102 41016 7109
rect 41198 7102 41208 7109
rect 41378 7109 41389 7155
rect 41378 7102 41388 7109
rect 40580 7100 40910 7102
rect 41450 6854 41508 7196
rect 42194 7162 42252 7196
rect 41570 7155 41580 7162
rect 41569 7109 41580 7155
rect 41750 7155 41760 7162
rect 41942 7155 41952 7162
rect 41570 7102 41580 7109
rect 41750 7109 41761 7155
rect 41941 7109 41952 7155
rect 41750 7102 41760 7109
rect 41942 7102 41952 7109
rect 42122 7102 42324 7162
rect 42494 7155 42504 7162
rect 42686 7155 42696 7162
rect 42494 7109 42505 7155
rect 42685 7109 42696 7155
rect 42866 7155 42876 7162
rect 42494 7102 42504 7109
rect 42686 7102 42696 7109
rect 42866 7109 42877 7155
rect 42866 7102 42876 7109
rect 42938 6854 42996 7196
rect 43682 7162 43740 7196
rect 43058 7155 43068 7162
rect 43057 7109 43068 7155
rect 43238 7155 43248 7162
rect 43430 7155 43440 7162
rect 43058 7102 43068 7109
rect 43238 7109 43249 7155
rect 43429 7109 43440 7155
rect 43238 7102 43248 7109
rect 43430 7102 43440 7109
rect 43610 7102 43812 7162
rect 43982 7155 43992 7162
rect 44174 7155 44184 7162
rect 43982 7109 43993 7155
rect 44173 7109 44184 7155
rect 44354 7155 44364 7162
rect 43982 7102 43992 7109
rect 44174 7102 44184 7109
rect 44354 7109 44365 7155
rect 44354 7102 44364 7109
rect 44426 6854 44484 7196
rect 45118 7162 45170 7208
rect 45208 8868 45260 8992
rect 45294 8902 45300 8962
rect 45470 8955 45480 8962
rect 45662 8955 45672 8962
rect 45470 8909 45481 8955
rect 45661 8909 45672 8955
rect 45842 8955 45852 8962
rect 45470 8902 45480 8909
rect 45662 8902 45672 8909
rect 45842 8909 45853 8955
rect 45842 8902 45852 8909
rect 45914 8868 45972 8992
rect 46034 8955 46044 8962
rect 46033 8909 46044 8955
rect 46214 8955 46224 8962
rect 46406 8955 46416 8962
rect 46034 8902 46044 8909
rect 46214 8909 46225 8955
rect 46405 8909 46416 8955
rect 46586 8955 46596 8962
rect 46214 8902 46224 8909
rect 46406 8902 46416 8909
rect 46586 8909 46597 8955
rect 46586 8902 46596 8909
rect 46658 8868 46716 8992
rect 46778 8955 46788 8962
rect 46777 8909 46788 8955
rect 46958 8955 46968 8962
rect 47150 8955 47160 8962
rect 46778 8902 46788 8909
rect 46958 8909 46969 8955
rect 47149 8909 47160 8955
rect 47330 8955 47340 8962
rect 46958 8902 46968 8909
rect 47150 8902 47160 8909
rect 47330 8909 47341 8955
rect 47330 8902 47340 8909
rect 47402 8868 47460 8992
rect 47522 8955 47532 8962
rect 47521 8909 47532 8955
rect 47702 8955 47712 8962
rect 47894 8955 47904 8962
rect 47522 8902 47532 8909
rect 47702 8909 47713 8955
rect 47893 8909 47904 8955
rect 48074 8955 48084 8962
rect 47702 8902 47712 8909
rect 47894 8902 47904 8909
rect 48074 8909 48085 8955
rect 48074 8902 48084 8909
rect 48146 8868 48204 8992
rect 48266 8955 48276 8962
rect 48265 8909 48276 8955
rect 48446 8955 48456 8962
rect 48638 8955 48648 8962
rect 48266 8902 48276 8909
rect 48446 8909 48457 8955
rect 48637 8909 48648 8955
rect 48818 8955 48828 8962
rect 48446 8902 48456 8909
rect 48638 8902 48648 8909
rect 48818 8909 48829 8955
rect 48818 8902 48828 8909
rect 48890 8868 48948 8992
rect 49010 8955 49020 8962
rect 49009 8909 49020 8955
rect 49190 8955 49200 8962
rect 49382 8955 49392 8962
rect 49010 8902 49020 8909
rect 49190 8909 49201 8955
rect 49381 8909 49392 8955
rect 49562 8955 49572 8962
rect 49190 8902 49200 8909
rect 49382 8902 49392 8909
rect 49562 8909 49573 8955
rect 49562 8902 49572 8909
rect 49634 8868 49692 8992
rect 49754 8955 49764 8962
rect 49753 8909 49764 8955
rect 49934 8955 49944 8962
rect 50126 8955 50136 8962
rect 49754 8902 49764 8909
rect 49934 8909 49945 8955
rect 50125 8909 50136 8955
rect 50306 8955 50316 8962
rect 49934 8902 49944 8909
rect 50126 8902 50136 8909
rect 50306 8909 50317 8955
rect 50306 8902 50316 8909
rect 50378 8868 50436 8992
rect 50498 8955 50508 8962
rect 50497 8909 50508 8955
rect 50678 8955 50688 8962
rect 50870 8955 50880 8962
rect 50498 8902 50508 8909
rect 50678 8909 50689 8955
rect 50869 8909 50880 8955
rect 51050 8955 51060 8962
rect 50678 8902 50688 8909
rect 50870 8902 50880 8909
rect 51050 8909 51061 8955
rect 51050 8902 51060 8909
rect 51104 8868 51162 8992
rect 45208 8856 45279 8868
rect 45208 8480 45239 8856
rect 45273 8480 45279 8856
rect 45208 8468 45279 8480
rect 45491 8856 45651 8868
rect 45491 8480 45497 8856
rect 45531 8480 45611 8856
rect 45645 8480 45651 8856
rect 45491 8468 45651 8480
rect 45863 8856 46023 8868
rect 45863 8480 45869 8856
rect 45903 8480 45983 8856
rect 46017 8480 46023 8856
rect 45863 8468 46023 8480
rect 46235 8856 46395 8868
rect 46235 8480 46241 8856
rect 46275 8480 46355 8856
rect 46389 8480 46395 8856
rect 46235 8468 46395 8480
rect 46607 8856 46767 8868
rect 46607 8480 46613 8856
rect 46647 8480 46727 8856
rect 46761 8480 46767 8856
rect 46607 8468 46767 8480
rect 46979 8856 47139 8868
rect 46979 8480 46985 8856
rect 47019 8480 47099 8856
rect 47133 8480 47139 8856
rect 46979 8468 47139 8480
rect 47351 8856 47511 8868
rect 47351 8480 47357 8856
rect 47391 8480 47471 8856
rect 47505 8480 47511 8856
rect 47351 8468 47511 8480
rect 47723 8856 47883 8868
rect 47723 8480 47729 8856
rect 47763 8480 47843 8856
rect 47877 8480 47883 8856
rect 47723 8468 47883 8480
rect 48095 8856 48255 8868
rect 48095 8480 48101 8856
rect 48135 8480 48215 8856
rect 48249 8480 48255 8856
rect 48095 8468 48255 8480
rect 48467 8856 48627 8868
rect 48467 8480 48473 8856
rect 48507 8480 48587 8856
rect 48621 8480 48627 8856
rect 48467 8468 48627 8480
rect 48839 8856 48999 8868
rect 48839 8480 48845 8856
rect 48879 8480 48959 8856
rect 48993 8480 48999 8856
rect 48839 8468 48999 8480
rect 49211 8856 49371 8868
rect 49211 8480 49217 8856
rect 49251 8480 49331 8856
rect 49365 8480 49371 8856
rect 49211 8468 49371 8480
rect 49583 8856 49743 8868
rect 49583 8480 49589 8856
rect 49623 8480 49703 8856
rect 49737 8480 49743 8856
rect 49583 8468 49743 8480
rect 49955 8856 50115 8868
rect 49955 8480 49961 8856
rect 49995 8480 50075 8856
rect 50109 8480 50115 8856
rect 49955 8468 50115 8480
rect 50327 8856 50487 8868
rect 50327 8480 50333 8856
rect 50367 8480 50447 8856
rect 50481 8480 50487 8856
rect 50327 8468 50487 8480
rect 50699 8856 50859 8868
rect 50699 8480 50705 8856
rect 50739 8480 50819 8856
rect 50853 8480 50859 8856
rect 50699 8468 50859 8480
rect 51071 8856 51162 8868
rect 51071 8480 51077 8856
rect 51111 8480 51162 8856
rect 51071 8468 51162 8480
rect 45208 8232 45260 8468
rect 45288 8427 45414 8428
rect 45288 8422 45481 8427
rect 45288 8278 45300 8422
rect 45470 8381 45481 8422
rect 45470 8319 45480 8381
rect 45470 8278 45481 8319
rect 45288 8273 45481 8278
rect 45288 8272 45414 8273
rect 45536 8232 45606 8468
rect 45661 8422 45853 8427
rect 45661 8381 45672 8422
rect 45662 8319 45672 8381
rect 45661 8278 45672 8319
rect 45842 8381 45853 8422
rect 45842 8319 45852 8381
rect 45842 8278 45853 8319
rect 45661 8273 45853 8278
rect 45908 8232 45978 8468
rect 46033 8422 46225 8427
rect 46033 8381 46044 8422
rect 46034 8319 46044 8381
rect 46033 8278 46044 8319
rect 46214 8381 46225 8422
rect 46214 8319 46224 8381
rect 46214 8278 46225 8319
rect 46033 8273 46225 8278
rect 46280 8232 46350 8468
rect 46405 8422 46597 8427
rect 46405 8381 46416 8422
rect 46406 8319 46416 8381
rect 46405 8278 46416 8319
rect 46586 8381 46597 8422
rect 46586 8319 46596 8381
rect 46586 8278 46597 8319
rect 46405 8273 46597 8278
rect 46652 8232 46722 8468
rect 46777 8422 46969 8427
rect 46777 8381 46788 8422
rect 46778 8319 46788 8381
rect 46777 8278 46788 8319
rect 46958 8381 46969 8422
rect 46958 8319 46968 8381
rect 46958 8278 46969 8319
rect 46777 8273 46969 8278
rect 47024 8232 47094 8468
rect 47149 8422 47341 8427
rect 47149 8381 47160 8422
rect 47150 8319 47160 8381
rect 47149 8278 47160 8319
rect 47330 8381 47341 8422
rect 47330 8319 47340 8381
rect 47330 8278 47341 8319
rect 47149 8273 47341 8278
rect 47396 8232 47466 8468
rect 47521 8422 47713 8427
rect 47521 8381 47532 8422
rect 47522 8319 47532 8381
rect 47521 8278 47532 8319
rect 47702 8381 47713 8422
rect 47702 8319 47712 8381
rect 47702 8278 47713 8319
rect 47521 8273 47713 8278
rect 47768 8232 47838 8468
rect 47893 8422 48085 8427
rect 47893 8381 47904 8422
rect 47894 8319 47904 8381
rect 47893 8278 47904 8319
rect 48074 8381 48085 8422
rect 48074 8319 48084 8381
rect 48074 8278 48085 8319
rect 47893 8273 48085 8278
rect 48140 8232 48210 8468
rect 48265 8422 48457 8427
rect 48265 8381 48276 8422
rect 48266 8319 48276 8381
rect 48265 8278 48276 8319
rect 48446 8381 48457 8422
rect 48446 8319 48456 8381
rect 48446 8278 48457 8319
rect 48265 8273 48457 8278
rect 48512 8232 48582 8468
rect 48637 8422 48829 8427
rect 48637 8381 48648 8422
rect 48638 8319 48648 8381
rect 48637 8278 48648 8319
rect 48818 8381 48829 8422
rect 48818 8319 48828 8381
rect 48818 8278 48829 8319
rect 48637 8273 48829 8278
rect 48884 8232 48954 8468
rect 49009 8422 49201 8427
rect 49009 8381 49020 8422
rect 49010 8319 49020 8381
rect 49009 8278 49020 8319
rect 49190 8381 49201 8422
rect 49190 8319 49200 8381
rect 49190 8278 49201 8319
rect 49009 8273 49201 8278
rect 49256 8232 49326 8468
rect 49381 8422 49573 8427
rect 49381 8381 49392 8422
rect 49382 8319 49392 8381
rect 49381 8278 49392 8319
rect 49562 8381 49573 8422
rect 49562 8319 49572 8381
rect 49562 8278 49573 8319
rect 49381 8273 49573 8278
rect 49628 8232 49698 8468
rect 49753 8422 49945 8427
rect 49753 8381 49764 8422
rect 49754 8319 49764 8381
rect 49753 8278 49764 8319
rect 49934 8381 49945 8422
rect 49934 8319 49944 8381
rect 49934 8278 49945 8319
rect 49753 8273 49945 8278
rect 50000 8232 50070 8468
rect 50125 8422 50317 8427
rect 50125 8381 50136 8422
rect 50126 8319 50136 8381
rect 50125 8278 50136 8319
rect 50306 8381 50317 8422
rect 50306 8319 50316 8381
rect 50306 8278 50317 8319
rect 50125 8273 50317 8278
rect 50372 8232 50442 8468
rect 50497 8422 50689 8427
rect 50497 8381 50508 8422
rect 50498 8319 50508 8381
rect 50497 8278 50508 8319
rect 50678 8381 50689 8422
rect 50678 8319 50688 8381
rect 50678 8278 50689 8319
rect 50497 8273 50689 8278
rect 50744 8232 50814 8468
rect 50869 8422 51061 8427
rect 50869 8381 50880 8422
rect 50870 8319 50880 8381
rect 50869 8278 50880 8319
rect 51050 8381 51061 8422
rect 51050 8319 51060 8381
rect 51050 8278 51061 8319
rect 50869 8273 51061 8278
rect 51104 8232 51162 8468
rect 45208 8220 45279 8232
rect 45208 7844 45239 8220
rect 45273 7844 45279 8220
rect 45208 7832 45279 7844
rect 45491 8220 45651 8232
rect 45491 7844 45497 8220
rect 45531 7844 45611 8220
rect 45645 7844 45651 8220
rect 45491 7832 45651 7844
rect 45863 8220 46023 8232
rect 45863 7844 45869 8220
rect 45903 7844 45983 8220
rect 46017 7844 46023 8220
rect 45863 7832 46023 7844
rect 46235 8220 46395 8232
rect 46235 7844 46241 8220
rect 46275 7844 46355 8220
rect 46389 7844 46395 8220
rect 46235 7832 46395 7844
rect 46607 8220 46767 8232
rect 46607 7844 46613 8220
rect 46647 7844 46727 8220
rect 46761 7844 46767 8220
rect 46607 7832 46767 7844
rect 46979 8220 47139 8232
rect 46979 7844 46985 8220
rect 47019 7844 47099 8220
rect 47133 7844 47139 8220
rect 46979 7832 47139 7844
rect 47351 8220 47511 8232
rect 47351 7844 47357 8220
rect 47391 7844 47471 8220
rect 47505 7844 47511 8220
rect 47351 7832 47511 7844
rect 47723 8220 47883 8232
rect 47723 7844 47729 8220
rect 47763 7844 47843 8220
rect 47877 7844 47883 8220
rect 47723 7832 47883 7844
rect 48095 8220 48255 8232
rect 48095 7844 48101 8220
rect 48135 7844 48215 8220
rect 48249 7844 48255 8220
rect 48095 7832 48255 7844
rect 48467 8220 48627 8232
rect 48467 7844 48473 8220
rect 48507 7844 48587 8220
rect 48621 7844 48627 8220
rect 48467 7832 48627 7844
rect 48839 8220 48999 8232
rect 48839 7844 48845 8220
rect 48879 7844 48959 8220
rect 48993 7844 48999 8220
rect 48839 7832 48999 7844
rect 49211 8220 49371 8232
rect 49211 7844 49217 8220
rect 49251 7844 49331 8220
rect 49365 7844 49371 8220
rect 49211 7832 49371 7844
rect 49583 8220 49743 8232
rect 49583 7844 49589 8220
rect 49623 7844 49703 8220
rect 49737 7844 49743 8220
rect 49583 7832 49743 7844
rect 49955 8220 50115 8232
rect 49955 7844 49961 8220
rect 49995 7844 50075 8220
rect 50109 7844 50115 8220
rect 49955 7832 50115 7844
rect 50327 8220 50487 8232
rect 50327 7844 50333 8220
rect 50367 7844 50447 8220
rect 50481 7844 50487 8220
rect 50327 7832 50487 7844
rect 50699 8220 50859 8232
rect 50699 7844 50705 8220
rect 50739 7844 50819 8220
rect 50853 7844 50859 8220
rect 50699 7832 50859 7844
rect 51071 8220 51162 8232
rect 51071 7844 51077 8220
rect 51111 7844 51162 8220
rect 51071 7832 51162 7844
rect 45208 7596 45260 7832
rect 45288 7791 45430 7792
rect 45288 7786 45481 7791
rect 45288 7642 45300 7786
rect 45470 7745 45481 7786
rect 45470 7683 45480 7745
rect 45470 7642 45481 7683
rect 45288 7637 45481 7642
rect 45288 7636 45430 7637
rect 45536 7596 45606 7832
rect 45661 7786 45853 7791
rect 45661 7745 45672 7786
rect 45662 7683 45672 7745
rect 45661 7642 45672 7683
rect 45842 7745 45853 7786
rect 45842 7683 45852 7745
rect 45842 7642 45853 7683
rect 45661 7637 45853 7642
rect 45908 7596 45978 7832
rect 46033 7786 46225 7791
rect 46033 7745 46044 7786
rect 46034 7683 46044 7745
rect 46033 7642 46044 7683
rect 46214 7745 46225 7786
rect 46214 7683 46224 7745
rect 46214 7642 46225 7683
rect 46033 7637 46225 7642
rect 46280 7596 46350 7832
rect 46405 7786 46597 7791
rect 46405 7745 46416 7786
rect 46406 7683 46416 7745
rect 46405 7642 46416 7683
rect 46586 7745 46597 7786
rect 46586 7683 46596 7745
rect 46586 7642 46597 7683
rect 46405 7637 46597 7642
rect 46652 7596 46722 7832
rect 46777 7786 46969 7791
rect 46777 7745 46788 7786
rect 46778 7683 46788 7745
rect 46777 7642 46788 7683
rect 46958 7745 46969 7786
rect 46958 7683 46968 7745
rect 46958 7642 46969 7683
rect 46777 7637 46969 7642
rect 47024 7596 47094 7832
rect 47149 7786 47341 7791
rect 47149 7745 47160 7786
rect 47150 7683 47160 7745
rect 47149 7642 47160 7683
rect 47330 7745 47341 7786
rect 47330 7683 47340 7745
rect 47330 7642 47341 7683
rect 47149 7637 47341 7642
rect 47396 7596 47466 7832
rect 47521 7786 47713 7791
rect 47521 7745 47532 7786
rect 47522 7683 47532 7745
rect 47521 7642 47532 7683
rect 47702 7745 47713 7786
rect 47702 7683 47712 7745
rect 47702 7642 47713 7683
rect 47521 7637 47713 7642
rect 47768 7596 47838 7832
rect 47893 7786 48085 7791
rect 47893 7745 47904 7786
rect 47894 7683 47904 7745
rect 47893 7642 47904 7683
rect 48074 7745 48085 7786
rect 48074 7683 48084 7745
rect 48074 7642 48085 7683
rect 47893 7637 48085 7642
rect 48140 7596 48210 7832
rect 48265 7786 48457 7791
rect 48265 7745 48276 7786
rect 48266 7683 48276 7745
rect 48265 7642 48276 7683
rect 48446 7745 48457 7786
rect 48446 7683 48456 7745
rect 48446 7642 48457 7683
rect 48265 7637 48457 7642
rect 48512 7596 48582 7832
rect 48637 7786 48829 7791
rect 48637 7745 48648 7786
rect 48638 7683 48648 7745
rect 48637 7642 48648 7683
rect 48818 7745 48829 7786
rect 48818 7683 48828 7745
rect 48818 7642 48829 7683
rect 48637 7637 48829 7642
rect 48884 7596 48954 7832
rect 49009 7786 49201 7791
rect 49009 7745 49020 7786
rect 49010 7683 49020 7745
rect 49009 7642 49020 7683
rect 49190 7745 49201 7786
rect 49190 7683 49200 7745
rect 49190 7642 49201 7683
rect 49009 7637 49201 7642
rect 49256 7596 49326 7832
rect 49381 7786 49573 7791
rect 49381 7745 49392 7786
rect 49382 7683 49392 7745
rect 49381 7642 49392 7683
rect 49562 7745 49573 7786
rect 49562 7683 49572 7745
rect 49562 7642 49573 7683
rect 49381 7637 49573 7642
rect 49628 7596 49698 7832
rect 49753 7786 49945 7791
rect 49753 7745 49764 7786
rect 49754 7683 49764 7745
rect 49753 7642 49764 7683
rect 49934 7745 49945 7786
rect 49934 7683 49944 7745
rect 49934 7642 49945 7683
rect 49753 7637 49945 7642
rect 50000 7596 50070 7832
rect 50125 7786 50317 7791
rect 50125 7745 50136 7786
rect 50126 7683 50136 7745
rect 50125 7642 50136 7683
rect 50306 7745 50317 7786
rect 50306 7683 50316 7745
rect 50306 7642 50317 7683
rect 50125 7637 50317 7642
rect 50372 7596 50442 7832
rect 50497 7786 50689 7791
rect 50497 7745 50508 7786
rect 50498 7683 50508 7745
rect 50497 7642 50508 7683
rect 50678 7745 50689 7786
rect 50678 7683 50688 7745
rect 50678 7642 50689 7683
rect 50497 7637 50689 7642
rect 50744 7596 50814 7832
rect 50869 7786 51061 7791
rect 50869 7745 50880 7786
rect 50870 7683 50880 7745
rect 50869 7642 50880 7683
rect 51050 7745 51061 7786
rect 51050 7683 51060 7745
rect 51050 7642 51061 7683
rect 50869 7637 51061 7642
rect 51104 7596 51162 7832
rect 45208 7584 45279 7596
rect 45208 7208 45239 7584
rect 45273 7208 45279 7584
rect 45208 7196 45279 7208
rect 45491 7584 45651 7596
rect 45491 7208 45497 7584
rect 45531 7208 45611 7584
rect 45645 7208 45651 7584
rect 45491 7196 45651 7208
rect 45863 7584 46023 7596
rect 45863 7208 45869 7584
rect 45903 7208 45983 7584
rect 46017 7208 46023 7584
rect 45863 7196 46023 7208
rect 46235 7584 46395 7596
rect 46235 7208 46241 7584
rect 46275 7208 46355 7584
rect 46389 7208 46395 7584
rect 46235 7196 46395 7208
rect 46607 7584 46767 7596
rect 46607 7208 46613 7584
rect 46647 7208 46727 7584
rect 46761 7208 46767 7584
rect 46607 7196 46767 7208
rect 46979 7584 47139 7596
rect 46979 7208 46985 7584
rect 47019 7208 47099 7584
rect 47133 7208 47139 7584
rect 46979 7196 47139 7208
rect 47351 7584 47511 7596
rect 47351 7208 47357 7584
rect 47391 7208 47471 7584
rect 47505 7208 47511 7584
rect 47351 7196 47511 7208
rect 47723 7584 47883 7596
rect 47723 7208 47729 7584
rect 47763 7208 47843 7584
rect 47877 7208 47883 7584
rect 47723 7196 47883 7208
rect 48095 7584 48255 7596
rect 48095 7208 48101 7584
rect 48135 7208 48215 7584
rect 48249 7208 48255 7584
rect 48095 7196 48255 7208
rect 48467 7584 48627 7596
rect 48467 7208 48473 7584
rect 48507 7208 48587 7584
rect 48621 7208 48627 7584
rect 48467 7196 48627 7208
rect 48839 7584 48999 7596
rect 48839 7208 48845 7584
rect 48879 7208 48959 7584
rect 48993 7208 48999 7584
rect 48839 7196 48999 7208
rect 49211 7584 49371 7596
rect 49211 7208 49217 7584
rect 49251 7208 49331 7584
rect 49365 7208 49371 7584
rect 49211 7196 49371 7208
rect 49583 7584 49743 7596
rect 49583 7208 49589 7584
rect 49623 7208 49703 7584
rect 49737 7208 49743 7584
rect 49583 7196 49743 7208
rect 49955 7584 50115 7596
rect 49955 7208 49961 7584
rect 49995 7208 50075 7584
rect 50109 7208 50115 7584
rect 49955 7196 50115 7208
rect 50327 7584 50487 7596
rect 50327 7208 50333 7584
rect 50367 7208 50447 7584
rect 50481 7208 50487 7584
rect 50327 7196 50487 7208
rect 50699 7584 50859 7596
rect 50699 7208 50705 7584
rect 50739 7208 50819 7584
rect 50853 7208 50859 7584
rect 50699 7196 50859 7208
rect 51071 7584 51162 7596
rect 51071 7208 51077 7584
rect 51111 7208 51162 7584
rect 51071 7196 51162 7208
rect 44546 7155 44556 7162
rect 44545 7109 44556 7155
rect 44726 7155 44736 7162
rect 44918 7155 44928 7162
rect 44546 7102 44556 7109
rect 44726 7109 44737 7155
rect 44917 7109 44928 7155
rect 44726 7102 44736 7109
rect 44918 7102 44928 7109
rect 45098 7102 45170 7162
rect 45286 7102 45300 7162
rect 45470 7155 45480 7162
rect 45470 7109 45481 7155
rect 45470 7102 45480 7109
rect 39962 6790 44484 6854
rect 39504 6722 39576 6739
rect 38390 6697 39264 6698
rect 39504 6697 39521 6722
rect 38390 6381 39521 6697
rect 38390 6380 39264 6381
rect 39515 6325 39521 6381
rect 39559 6495 39576 6722
rect 39824 6722 39892 6739
rect 39559 6325 39565 6495
rect 39515 6313 39565 6325
rect 39824 6325 39839 6722
rect 39877 6647 39892 6722
rect 40722 6686 40776 6790
rect 41118 6686 41188 6790
rect 41450 6686 41508 6790
rect 41862 6686 41932 6790
rect 42194 6686 42252 6790
rect 42606 6686 42676 6790
rect 42938 6686 42996 6790
rect 43350 6686 43420 6790
rect 43670 6686 43724 6790
rect 40722 6680 40828 6686
rect 40112 6647 40122 6675
rect 39877 6441 40122 6647
rect 39877 6325 39892 6441
rect 40112 6401 40122 6441
rect 40404 6401 40414 6675
rect 40722 6610 40746 6680
rect 40816 6610 40828 6680
rect 40722 6604 40828 6610
rect 41106 6680 41200 6686
rect 41106 6610 41118 6680
rect 41188 6610 41200 6680
rect 41106 6604 41200 6610
rect 41450 6680 41572 6686
rect 41450 6610 41490 6680
rect 41560 6610 41572 6680
rect 41450 6604 41572 6610
rect 41850 6680 41944 6686
rect 41850 6610 41862 6680
rect 41932 6610 41944 6680
rect 41850 6604 41944 6610
rect 42194 6680 42316 6686
rect 42194 6610 42234 6680
rect 42304 6610 42316 6680
rect 42194 6604 42316 6610
rect 42594 6680 42688 6686
rect 42594 6610 42606 6680
rect 42676 6610 42688 6680
rect 42594 6604 42688 6610
rect 42938 6680 43060 6686
rect 42938 6610 42978 6680
rect 43048 6610 43060 6680
rect 42938 6604 43060 6610
rect 43338 6680 43432 6686
rect 43338 6610 43350 6680
rect 43420 6610 43432 6680
rect 43338 6604 43432 6610
rect 43600 6680 43724 6686
rect 43600 6610 43612 6680
rect 43682 6610 43724 6680
rect 43600 6604 43724 6610
rect 40722 6480 40776 6604
rect 40826 6567 40836 6576
rect 40825 6521 40836 6567
rect 41006 6567 41016 6576
rect 41198 6567 41208 6576
rect 40826 6512 40836 6521
rect 41006 6521 41017 6567
rect 41197 6521 41208 6567
rect 41378 6567 41388 6576
rect 41006 6512 41016 6521
rect 41198 6512 41208 6521
rect 41378 6521 41389 6567
rect 41378 6512 41388 6521
rect 41450 6480 41508 6604
rect 41570 6567 41580 6576
rect 41569 6521 41580 6567
rect 41750 6567 41760 6576
rect 41942 6567 41952 6576
rect 41570 6512 41580 6521
rect 41750 6521 41761 6567
rect 41941 6521 41952 6567
rect 42122 6567 42132 6576
rect 41750 6512 41760 6521
rect 41942 6512 41952 6521
rect 42122 6521 42133 6567
rect 42122 6512 42132 6521
rect 42194 6480 42252 6604
rect 42314 6567 42324 6576
rect 42313 6521 42324 6567
rect 42494 6567 42504 6576
rect 42686 6567 42696 6576
rect 42314 6512 42324 6521
rect 42494 6521 42505 6567
rect 42685 6521 42696 6567
rect 42866 6567 42876 6576
rect 42494 6512 42504 6521
rect 42686 6512 42696 6521
rect 42866 6521 42877 6567
rect 42866 6512 42876 6521
rect 42938 6480 42996 6604
rect 43058 6567 43068 6576
rect 43057 6521 43068 6567
rect 43238 6567 43248 6576
rect 43430 6567 43440 6576
rect 43058 6512 43068 6521
rect 43238 6521 43249 6567
rect 43429 6521 43440 6567
rect 43610 6567 43620 6576
rect 43238 6512 43248 6521
rect 43430 6512 43440 6521
rect 43610 6521 43621 6567
rect 43610 6512 43620 6521
rect 43670 6480 43724 6604
rect 44606 6557 44616 6831
rect 44898 6557 44908 6831
rect 45536 6794 45606 7196
rect 45662 7155 45672 7162
rect 45661 7109 45672 7155
rect 45842 7155 45852 7162
rect 46034 7155 46044 7162
rect 45662 7102 45672 7109
rect 45842 7109 45853 7155
rect 46033 7109 46044 7155
rect 46214 7155 46224 7162
rect 45842 7102 45852 7109
rect 46034 7102 46044 7109
rect 46214 7109 46225 7155
rect 46214 7102 46224 7109
rect 46280 6794 46350 7196
rect 46406 7155 46416 7162
rect 46405 7109 46416 7155
rect 46586 7155 46596 7162
rect 46778 7155 46788 7162
rect 46406 7102 46416 7109
rect 46586 7109 46597 7155
rect 46777 7109 46788 7155
rect 46958 7155 46968 7162
rect 46586 7102 46596 7109
rect 46778 7102 46788 7109
rect 46958 7109 46969 7155
rect 46958 7102 46968 7109
rect 47024 6794 47094 7196
rect 47150 7155 47160 7162
rect 47149 7109 47160 7155
rect 47330 7155 47340 7162
rect 47522 7155 47532 7162
rect 47150 7102 47160 7109
rect 47330 7109 47341 7155
rect 47521 7109 47532 7155
rect 47702 7155 47712 7162
rect 47330 7102 47340 7109
rect 47522 7102 47532 7109
rect 47702 7109 47713 7155
rect 47702 7102 47712 7109
rect 47768 6794 47838 7196
rect 47894 7155 47904 7162
rect 47893 7109 47904 7155
rect 48074 7155 48084 7162
rect 48266 7155 48276 7162
rect 47894 7102 47904 7109
rect 48074 7109 48085 7155
rect 48265 7109 48276 7155
rect 48446 7155 48456 7162
rect 48074 7102 48084 7109
rect 48266 7102 48276 7109
rect 48446 7109 48457 7155
rect 48446 7102 48456 7109
rect 48512 6794 48582 7196
rect 48638 7155 48648 7162
rect 48637 7109 48648 7155
rect 48818 7155 48828 7162
rect 49010 7155 49020 7162
rect 48638 7102 48648 7109
rect 48818 7109 48829 7155
rect 49009 7109 49020 7155
rect 49190 7155 49200 7162
rect 48818 7102 48828 7109
rect 49010 7102 49020 7109
rect 49190 7109 49201 7155
rect 49190 7102 49200 7109
rect 49256 6794 49326 7196
rect 49382 7155 49392 7162
rect 49381 7109 49392 7155
rect 49562 7155 49572 7162
rect 49754 7155 49764 7162
rect 49382 7102 49392 7109
rect 49562 7109 49573 7155
rect 49753 7109 49764 7155
rect 49934 7155 49944 7162
rect 49562 7102 49572 7109
rect 49754 7102 49764 7109
rect 49934 7109 49945 7155
rect 49934 7102 49944 7109
rect 50000 6794 50070 7196
rect 50126 7155 50136 7162
rect 50125 7109 50136 7155
rect 50306 7155 50316 7162
rect 50498 7155 50508 7162
rect 50126 7102 50136 7109
rect 50306 7109 50317 7155
rect 50497 7109 50508 7155
rect 50678 7155 50688 7162
rect 50306 7102 50316 7109
rect 50498 7102 50508 7109
rect 50678 7109 50689 7155
rect 50678 7102 50688 7109
rect 50744 6794 50814 7196
rect 50870 7155 50880 7162
rect 50869 7109 50880 7155
rect 51050 7155 51060 7162
rect 50870 7102 50880 7109
rect 51050 7109 51061 7155
rect 51050 7102 51060 7109
rect 40722 6468 40815 6480
rect 39824 6309 39892 6325
rect 40236 6225 40246 6259
rect 39958 6219 40246 6225
rect 39958 6153 39970 6219
rect 40042 6153 40246 6219
rect 39958 6149 40246 6153
rect 39958 6147 40054 6149
rect 40236 6109 40246 6149
rect 40392 6109 40402 6259
rect 40236 5825 40246 5859
rect 39958 5819 40246 5825
rect 39958 5755 39970 5819
rect 40042 5755 40246 5819
rect 39958 5749 40246 5755
rect 40236 5709 40246 5749
rect 40392 5709 40402 5859
rect 40722 5692 40775 6468
rect 40809 5692 40815 6468
rect 40722 5680 40815 5692
rect 41027 6468 41187 6480
rect 41027 5692 41033 6468
rect 41067 5692 41147 6468
rect 41181 5692 41187 6468
rect 41027 5680 41187 5692
rect 41399 6468 41559 6480
rect 41399 5692 41405 6468
rect 41439 5692 41519 6468
rect 41553 5692 41559 6468
rect 41399 5680 41559 5692
rect 41771 6468 41931 6480
rect 41771 5692 41777 6468
rect 41811 5692 41891 6468
rect 41925 5692 41931 6468
rect 41771 5680 41931 5692
rect 42143 6468 42303 6480
rect 42143 5692 42149 6468
rect 42183 5692 42263 6468
rect 42297 5692 42303 6468
rect 42143 5680 42303 5692
rect 42515 6468 42675 6480
rect 42515 5692 42521 6468
rect 42555 5692 42635 6468
rect 42669 5692 42675 6468
rect 42515 5680 42675 5692
rect 42887 6468 43047 6480
rect 42887 5692 42893 6468
rect 42927 5692 43007 6468
rect 43041 5692 43047 6468
rect 42887 5680 43047 5692
rect 43259 6468 43419 6480
rect 43259 5692 43265 6468
rect 43299 5692 43379 6468
rect 43413 5692 43419 6468
rect 43259 5680 43419 5692
rect 43631 6468 43724 6480
rect 43631 5692 43637 6468
rect 43671 5692 43724 6468
rect 44660 6082 44732 6557
rect 45422 6522 45432 6794
rect 45714 6522 45724 6794
rect 46166 6522 46176 6794
rect 46458 6522 46468 6794
rect 46910 6522 46920 6794
rect 47202 6522 47212 6794
rect 47654 6522 47664 6794
rect 47946 6522 47956 6794
rect 48398 6522 48408 6794
rect 48690 6522 48700 6794
rect 49142 6522 49152 6794
rect 49434 6522 49444 6794
rect 49886 6522 49896 6794
rect 50178 6522 50188 6794
rect 50630 6522 50640 6794
rect 50922 6522 50932 6794
rect 45628 6101 45638 6135
rect 44660 5855 44677 6082
rect 43631 5680 43724 5692
rect 40236 5425 40246 5459
rect 39958 5419 40246 5425
rect 39958 5355 39970 5419
rect 40042 5355 40246 5419
rect 39958 5349 40246 5355
rect 40236 5309 40246 5349
rect 40392 5309 40402 5459
rect 40722 5444 40770 5680
rect 40825 5634 41017 5639
rect 40825 5593 40836 5634
rect 40826 5531 40836 5593
rect 40825 5490 40836 5531
rect 41006 5593 41017 5634
rect 41006 5531 41016 5593
rect 41006 5490 41017 5531
rect 40825 5485 41017 5490
rect 41072 5444 41142 5680
rect 41197 5634 41389 5639
rect 41197 5593 41208 5634
rect 41198 5531 41208 5593
rect 41197 5490 41208 5531
rect 41378 5593 41389 5634
rect 41378 5531 41388 5593
rect 41378 5490 41389 5531
rect 41197 5485 41389 5490
rect 41444 5444 41514 5680
rect 41569 5634 41761 5639
rect 41569 5593 41580 5634
rect 41570 5531 41580 5593
rect 41569 5490 41580 5531
rect 41750 5593 41761 5634
rect 41750 5531 41760 5593
rect 41750 5490 41761 5531
rect 41569 5485 41761 5490
rect 41816 5444 41886 5680
rect 41941 5634 42133 5639
rect 41941 5593 41952 5634
rect 41942 5531 41952 5593
rect 41941 5490 41952 5531
rect 42122 5593 42133 5634
rect 42122 5531 42132 5593
rect 42122 5490 42133 5531
rect 41941 5485 42133 5490
rect 42188 5444 42258 5680
rect 42313 5634 42505 5639
rect 42313 5593 42324 5634
rect 42314 5531 42324 5593
rect 42313 5490 42324 5531
rect 42494 5593 42505 5634
rect 42494 5531 42504 5593
rect 42494 5490 42505 5531
rect 42313 5485 42505 5490
rect 42560 5444 42630 5680
rect 42685 5634 42877 5639
rect 42685 5593 42696 5634
rect 42686 5531 42696 5593
rect 42685 5490 42696 5531
rect 42866 5593 42877 5634
rect 42866 5531 42876 5593
rect 42866 5490 42877 5531
rect 42685 5485 42877 5490
rect 42932 5444 43002 5680
rect 43057 5634 43249 5639
rect 43057 5593 43068 5634
rect 43058 5531 43068 5593
rect 43057 5490 43068 5531
rect 43238 5593 43249 5634
rect 43238 5531 43248 5593
rect 43238 5490 43249 5531
rect 43057 5485 43249 5490
rect 43304 5444 43374 5680
rect 43429 5634 43621 5639
rect 43429 5593 43440 5634
rect 43430 5531 43440 5593
rect 43429 5490 43440 5531
rect 43610 5593 43621 5634
rect 43610 5531 43620 5593
rect 43610 5490 43621 5531
rect 43429 5485 43621 5490
rect 43670 5444 43724 5680
rect 44152 5569 44162 5719
rect 44308 5685 44318 5719
rect 44671 5685 44677 5855
rect 44715 5855 44732 6082
rect 44978 6082 45638 6101
rect 44715 5685 44721 5855
rect 44308 5679 44596 5685
rect 44308 5613 44512 5679
rect 44584 5613 44596 5679
rect 44671 5673 44721 5685
rect 44978 5685 44995 6082
rect 45033 5685 45638 6082
rect 44978 5667 45638 5685
rect 45628 5635 45638 5667
rect 46122 5635 46132 6135
rect 44308 5609 44596 5613
rect 44308 5569 44318 5609
rect 44500 5607 44596 5609
rect 40722 5432 40815 5444
rect 39504 5291 39894 5309
rect 39504 4894 39521 5291
rect 39559 4894 39839 5291
rect 39877 4894 39894 5291
rect 40236 5025 40246 5059
rect 39958 5019 40246 5025
rect 39958 4955 39970 5019
rect 40042 4955 40246 5019
rect 39958 4949 40246 4955
rect 40236 4909 40246 4949
rect 40392 4909 40402 5059
rect 39504 4875 39894 4894
rect 40722 4656 40775 5432
rect 40809 4656 40815 5432
rect 40722 4644 40815 4656
rect 41027 5432 41187 5444
rect 41027 4656 41033 5432
rect 41067 4656 41147 5432
rect 41181 4656 41187 5432
rect 41027 4644 41187 4656
rect 41399 5432 41559 5444
rect 41399 4656 41405 5432
rect 41439 4656 41519 5432
rect 41553 4656 41559 5432
rect 41399 4644 41559 4656
rect 41771 5432 41931 5444
rect 41771 4656 41777 5432
rect 41811 4656 41891 5432
rect 41925 4656 41931 5432
rect 41771 4644 41931 4656
rect 42143 5432 42303 5444
rect 42143 4656 42149 5432
rect 42183 4656 42263 5432
rect 42297 4656 42303 5432
rect 42143 4644 42303 4656
rect 42515 5432 42675 5444
rect 42515 4656 42521 5432
rect 42555 4656 42635 5432
rect 42669 4656 42675 5432
rect 42515 4644 42675 4656
rect 42887 5432 43047 5444
rect 42887 4656 42893 5432
rect 42927 4656 43007 5432
rect 43041 4656 43047 5432
rect 42887 4644 43047 4656
rect 43259 5432 43419 5444
rect 43259 4656 43265 5432
rect 43299 4656 43379 5432
rect 43413 4656 43419 5432
rect 43259 4644 43419 4656
rect 43631 5432 43724 5444
rect 43631 4656 43637 5432
rect 43671 4656 43724 5432
rect 44152 5169 44162 5319
rect 44308 5285 44318 5319
rect 44308 5279 44596 5285
rect 44308 5215 44512 5279
rect 44584 5215 44596 5279
rect 44308 5209 44596 5215
rect 44308 5169 44318 5209
rect 44152 4769 44162 4919
rect 44308 4885 44318 4919
rect 44308 4879 44596 4885
rect 44308 4815 44512 4879
rect 44584 4815 44596 4879
rect 44308 4809 44596 4815
rect 44308 4769 44318 4809
rect 45842 4748 45852 5020
rect 46134 4748 46144 5020
rect 43631 4644 43724 4656
rect 40722 4408 40770 4644
rect 40825 4598 41017 4603
rect 40825 4557 40836 4598
rect 40826 4495 40836 4557
rect 40825 4454 40836 4495
rect 41006 4557 41017 4598
rect 41006 4495 41016 4557
rect 41006 4454 41017 4495
rect 40825 4449 41017 4454
rect 41072 4408 41142 4644
rect 41197 4598 41389 4603
rect 41197 4557 41208 4598
rect 41198 4495 41208 4557
rect 41197 4454 41208 4495
rect 41378 4557 41389 4598
rect 41378 4495 41388 4557
rect 41378 4454 41389 4495
rect 41197 4449 41389 4454
rect 41444 4408 41514 4644
rect 41569 4598 41761 4603
rect 41569 4557 41580 4598
rect 41570 4495 41580 4557
rect 41569 4454 41580 4495
rect 41750 4557 41761 4598
rect 41750 4495 41760 4557
rect 41750 4454 41761 4495
rect 41569 4449 41761 4454
rect 41816 4408 41886 4644
rect 41941 4598 42133 4603
rect 41941 4557 41952 4598
rect 41942 4495 41952 4557
rect 41941 4454 41952 4495
rect 42122 4557 42133 4598
rect 42122 4495 42132 4557
rect 42122 4454 42133 4495
rect 41941 4449 42133 4454
rect 42188 4408 42258 4644
rect 42313 4598 42505 4603
rect 42313 4557 42324 4598
rect 42314 4495 42324 4557
rect 42313 4454 42324 4495
rect 42494 4557 42505 4598
rect 42494 4495 42504 4557
rect 42494 4454 42505 4495
rect 42313 4449 42505 4454
rect 42560 4408 42630 4644
rect 42685 4598 42877 4603
rect 42685 4557 42696 4598
rect 42686 4495 42696 4557
rect 42685 4454 42696 4495
rect 42866 4557 42877 4598
rect 42866 4495 42876 4557
rect 42866 4454 42877 4495
rect 42685 4449 42877 4454
rect 42932 4408 43002 4644
rect 43057 4598 43249 4603
rect 43057 4557 43068 4598
rect 43058 4495 43068 4557
rect 43057 4454 43068 4495
rect 43238 4557 43249 4598
rect 43238 4495 43248 4557
rect 43238 4454 43249 4495
rect 43057 4449 43249 4454
rect 43304 4408 43374 4644
rect 43429 4598 43621 4603
rect 43429 4557 43440 4598
rect 43430 4495 43440 4557
rect 43429 4454 43440 4495
rect 43610 4557 43621 4598
rect 43610 4495 43620 4557
rect 43610 4454 43621 4495
rect 43429 4449 43621 4454
rect 43670 4408 43724 4644
rect 44660 4651 45050 4669
rect 40722 4396 40815 4408
rect 40722 3620 40775 4396
rect 40809 3620 40815 4396
rect 40722 3608 40815 3620
rect 41027 4396 41187 4408
rect 41027 3620 41033 4396
rect 41067 3620 41147 4396
rect 41181 3620 41187 4396
rect 41027 3608 41187 3620
rect 41399 4396 41559 4408
rect 41399 3620 41405 4396
rect 41439 3620 41519 4396
rect 41553 3620 41559 4396
rect 41399 3608 41559 3620
rect 41771 4396 41931 4408
rect 41771 3620 41777 4396
rect 41811 3620 41891 4396
rect 41925 3620 41931 4396
rect 41771 3608 41931 3620
rect 42143 4396 42303 4408
rect 42143 3620 42149 4396
rect 42183 3620 42263 4396
rect 42297 3620 42303 4396
rect 42143 3608 42303 3620
rect 42515 4396 42675 4408
rect 42515 3620 42521 4396
rect 42555 3620 42635 4396
rect 42669 3620 42675 4396
rect 42515 3608 42675 3620
rect 42887 4396 43047 4408
rect 42887 3620 42893 4396
rect 42927 3620 43007 4396
rect 43041 3620 43047 4396
rect 42887 3608 43047 3620
rect 43259 4396 43419 4408
rect 43259 3620 43265 4396
rect 43299 3620 43379 4396
rect 43413 3620 43419 4396
rect 43259 3608 43419 3620
rect 43631 4396 43724 4408
rect 43631 3620 43637 4396
rect 43671 3620 43724 4396
rect 44152 4369 44162 4519
rect 44308 4485 44318 4519
rect 44308 4479 44596 4485
rect 44308 4415 44512 4479
rect 44584 4415 44596 4479
rect 44308 4409 44596 4415
rect 44308 4369 44318 4409
rect 44660 4254 44677 4651
rect 44715 4254 44995 4651
rect 45033 4254 45050 4651
rect 45954 4359 46026 4748
rect 44660 4235 45050 4254
rect 45546 4132 45556 4306
rect 45730 4246 45740 4306
rect 45730 4240 45882 4246
rect 45730 4186 45812 4240
rect 45870 4186 45882 4240
rect 45730 4180 45882 4186
rect 45730 4132 45740 4180
rect 45954 3962 45971 4359
rect 46009 3962 46026 4359
rect 45954 3944 46026 3962
rect 45546 3732 45556 3906
rect 45730 3846 45740 3906
rect 45730 3840 45882 3846
rect 45730 3786 45812 3840
rect 45870 3786 45882 3840
rect 45730 3780 45882 3786
rect 45954 3828 46026 3846
rect 45730 3732 45740 3780
rect 43631 3608 43724 3620
rect 40722 3372 40770 3608
rect 40825 3562 41017 3567
rect 40825 3521 40836 3562
rect 40826 3459 40836 3521
rect 40825 3418 40836 3459
rect 41006 3521 41017 3562
rect 41006 3459 41016 3521
rect 41006 3418 41017 3459
rect 40825 3413 41017 3418
rect 41072 3372 41142 3608
rect 41197 3562 41389 3567
rect 41197 3521 41208 3562
rect 41198 3459 41208 3521
rect 41197 3418 41208 3459
rect 41378 3521 41389 3562
rect 41378 3459 41388 3521
rect 41378 3418 41389 3459
rect 41197 3413 41389 3418
rect 41444 3372 41514 3608
rect 41569 3562 41761 3567
rect 41569 3521 41580 3562
rect 41570 3459 41580 3521
rect 41569 3418 41580 3459
rect 41750 3521 41761 3562
rect 41750 3459 41760 3521
rect 41750 3418 41761 3459
rect 41569 3413 41761 3418
rect 41816 3372 41886 3608
rect 41941 3562 42133 3567
rect 41941 3521 41952 3562
rect 41942 3459 41952 3521
rect 41941 3418 41952 3459
rect 42122 3521 42133 3562
rect 42122 3459 42132 3521
rect 42122 3418 42133 3459
rect 41941 3413 42133 3418
rect 42188 3372 42258 3608
rect 42313 3562 42505 3567
rect 42313 3521 42324 3562
rect 42314 3459 42324 3521
rect 42313 3418 42324 3459
rect 42494 3521 42505 3562
rect 42494 3459 42504 3521
rect 42494 3418 42505 3459
rect 42313 3413 42505 3418
rect 42560 3372 42630 3608
rect 42685 3562 42877 3567
rect 42685 3521 42696 3562
rect 42686 3459 42696 3521
rect 42685 3418 42696 3459
rect 42866 3521 42877 3562
rect 42866 3459 42876 3521
rect 42866 3418 42877 3459
rect 42685 3413 42877 3418
rect 42932 3372 43002 3608
rect 43057 3562 43249 3567
rect 43057 3521 43068 3562
rect 43058 3459 43068 3521
rect 43057 3418 43068 3459
rect 43238 3521 43249 3562
rect 43238 3459 43248 3521
rect 43238 3418 43249 3459
rect 43057 3413 43249 3418
rect 43304 3372 43374 3608
rect 43429 3562 43621 3567
rect 43429 3521 43440 3562
rect 43430 3459 43440 3521
rect 43429 3418 43440 3459
rect 43610 3521 43621 3562
rect 43610 3459 43620 3521
rect 43610 3418 43621 3459
rect 43429 3413 43621 3418
rect 43670 3372 43724 3608
rect 40722 3360 40815 3372
rect 40722 2584 40775 3360
rect 40809 2584 40815 3360
rect 40722 2572 40815 2584
rect 41027 3360 41187 3372
rect 41027 2584 41033 3360
rect 41067 2584 41147 3360
rect 41181 2584 41187 3360
rect 41027 2572 41187 2584
rect 41399 3360 41559 3372
rect 41399 2584 41405 3360
rect 41439 2584 41519 3360
rect 41553 2584 41559 3360
rect 41399 2572 41559 2584
rect 41771 3360 41931 3372
rect 41771 2584 41777 3360
rect 41811 2584 41891 3360
rect 41925 2584 41931 3360
rect 41771 2572 41931 2584
rect 42143 3360 42303 3372
rect 42143 2584 42149 3360
rect 42183 2584 42263 3360
rect 42297 2584 42303 3360
rect 42143 2572 42303 2584
rect 42515 3360 42675 3372
rect 42515 2584 42521 3360
rect 42555 2584 42635 3360
rect 42669 2584 42675 3360
rect 42515 2572 42675 2584
rect 42887 3360 43047 3372
rect 42887 2584 42893 3360
rect 42927 2584 43007 3360
rect 43041 2584 43047 3360
rect 42887 2572 43047 2584
rect 43259 3360 43419 3372
rect 43259 2584 43265 3360
rect 43299 2584 43379 3360
rect 43413 2584 43419 3360
rect 43259 2572 43419 2584
rect 43631 3360 43724 3372
rect 43631 2584 43637 3360
rect 43671 2584 43724 3360
rect 45546 3332 45556 3506
rect 45730 3446 45740 3506
rect 45730 3440 45882 3446
rect 45730 3386 45812 3440
rect 45870 3386 45882 3440
rect 45730 3380 45882 3386
rect 45954 3431 45971 3828
rect 46009 3431 46026 3828
rect 45730 3332 45740 3380
rect 43631 2572 43724 2584
rect 40826 2531 40836 2536
rect 40825 2485 40836 2531
rect 41006 2531 41016 2536
rect 40826 2482 40836 2485
rect 41006 2485 41017 2531
rect 41006 2482 41016 2485
rect 41072 1888 41142 2572
rect 41198 2531 41208 2536
rect 41197 2485 41208 2531
rect 41378 2531 41388 2536
rect 41570 2531 41580 2536
rect 41198 2482 41208 2485
rect 41378 2485 41389 2531
rect 41569 2485 41580 2531
rect 41750 2531 41760 2536
rect 41378 2482 41388 2485
rect 41570 2482 41580 2485
rect 41750 2485 41761 2531
rect 41750 2482 41760 2485
rect 41816 2196 41886 2572
rect 41942 2531 41952 2536
rect 41941 2485 41952 2531
rect 42122 2531 42132 2536
rect 42314 2531 42324 2536
rect 41942 2482 41952 2485
rect 42122 2485 42133 2531
rect 42313 2485 42324 2531
rect 42494 2531 42504 2536
rect 42122 2482 42132 2485
rect 42314 2482 42324 2485
rect 42494 2485 42505 2531
rect 42494 2482 42504 2485
rect 42560 2196 42630 2572
rect 42686 2531 42696 2536
rect 42685 2485 42696 2531
rect 42866 2531 42876 2536
rect 43058 2531 43068 2536
rect 42686 2482 42696 2485
rect 42866 2485 42877 2531
rect 43057 2485 43068 2531
rect 43238 2531 43248 2536
rect 42866 2482 42876 2485
rect 43058 2482 43068 2485
rect 43238 2485 43249 2531
rect 43238 2482 43248 2485
rect 41806 2016 41816 2196
rect 42630 2016 42640 2196
rect 40824 1878 41390 1888
rect 40824 1832 40836 1878
rect 40825 1827 40836 1832
rect 40826 1822 40836 1827
rect 41006 1832 41208 1878
rect 41006 1827 41017 1832
rect 41006 1822 41016 1827
rect 40720 1795 40794 1796
rect 41072 1795 41142 1832
rect 41197 1827 41208 1832
rect 41198 1822 41208 1827
rect 41378 1832 41390 1878
rect 41570 1873 41580 1878
rect 41378 1827 41389 1832
rect 41569 1827 41580 1873
rect 41750 1873 41760 1878
rect 41378 1822 41388 1827
rect 41570 1822 41580 1827
rect 41750 1827 41761 1873
rect 41750 1822 41760 1827
rect 41444 1795 41514 1796
rect 41816 1795 41886 2016
rect 41942 1873 41952 1878
rect 41941 1827 41952 1873
rect 42122 1873 42132 1878
rect 42314 1873 42324 1878
rect 41942 1822 41952 1827
rect 42122 1827 42133 1873
rect 42313 1827 42324 1873
rect 42494 1873 42504 1878
rect 42122 1822 42132 1827
rect 42314 1822 42324 1827
rect 42494 1827 42505 1873
rect 42494 1822 42504 1827
rect 42188 1795 42258 1796
rect 42560 1795 42630 2016
rect 43304 1888 43374 2572
rect 43430 2531 43440 2536
rect 43429 2485 43440 2531
rect 43610 2531 43620 2536
rect 43430 2482 43440 2485
rect 43610 2485 43621 2531
rect 43610 2482 43620 2485
rect 43932 2340 43942 2612
rect 44224 2340 44234 2612
rect 44676 2340 44686 2612
rect 44968 2340 44978 2612
rect 45420 2340 45430 2612
rect 45712 2340 45722 2612
rect 45954 2384 46026 3431
rect 43056 1878 43622 1888
rect 42686 1873 42696 1878
rect 42685 1827 42696 1873
rect 42866 1873 42876 1878
rect 42686 1822 42696 1827
rect 42866 1827 42877 1873
rect 43056 1832 43068 1878
rect 43057 1827 43068 1832
rect 42866 1822 42876 1827
rect 43058 1822 43068 1827
rect 43238 1832 43440 1878
rect 43238 1827 43249 1832
rect 43238 1822 43248 1827
rect 42932 1795 43002 1796
rect 43304 1795 43374 1832
rect 43429 1827 43440 1832
rect 43430 1822 43440 1827
rect 43610 1832 43622 1878
rect 43802 1873 43812 1878
rect 43610 1827 43621 1832
rect 43801 1827 43812 1873
rect 43982 1873 43992 1878
rect 43610 1822 43620 1827
rect 43802 1822 43812 1827
rect 43982 1827 43993 1873
rect 43982 1822 43992 1827
rect 43676 1795 43746 1796
rect 44048 1795 44118 2340
rect 44174 1873 44184 1878
rect 44173 1827 44184 1873
rect 44354 1873 44364 1878
rect 44546 1873 44556 1878
rect 44174 1822 44184 1827
rect 44354 1827 44365 1873
rect 44545 1827 44556 1873
rect 44726 1873 44736 1878
rect 44354 1822 44364 1827
rect 44546 1822 44556 1827
rect 44726 1827 44737 1873
rect 44726 1822 44736 1827
rect 44420 1795 44490 1796
rect 44792 1795 44862 2340
rect 44918 1873 44928 1878
rect 44917 1827 44928 1873
rect 45098 1873 45108 1878
rect 45290 1873 45300 1878
rect 44918 1822 44928 1827
rect 45098 1827 45109 1873
rect 45289 1827 45300 1873
rect 45470 1873 45480 1878
rect 45098 1822 45108 1827
rect 45290 1822 45300 1827
rect 45470 1827 45481 1873
rect 45470 1822 45480 1827
rect 45164 1795 45234 1796
rect 45536 1795 45606 2340
rect 45952 2336 46026 2384
rect 46164 2340 46174 2612
rect 46456 2340 46466 2612
rect 46908 2340 46918 2612
rect 47200 2340 47210 2612
rect 47652 2340 47662 2612
rect 47944 2340 47954 2612
rect 48396 2340 48406 2612
rect 48688 2340 48698 2612
rect 49140 2340 49150 2612
rect 49432 2340 49442 2612
rect 45912 2324 46026 2336
rect 45816 2050 45826 2324
rect 46104 2050 46114 2324
rect 45662 1873 45672 1878
rect 45661 1827 45672 1873
rect 45842 1873 45852 1878
rect 46034 1873 46044 1878
rect 45662 1822 45672 1827
rect 45842 1827 45853 1873
rect 46033 1827 46044 1873
rect 46214 1873 46224 1878
rect 45842 1822 45852 1827
rect 46034 1822 46044 1827
rect 46214 1827 46225 1873
rect 46214 1822 46224 1827
rect 45908 1795 45978 1796
rect 46280 1795 46350 2340
rect 46406 1873 46416 1878
rect 46405 1827 46416 1873
rect 46586 1873 46596 1878
rect 46778 1873 46788 1878
rect 46406 1822 46416 1827
rect 46586 1827 46597 1873
rect 46777 1827 46788 1873
rect 46958 1873 46968 1878
rect 46586 1822 46596 1827
rect 46778 1822 46788 1827
rect 46958 1827 46969 1873
rect 46958 1822 46968 1827
rect 46652 1795 46722 1796
rect 47024 1795 47094 2340
rect 47150 1873 47160 1878
rect 47149 1827 47160 1873
rect 47330 1873 47340 1878
rect 47522 1873 47532 1878
rect 47150 1822 47160 1827
rect 47330 1827 47341 1873
rect 47521 1827 47532 1873
rect 47702 1873 47712 1878
rect 47330 1822 47340 1827
rect 47522 1822 47532 1827
rect 47702 1827 47713 1873
rect 47702 1822 47712 1827
rect 47396 1795 47466 1796
rect 47768 1795 47838 2340
rect 47894 1873 47904 1878
rect 47893 1827 47904 1873
rect 48074 1873 48084 1878
rect 48266 1873 48276 1878
rect 47894 1822 47904 1827
rect 48074 1827 48085 1873
rect 48265 1827 48276 1873
rect 48446 1873 48456 1878
rect 48074 1822 48084 1827
rect 48266 1822 48276 1827
rect 48446 1827 48457 1873
rect 48446 1822 48456 1827
rect 48140 1795 48210 1796
rect 48512 1795 48582 2340
rect 48638 1873 48648 1878
rect 48637 1827 48648 1873
rect 48818 1873 48828 1878
rect 49010 1873 49020 1878
rect 48638 1822 48648 1827
rect 48818 1827 48829 1873
rect 49009 1827 49020 1873
rect 49190 1873 49200 1878
rect 48818 1822 48828 1827
rect 49010 1822 49020 1827
rect 49190 1827 49201 1873
rect 49190 1822 49200 1827
rect 48884 1795 48954 1796
rect 49256 1795 49326 2340
rect 49382 1873 49392 1878
rect 49381 1827 49392 1873
rect 49562 1873 49572 1878
rect 49382 1822 49392 1827
rect 49562 1827 49573 1873
rect 49562 1822 49572 1827
rect 49604 1795 49678 1808
rect 40720 1783 40815 1795
rect 40720 1607 40775 1783
rect 40809 1607 40815 1783
rect 40720 1595 40815 1607
rect 41027 1783 41187 1795
rect 41027 1607 41033 1783
rect 41067 1607 41147 1783
rect 41181 1607 41187 1783
rect 41027 1595 41187 1607
rect 41399 1783 41559 1795
rect 41399 1607 41405 1783
rect 41439 1607 41519 1783
rect 41553 1607 41559 1783
rect 41399 1595 41559 1607
rect 41771 1783 41931 1795
rect 41771 1607 41777 1783
rect 41811 1607 41891 1783
rect 41925 1607 41931 1783
rect 41771 1595 41931 1607
rect 42143 1783 42303 1795
rect 42143 1607 42149 1783
rect 42183 1607 42263 1783
rect 42297 1607 42303 1783
rect 42143 1595 42303 1607
rect 42515 1783 42675 1795
rect 42515 1607 42521 1783
rect 42555 1607 42635 1783
rect 42669 1607 42675 1783
rect 42515 1595 42675 1607
rect 42887 1783 43047 1795
rect 42887 1607 42893 1783
rect 42927 1607 43007 1783
rect 43041 1607 43047 1783
rect 42887 1595 43047 1607
rect 43259 1783 43419 1795
rect 43259 1607 43265 1783
rect 43299 1607 43379 1783
rect 43413 1607 43419 1783
rect 43259 1595 43419 1607
rect 43631 1783 43791 1795
rect 43631 1607 43637 1783
rect 43671 1607 43751 1783
rect 43785 1607 43791 1783
rect 43631 1595 43791 1607
rect 44003 1783 44163 1795
rect 44003 1607 44009 1783
rect 44043 1607 44123 1783
rect 44157 1607 44163 1783
rect 44003 1595 44163 1607
rect 44375 1783 44535 1795
rect 44375 1607 44381 1783
rect 44415 1607 44495 1783
rect 44529 1607 44535 1783
rect 44375 1595 44535 1607
rect 44747 1783 44907 1795
rect 44747 1607 44753 1783
rect 44787 1607 44867 1783
rect 44901 1607 44907 1783
rect 44747 1595 44907 1607
rect 45119 1783 45279 1795
rect 45119 1607 45125 1783
rect 45159 1607 45239 1783
rect 45273 1607 45279 1783
rect 45119 1595 45279 1607
rect 45491 1783 45651 1795
rect 45491 1607 45497 1783
rect 45531 1607 45611 1783
rect 45645 1607 45651 1783
rect 45491 1595 45651 1607
rect 45863 1783 46023 1795
rect 45863 1607 45869 1783
rect 45903 1607 45983 1783
rect 46017 1607 46023 1783
rect 45863 1595 46023 1607
rect 46235 1783 46395 1795
rect 46235 1607 46241 1783
rect 46275 1607 46355 1783
rect 46389 1607 46395 1783
rect 46235 1595 46395 1607
rect 46607 1783 46767 1795
rect 46607 1607 46613 1783
rect 46647 1607 46727 1783
rect 46761 1607 46767 1783
rect 46607 1595 46767 1607
rect 46979 1783 47139 1795
rect 46979 1607 46985 1783
rect 47019 1607 47099 1783
rect 47133 1607 47139 1783
rect 46979 1595 47139 1607
rect 47351 1783 47511 1795
rect 47351 1607 47357 1783
rect 47391 1607 47471 1783
rect 47505 1607 47511 1783
rect 47351 1595 47511 1607
rect 47723 1783 47883 1795
rect 47723 1607 47729 1783
rect 47763 1607 47843 1783
rect 47877 1607 47883 1783
rect 47723 1595 47883 1607
rect 48095 1783 48255 1795
rect 48095 1607 48101 1783
rect 48135 1607 48215 1783
rect 48249 1607 48255 1783
rect 48095 1595 48255 1607
rect 48467 1783 48627 1795
rect 48467 1607 48473 1783
rect 48507 1607 48587 1783
rect 48621 1607 48627 1783
rect 48467 1595 48627 1607
rect 48839 1783 48999 1795
rect 48839 1607 48845 1783
rect 48879 1607 48959 1783
rect 48993 1607 48999 1783
rect 48839 1595 48999 1607
rect 49211 1783 49371 1795
rect 49211 1607 49217 1783
rect 49251 1607 49331 1783
rect 49365 1607 49371 1783
rect 49211 1595 49371 1607
rect 49583 1783 49678 1795
rect 49583 1607 49589 1783
rect 49623 1607 49678 1783
rect 49583 1595 49678 1607
rect 40720 1377 40794 1595
rect 41072 1564 41142 1595
rect 40824 1558 41390 1564
rect 40824 1414 40836 1558
rect 41006 1414 41208 1558
rect 41378 1414 41390 1558
rect 40824 1408 41390 1414
rect 41072 1377 41142 1408
rect 41444 1377 41514 1595
rect 41569 1558 41761 1563
rect 41569 1517 41580 1558
rect 41570 1455 41580 1517
rect 41569 1414 41580 1455
rect 41750 1517 41761 1558
rect 41750 1455 41760 1517
rect 41750 1414 41761 1455
rect 41569 1409 41761 1414
rect 41816 1377 41886 1595
rect 41941 1558 42133 1563
rect 41941 1517 41952 1558
rect 41942 1455 41952 1517
rect 41941 1414 41952 1455
rect 42122 1517 42133 1558
rect 42122 1455 42132 1517
rect 42122 1414 42133 1455
rect 41941 1409 42133 1414
rect 42188 1377 42258 1595
rect 42313 1558 42505 1563
rect 42313 1517 42324 1558
rect 42314 1455 42324 1517
rect 42313 1414 42324 1455
rect 42494 1517 42505 1558
rect 42494 1455 42504 1517
rect 42494 1414 42505 1455
rect 42313 1409 42505 1414
rect 42560 1377 42630 1595
rect 42685 1558 42877 1563
rect 42685 1517 42696 1558
rect 42686 1455 42696 1517
rect 42685 1414 42696 1455
rect 42866 1517 42877 1558
rect 42866 1455 42876 1517
rect 42866 1414 42877 1455
rect 42685 1409 42877 1414
rect 42932 1377 43002 1595
rect 43304 1564 43374 1595
rect 43056 1558 43622 1564
rect 43056 1414 43068 1558
rect 43238 1414 43440 1558
rect 43610 1414 43622 1558
rect 43056 1408 43622 1414
rect 43304 1377 43374 1408
rect 43676 1377 43746 1595
rect 43801 1558 43993 1563
rect 43801 1517 43812 1558
rect 43802 1455 43812 1517
rect 43801 1414 43812 1455
rect 43982 1517 43993 1558
rect 43982 1455 43992 1517
rect 43982 1414 43993 1455
rect 43801 1409 43993 1414
rect 44048 1377 44118 1595
rect 44173 1558 44365 1563
rect 44173 1517 44184 1558
rect 44174 1455 44184 1517
rect 44173 1414 44184 1455
rect 44354 1517 44365 1558
rect 44354 1455 44364 1517
rect 44354 1414 44365 1455
rect 44173 1409 44365 1414
rect 44420 1377 44490 1595
rect 44545 1558 44737 1563
rect 44545 1517 44556 1558
rect 44546 1455 44556 1517
rect 44545 1414 44556 1455
rect 44726 1517 44737 1558
rect 44726 1455 44736 1517
rect 44726 1414 44737 1455
rect 44545 1409 44737 1414
rect 44792 1377 44862 1595
rect 44917 1558 45109 1563
rect 44917 1517 44928 1558
rect 44918 1455 44928 1517
rect 44917 1414 44928 1455
rect 45098 1517 45109 1558
rect 45098 1455 45108 1517
rect 45098 1414 45109 1455
rect 44917 1409 45109 1414
rect 45164 1377 45234 1595
rect 45289 1558 45481 1563
rect 45289 1517 45300 1558
rect 45290 1455 45300 1517
rect 45289 1414 45300 1455
rect 45470 1517 45481 1558
rect 45470 1455 45480 1517
rect 45470 1414 45481 1455
rect 45289 1409 45481 1414
rect 45536 1377 45606 1595
rect 45661 1558 45853 1563
rect 45661 1517 45672 1558
rect 45662 1455 45672 1517
rect 45661 1414 45672 1455
rect 45842 1517 45853 1558
rect 45842 1455 45852 1517
rect 45842 1414 45853 1455
rect 45661 1409 45853 1414
rect 45908 1377 45978 1595
rect 46033 1558 46225 1563
rect 46033 1517 46044 1558
rect 46034 1455 46044 1517
rect 46033 1414 46044 1455
rect 46214 1517 46225 1558
rect 46214 1455 46224 1517
rect 46214 1414 46225 1455
rect 46033 1409 46225 1414
rect 46280 1377 46350 1595
rect 46405 1558 46597 1563
rect 46405 1517 46416 1558
rect 46406 1455 46416 1517
rect 46405 1414 46416 1455
rect 46586 1517 46597 1558
rect 46586 1455 46596 1517
rect 46586 1414 46597 1455
rect 46405 1409 46597 1414
rect 46652 1377 46722 1595
rect 46777 1558 46969 1563
rect 46777 1517 46788 1558
rect 46778 1455 46788 1517
rect 46777 1414 46788 1455
rect 46958 1517 46969 1558
rect 46958 1455 46968 1517
rect 46958 1414 46969 1455
rect 46777 1409 46969 1414
rect 47024 1377 47094 1595
rect 47149 1558 47341 1563
rect 47149 1517 47160 1558
rect 47150 1455 47160 1517
rect 47149 1414 47160 1455
rect 47330 1517 47341 1558
rect 47330 1455 47340 1517
rect 47330 1414 47341 1455
rect 47149 1409 47341 1414
rect 47396 1377 47466 1595
rect 47521 1558 47713 1563
rect 47521 1517 47532 1558
rect 47522 1455 47532 1517
rect 47521 1414 47532 1455
rect 47702 1517 47713 1558
rect 47702 1455 47712 1517
rect 47702 1414 47713 1455
rect 47521 1409 47713 1414
rect 47768 1377 47838 1595
rect 47893 1558 48085 1563
rect 47893 1517 47904 1558
rect 47894 1455 47904 1517
rect 47893 1414 47904 1455
rect 48074 1517 48085 1558
rect 48074 1455 48084 1517
rect 48074 1414 48085 1455
rect 47893 1409 48085 1414
rect 48140 1377 48210 1595
rect 48265 1558 48457 1563
rect 48265 1517 48276 1558
rect 48266 1455 48276 1517
rect 48265 1414 48276 1455
rect 48446 1517 48457 1558
rect 48446 1455 48456 1517
rect 48446 1414 48457 1455
rect 48265 1409 48457 1414
rect 48512 1377 48582 1595
rect 48637 1558 48829 1563
rect 48637 1517 48648 1558
rect 48638 1455 48648 1517
rect 48637 1414 48648 1455
rect 48818 1517 48829 1558
rect 48818 1455 48828 1517
rect 48818 1414 48829 1455
rect 48637 1409 48829 1414
rect 48884 1377 48954 1595
rect 49009 1558 49201 1563
rect 49009 1517 49020 1558
rect 49010 1455 49020 1517
rect 49009 1414 49020 1455
rect 49190 1517 49201 1558
rect 49190 1455 49200 1517
rect 49190 1414 49201 1455
rect 49009 1409 49201 1414
rect 49256 1377 49326 1595
rect 49381 1558 49573 1563
rect 49381 1517 49392 1558
rect 49382 1455 49392 1517
rect 49381 1414 49392 1455
rect 49562 1517 49573 1558
rect 49562 1455 49572 1517
rect 49562 1414 49573 1455
rect 49381 1409 49573 1414
rect 49604 1377 49678 1595
rect 40720 1365 40815 1377
rect 40720 1189 40775 1365
rect 40809 1189 40815 1365
rect 40720 1177 40815 1189
rect 41027 1365 41187 1377
rect 41027 1189 41033 1365
rect 41067 1189 41147 1365
rect 41181 1189 41187 1365
rect 41027 1177 41187 1189
rect 41399 1365 41559 1377
rect 41399 1189 41405 1365
rect 41439 1189 41519 1365
rect 41553 1189 41559 1365
rect 41399 1177 41559 1189
rect 41771 1365 41931 1377
rect 41771 1189 41777 1365
rect 41811 1189 41891 1365
rect 41925 1189 41931 1365
rect 41771 1177 41931 1189
rect 42143 1365 42303 1377
rect 42143 1189 42149 1365
rect 42183 1189 42263 1365
rect 42297 1189 42303 1365
rect 42143 1177 42303 1189
rect 42515 1365 42675 1377
rect 42515 1189 42521 1365
rect 42555 1189 42635 1365
rect 42669 1189 42675 1365
rect 42515 1177 42675 1189
rect 42887 1365 43047 1377
rect 42887 1189 42893 1365
rect 42927 1189 43007 1365
rect 43041 1189 43047 1365
rect 42887 1177 43047 1189
rect 43259 1365 43419 1377
rect 43259 1189 43265 1365
rect 43299 1189 43379 1365
rect 43413 1189 43419 1365
rect 43259 1177 43419 1189
rect 43631 1365 43791 1377
rect 43631 1189 43637 1365
rect 43671 1189 43751 1365
rect 43785 1189 43791 1365
rect 43631 1177 43791 1189
rect 44003 1365 44163 1377
rect 44003 1189 44009 1365
rect 44043 1189 44123 1365
rect 44157 1189 44163 1365
rect 44003 1177 44163 1189
rect 44375 1365 44535 1377
rect 44375 1189 44381 1365
rect 44415 1189 44495 1365
rect 44529 1189 44535 1365
rect 44375 1177 44535 1189
rect 44747 1365 44907 1377
rect 44747 1189 44753 1365
rect 44787 1189 44867 1365
rect 44901 1189 44907 1365
rect 44747 1177 44907 1189
rect 45119 1365 45279 1377
rect 45119 1189 45125 1365
rect 45159 1189 45239 1365
rect 45273 1189 45279 1365
rect 45119 1177 45279 1189
rect 45491 1365 45651 1377
rect 45491 1189 45497 1365
rect 45531 1189 45611 1365
rect 45645 1189 45651 1365
rect 45491 1177 45651 1189
rect 45863 1365 46023 1377
rect 45863 1189 45869 1365
rect 45903 1189 45983 1365
rect 46017 1189 46023 1365
rect 45863 1177 46023 1189
rect 46235 1365 46395 1377
rect 46235 1189 46241 1365
rect 46275 1189 46355 1365
rect 46389 1189 46395 1365
rect 46235 1177 46395 1189
rect 46607 1365 46767 1377
rect 46607 1189 46613 1365
rect 46647 1189 46727 1365
rect 46761 1189 46767 1365
rect 46607 1177 46767 1189
rect 46979 1365 47139 1377
rect 46979 1189 46985 1365
rect 47019 1189 47099 1365
rect 47133 1189 47139 1365
rect 46979 1177 47139 1189
rect 47351 1365 47511 1377
rect 47351 1189 47357 1365
rect 47391 1189 47471 1365
rect 47505 1189 47511 1365
rect 47351 1177 47511 1189
rect 47723 1365 47883 1377
rect 47723 1189 47729 1365
rect 47763 1189 47843 1365
rect 47877 1189 47883 1365
rect 47723 1177 47883 1189
rect 48095 1365 48255 1377
rect 48095 1189 48101 1365
rect 48135 1189 48215 1365
rect 48249 1189 48255 1365
rect 48095 1177 48255 1189
rect 48467 1365 48627 1377
rect 48467 1189 48473 1365
rect 48507 1189 48587 1365
rect 48621 1189 48627 1365
rect 48467 1177 48627 1189
rect 48839 1365 48999 1377
rect 48839 1189 48845 1365
rect 48879 1189 48959 1365
rect 48993 1189 48999 1365
rect 48839 1177 48999 1189
rect 49211 1365 49371 1377
rect 49211 1189 49217 1365
rect 49251 1189 49331 1365
rect 49365 1189 49371 1365
rect 49211 1177 49371 1189
rect 49583 1365 49678 1377
rect 49583 1189 49589 1365
rect 49623 1189 49678 1365
rect 49583 1177 49678 1189
rect 40720 959 40794 1177
rect 41072 1146 41142 1177
rect 40824 1140 41390 1146
rect 40824 996 40836 1140
rect 41006 996 41208 1140
rect 41378 996 41390 1140
rect 40824 990 41390 996
rect 41072 959 41142 990
rect 41444 959 41514 1177
rect 41569 1140 41761 1145
rect 41569 1099 41580 1140
rect 41570 1037 41580 1099
rect 41569 996 41580 1037
rect 41750 1099 41761 1140
rect 41750 1037 41760 1099
rect 41750 996 41761 1037
rect 41569 991 41761 996
rect 41816 959 41886 1177
rect 41941 1140 42133 1145
rect 41941 1099 41952 1140
rect 41942 1037 41952 1099
rect 41941 996 41952 1037
rect 42122 1099 42133 1140
rect 42122 1037 42132 1099
rect 42122 996 42133 1037
rect 41941 991 42133 996
rect 42188 959 42258 1177
rect 42313 1140 42505 1145
rect 42313 1099 42324 1140
rect 42314 1037 42324 1099
rect 42313 996 42324 1037
rect 42494 1099 42505 1140
rect 42494 1037 42504 1099
rect 42494 996 42505 1037
rect 42313 991 42505 996
rect 42560 959 42630 1177
rect 42685 1140 42877 1145
rect 42685 1099 42696 1140
rect 42686 1037 42696 1099
rect 42685 996 42696 1037
rect 42866 1099 42877 1140
rect 42866 1037 42876 1099
rect 42866 996 42877 1037
rect 42685 991 42877 996
rect 42932 959 43002 1177
rect 43304 1146 43374 1177
rect 43056 1140 43622 1146
rect 43056 996 43068 1140
rect 43238 996 43440 1140
rect 43610 996 43622 1140
rect 43056 990 43622 996
rect 43304 959 43374 990
rect 43676 959 43746 1177
rect 43801 1140 43993 1145
rect 43801 1099 43812 1140
rect 43802 1037 43812 1099
rect 43801 996 43812 1037
rect 43982 1099 43993 1140
rect 43982 1037 43992 1099
rect 43982 996 43993 1037
rect 43801 991 43993 996
rect 44048 959 44118 1177
rect 44173 1140 44365 1145
rect 44173 1099 44184 1140
rect 44174 1037 44184 1099
rect 44173 996 44184 1037
rect 44354 1099 44365 1140
rect 44354 1037 44364 1099
rect 44354 996 44365 1037
rect 44173 991 44365 996
rect 44420 959 44490 1177
rect 44545 1140 44737 1145
rect 44545 1099 44556 1140
rect 44546 1037 44556 1099
rect 44545 996 44556 1037
rect 44726 1099 44737 1140
rect 44726 1037 44736 1099
rect 44726 996 44737 1037
rect 44545 991 44737 996
rect 44792 959 44862 1177
rect 44917 1140 45109 1145
rect 44917 1099 44928 1140
rect 44918 1037 44928 1099
rect 44917 996 44928 1037
rect 45098 1099 45109 1140
rect 45098 1037 45108 1099
rect 45098 996 45109 1037
rect 44917 991 45109 996
rect 45164 959 45234 1177
rect 45289 1140 45481 1145
rect 45289 1099 45300 1140
rect 45290 1037 45300 1099
rect 45289 996 45300 1037
rect 45470 1099 45481 1140
rect 45470 1037 45480 1099
rect 45470 996 45481 1037
rect 45289 991 45481 996
rect 45536 959 45606 1177
rect 45661 1140 45853 1145
rect 45661 1099 45672 1140
rect 45662 1037 45672 1099
rect 45661 996 45672 1037
rect 45842 1099 45853 1140
rect 45842 1037 45852 1099
rect 45842 996 45853 1037
rect 45661 991 45853 996
rect 45908 959 45978 1177
rect 46033 1140 46225 1145
rect 46033 1099 46044 1140
rect 46034 1037 46044 1099
rect 46033 996 46044 1037
rect 46214 1099 46225 1140
rect 46214 1037 46224 1099
rect 46214 996 46225 1037
rect 46033 991 46225 996
rect 46280 959 46350 1177
rect 46405 1140 46597 1145
rect 46405 1099 46416 1140
rect 46406 1037 46416 1099
rect 46405 996 46416 1037
rect 46586 1099 46597 1140
rect 46586 1037 46596 1099
rect 46586 996 46597 1037
rect 46405 991 46597 996
rect 46652 959 46722 1177
rect 46777 1140 46969 1145
rect 46777 1099 46788 1140
rect 46778 1037 46788 1099
rect 46777 996 46788 1037
rect 46958 1099 46969 1140
rect 46958 1037 46968 1099
rect 46958 996 46969 1037
rect 46777 991 46969 996
rect 47024 959 47094 1177
rect 47149 1140 47341 1145
rect 47149 1099 47160 1140
rect 47150 1037 47160 1099
rect 47149 996 47160 1037
rect 47330 1099 47341 1140
rect 47330 1037 47340 1099
rect 47330 996 47341 1037
rect 47149 991 47341 996
rect 47396 959 47466 1177
rect 47521 1140 47713 1145
rect 47521 1099 47532 1140
rect 47522 1037 47532 1099
rect 47521 996 47532 1037
rect 47702 1099 47713 1140
rect 47702 1037 47712 1099
rect 47702 996 47713 1037
rect 47521 991 47713 996
rect 47768 959 47838 1177
rect 47893 1140 48085 1145
rect 47893 1099 47904 1140
rect 47894 1037 47904 1099
rect 47893 996 47904 1037
rect 48074 1099 48085 1140
rect 48074 1037 48084 1099
rect 48074 996 48085 1037
rect 47893 991 48085 996
rect 48140 959 48210 1177
rect 48265 1140 48457 1145
rect 48265 1099 48276 1140
rect 48266 1037 48276 1099
rect 48265 996 48276 1037
rect 48446 1099 48457 1140
rect 48446 1037 48456 1099
rect 48446 996 48457 1037
rect 48265 991 48457 996
rect 48512 959 48582 1177
rect 48637 1140 48829 1145
rect 48637 1099 48648 1140
rect 48638 1037 48648 1099
rect 48637 996 48648 1037
rect 48818 1099 48829 1140
rect 48818 1037 48828 1099
rect 48818 996 48829 1037
rect 48637 991 48829 996
rect 48884 959 48954 1177
rect 49009 1140 49201 1145
rect 49009 1099 49020 1140
rect 49010 1037 49020 1099
rect 49009 996 49020 1037
rect 49190 1099 49201 1140
rect 49190 1037 49200 1099
rect 49190 996 49201 1037
rect 49009 991 49201 996
rect 49256 959 49326 1177
rect 49381 1140 49573 1145
rect 49381 1099 49392 1140
rect 49382 1037 49392 1099
rect 49381 996 49392 1037
rect 49562 1099 49573 1140
rect 49562 1037 49572 1099
rect 49562 996 49573 1037
rect 49381 991 49573 996
rect 49604 959 49678 1177
rect 40720 947 40815 959
rect 40720 771 40775 947
rect 40809 771 40815 947
rect 40720 759 40815 771
rect 41027 947 41187 959
rect 41027 771 41033 947
rect 41067 771 41147 947
rect 41181 771 41187 947
rect 41027 759 41187 771
rect 41399 947 41559 959
rect 41399 771 41405 947
rect 41439 771 41519 947
rect 41553 771 41559 947
rect 41399 759 41559 771
rect 41771 947 41931 959
rect 41771 771 41777 947
rect 41811 771 41891 947
rect 41925 771 41931 947
rect 41771 759 41931 771
rect 42143 947 42303 959
rect 42143 771 42149 947
rect 42183 771 42263 947
rect 42297 771 42303 947
rect 42143 759 42303 771
rect 42515 947 42675 959
rect 42515 771 42521 947
rect 42555 771 42635 947
rect 42669 771 42675 947
rect 42515 759 42675 771
rect 42887 947 43047 959
rect 42887 771 42893 947
rect 42927 771 43007 947
rect 43041 771 43047 947
rect 42887 759 43047 771
rect 43259 947 43419 959
rect 43259 771 43265 947
rect 43299 771 43379 947
rect 43413 771 43419 947
rect 43259 759 43419 771
rect 43631 947 43791 959
rect 43631 771 43637 947
rect 43671 771 43751 947
rect 43785 771 43791 947
rect 43631 759 43791 771
rect 44003 947 44163 959
rect 44003 771 44009 947
rect 44043 771 44123 947
rect 44157 771 44163 947
rect 44003 759 44163 771
rect 44375 947 44535 959
rect 44375 771 44381 947
rect 44415 771 44495 947
rect 44529 771 44535 947
rect 44375 759 44535 771
rect 44747 947 44907 959
rect 44747 771 44753 947
rect 44787 771 44867 947
rect 44901 771 44907 947
rect 44747 759 44907 771
rect 45119 947 45279 959
rect 45119 771 45125 947
rect 45159 771 45239 947
rect 45273 771 45279 947
rect 45119 759 45279 771
rect 45491 947 45651 959
rect 45491 771 45497 947
rect 45531 771 45611 947
rect 45645 771 45651 947
rect 45491 759 45651 771
rect 45863 947 46023 959
rect 45863 771 45869 947
rect 45903 771 45983 947
rect 46017 771 46023 947
rect 45863 759 46023 771
rect 46235 947 46395 959
rect 46235 771 46241 947
rect 46275 771 46355 947
rect 46389 771 46395 947
rect 46235 759 46395 771
rect 46607 947 46767 959
rect 46607 771 46613 947
rect 46647 771 46727 947
rect 46761 771 46767 947
rect 46607 759 46767 771
rect 46979 947 47139 959
rect 46979 771 46985 947
rect 47019 771 47099 947
rect 47133 771 47139 947
rect 46979 759 47139 771
rect 47351 947 47511 959
rect 47351 771 47357 947
rect 47391 771 47471 947
rect 47505 771 47511 947
rect 47351 759 47511 771
rect 47723 947 47883 959
rect 47723 771 47729 947
rect 47763 771 47843 947
rect 47877 771 47883 947
rect 47723 759 47883 771
rect 48095 947 48255 959
rect 48095 771 48101 947
rect 48135 771 48215 947
rect 48249 771 48255 947
rect 48095 759 48255 771
rect 48467 947 48627 959
rect 48467 771 48473 947
rect 48507 771 48587 947
rect 48621 771 48627 947
rect 48467 759 48627 771
rect 48839 947 48999 959
rect 48839 771 48845 947
rect 48879 771 48959 947
rect 48993 771 48999 947
rect 48839 759 48999 771
rect 49211 947 49371 959
rect 49211 771 49217 947
rect 49251 771 49331 947
rect 49365 771 49371 947
rect 49211 759 49371 771
rect 49583 947 49678 959
rect 49583 771 49589 947
rect 49623 771 49678 947
rect 49583 759 49678 771
rect 40720 541 40794 759
rect 41072 728 41142 759
rect 40824 722 41390 728
rect 40824 578 40836 722
rect 41006 578 41208 722
rect 41378 578 41390 722
rect 40824 572 41390 578
rect 41072 541 41142 572
rect 41444 541 41514 759
rect 41569 722 41761 727
rect 41569 681 41580 722
rect 41570 619 41580 681
rect 41569 578 41580 619
rect 41750 681 41761 722
rect 41750 619 41760 681
rect 41750 578 41761 619
rect 41569 573 41761 578
rect 41816 541 41886 759
rect 41941 722 42133 727
rect 41941 681 41952 722
rect 41942 619 41952 681
rect 41941 578 41952 619
rect 42122 681 42133 722
rect 42122 619 42132 681
rect 42122 578 42133 619
rect 41941 573 42133 578
rect 42188 541 42258 759
rect 42313 722 42505 727
rect 42313 681 42324 722
rect 42314 619 42324 681
rect 42313 578 42324 619
rect 42494 681 42505 722
rect 42494 619 42504 681
rect 42494 578 42505 619
rect 42313 573 42505 578
rect 42560 541 42630 759
rect 42685 722 42877 727
rect 42685 681 42696 722
rect 42686 619 42696 681
rect 42685 578 42696 619
rect 42866 681 42877 722
rect 42866 619 42876 681
rect 42866 578 42877 619
rect 42685 573 42877 578
rect 42932 541 43002 759
rect 43304 728 43374 759
rect 43056 722 43622 728
rect 43056 578 43068 722
rect 43238 578 43440 722
rect 43610 578 43622 722
rect 43056 572 43622 578
rect 43304 541 43374 572
rect 43676 541 43746 759
rect 43801 722 43993 727
rect 43801 681 43812 722
rect 43802 619 43812 681
rect 43801 578 43812 619
rect 43982 681 43993 722
rect 43982 619 43992 681
rect 43982 578 43993 619
rect 43801 573 43993 578
rect 44048 541 44118 759
rect 44173 722 44365 727
rect 44173 681 44184 722
rect 44174 619 44184 681
rect 44173 578 44184 619
rect 44354 681 44365 722
rect 44354 619 44364 681
rect 44354 578 44365 619
rect 44173 573 44365 578
rect 44420 541 44490 759
rect 44545 722 44737 727
rect 44545 681 44556 722
rect 44546 619 44556 681
rect 44545 578 44556 619
rect 44726 681 44737 722
rect 44726 619 44736 681
rect 44726 578 44737 619
rect 44545 573 44737 578
rect 44792 541 44862 759
rect 44917 722 45109 727
rect 44917 681 44928 722
rect 44918 619 44928 681
rect 44917 578 44928 619
rect 45098 681 45109 722
rect 45098 619 45108 681
rect 45098 578 45109 619
rect 44917 573 45109 578
rect 45164 541 45234 759
rect 45289 722 45481 727
rect 45289 681 45300 722
rect 45290 619 45300 681
rect 45289 578 45300 619
rect 45470 681 45481 722
rect 45470 619 45480 681
rect 45470 578 45481 619
rect 45289 573 45481 578
rect 45536 541 45606 759
rect 45661 722 45853 727
rect 45661 681 45672 722
rect 45662 619 45672 681
rect 45661 578 45672 619
rect 45842 681 45853 722
rect 45842 619 45852 681
rect 45842 578 45853 619
rect 45661 573 45853 578
rect 45908 541 45978 759
rect 46033 722 46225 727
rect 46033 681 46044 722
rect 46034 619 46044 681
rect 46033 578 46044 619
rect 46214 681 46225 722
rect 46214 619 46224 681
rect 46214 578 46225 619
rect 46033 573 46225 578
rect 46280 541 46350 759
rect 46405 722 46597 727
rect 46405 681 46416 722
rect 46406 619 46416 681
rect 46405 578 46416 619
rect 46586 681 46597 722
rect 46586 619 46596 681
rect 46586 578 46597 619
rect 46405 573 46597 578
rect 46652 541 46722 759
rect 46777 722 46969 727
rect 46777 681 46788 722
rect 46778 619 46788 681
rect 46777 578 46788 619
rect 46958 681 46969 722
rect 46958 619 46968 681
rect 46958 578 46969 619
rect 46777 573 46969 578
rect 47024 541 47094 759
rect 47149 722 47341 727
rect 47149 681 47160 722
rect 47150 619 47160 681
rect 47149 578 47160 619
rect 47330 681 47341 722
rect 47330 619 47340 681
rect 47330 578 47341 619
rect 47149 573 47341 578
rect 47396 541 47466 759
rect 47521 722 47713 727
rect 47521 681 47532 722
rect 47522 619 47532 681
rect 47521 578 47532 619
rect 47702 681 47713 722
rect 47702 619 47712 681
rect 47702 578 47713 619
rect 47521 573 47713 578
rect 47768 541 47838 759
rect 47893 722 48085 727
rect 47893 681 47904 722
rect 47894 619 47904 681
rect 47893 578 47904 619
rect 48074 681 48085 722
rect 48074 619 48084 681
rect 48074 578 48085 619
rect 47893 573 48085 578
rect 48140 541 48210 759
rect 48265 722 48457 727
rect 48265 681 48276 722
rect 48266 619 48276 681
rect 48265 578 48276 619
rect 48446 681 48457 722
rect 48446 619 48456 681
rect 48446 578 48457 619
rect 48265 573 48457 578
rect 48512 541 48582 759
rect 48637 722 48829 727
rect 48637 681 48648 722
rect 48638 619 48648 681
rect 48637 578 48648 619
rect 48818 681 48829 722
rect 48818 619 48828 681
rect 48818 578 48829 619
rect 48637 573 48829 578
rect 48884 541 48954 759
rect 49009 722 49201 727
rect 49009 681 49020 722
rect 49010 619 49020 681
rect 49009 578 49020 619
rect 49190 681 49201 722
rect 49190 619 49200 681
rect 49190 578 49201 619
rect 49009 573 49201 578
rect 49256 541 49326 759
rect 49381 722 49573 727
rect 49381 681 49392 722
rect 49382 619 49392 681
rect 49381 578 49392 619
rect 49562 681 49573 722
rect 49562 619 49572 681
rect 49562 578 49573 619
rect 49381 573 49573 578
rect 49604 541 49678 759
rect 40720 529 40815 541
rect 40720 353 40775 529
rect 40809 353 40815 529
rect 40720 341 40815 353
rect 41027 529 41187 541
rect 41027 353 41033 529
rect 41067 353 41147 529
rect 41181 353 41187 529
rect 41027 341 41187 353
rect 41399 529 41559 541
rect 41399 353 41405 529
rect 41439 353 41519 529
rect 41553 353 41559 529
rect 41399 341 41559 353
rect 41771 529 41931 541
rect 41771 353 41777 529
rect 41811 353 41891 529
rect 41925 353 41931 529
rect 41771 341 41931 353
rect 42143 529 42303 541
rect 42143 353 42149 529
rect 42183 353 42263 529
rect 42297 353 42303 529
rect 42143 341 42303 353
rect 42515 529 42675 541
rect 42515 353 42521 529
rect 42555 353 42635 529
rect 42669 353 42675 529
rect 42515 341 42675 353
rect 42887 529 43047 541
rect 42887 353 42893 529
rect 42927 353 43007 529
rect 43041 353 43047 529
rect 42887 341 43047 353
rect 43259 529 43419 541
rect 43259 353 43265 529
rect 43299 353 43379 529
rect 43413 353 43419 529
rect 43259 341 43419 353
rect 43631 529 43791 541
rect 43631 353 43637 529
rect 43671 353 43751 529
rect 43785 353 43791 529
rect 43631 341 43791 353
rect 44003 529 44163 541
rect 44003 353 44009 529
rect 44043 353 44123 529
rect 44157 353 44163 529
rect 44003 341 44163 353
rect 44375 529 44535 541
rect 44375 353 44381 529
rect 44415 353 44495 529
rect 44529 353 44535 529
rect 44375 341 44535 353
rect 44747 529 44907 541
rect 44747 353 44753 529
rect 44787 353 44867 529
rect 44901 353 44907 529
rect 44747 341 44907 353
rect 45119 529 45279 541
rect 45119 353 45125 529
rect 45159 353 45239 529
rect 45273 353 45279 529
rect 45119 341 45279 353
rect 45491 529 45651 541
rect 45491 353 45497 529
rect 45531 353 45611 529
rect 45645 353 45651 529
rect 45491 341 45651 353
rect 45863 529 46023 541
rect 45863 353 45869 529
rect 45903 353 45983 529
rect 46017 353 46023 529
rect 45863 341 46023 353
rect 46235 529 46395 541
rect 46235 353 46241 529
rect 46275 353 46355 529
rect 46389 353 46395 529
rect 46235 341 46395 353
rect 46607 529 46767 541
rect 46607 353 46613 529
rect 46647 353 46727 529
rect 46761 353 46767 529
rect 46607 341 46767 353
rect 46979 529 47139 541
rect 46979 353 46985 529
rect 47019 353 47099 529
rect 47133 353 47139 529
rect 46979 341 47139 353
rect 47351 529 47511 541
rect 47351 353 47357 529
rect 47391 353 47471 529
rect 47505 353 47511 529
rect 47351 341 47511 353
rect 47723 529 47883 541
rect 47723 353 47729 529
rect 47763 353 47843 529
rect 47877 353 47883 529
rect 47723 341 47883 353
rect 48095 529 48255 541
rect 48095 353 48101 529
rect 48135 353 48215 529
rect 48249 353 48255 529
rect 48095 341 48255 353
rect 48467 529 48627 541
rect 48467 353 48473 529
rect 48507 353 48587 529
rect 48621 353 48627 529
rect 48467 341 48627 353
rect 48839 529 48999 541
rect 48839 353 48845 529
rect 48879 353 48959 529
rect 48993 353 48999 529
rect 48839 341 48999 353
rect 49211 529 49371 541
rect 49211 353 49217 529
rect 49251 353 49331 529
rect 49365 353 49371 529
rect 49211 341 49371 353
rect 49583 529 49678 541
rect 49583 353 49589 529
rect 49623 353 49678 529
rect 49583 341 49678 353
rect 40720 218 40794 341
rect 40826 309 40836 314
rect 40825 304 40836 309
rect 40824 258 40836 304
rect 41006 309 41016 314
rect 41006 304 41017 309
rect 41072 304 41142 341
rect 41444 340 41514 341
rect 41816 340 41886 341
rect 42188 340 42258 341
rect 42560 340 42630 341
rect 42932 340 43002 341
rect 41198 309 41208 314
rect 41197 304 41208 309
rect 41006 258 41208 304
rect 41378 309 41388 314
rect 41378 304 41389 309
rect 41378 258 41390 304
rect 40824 246 41390 258
rect 41450 226 41508 340
rect 41570 309 41580 314
rect 41569 263 41580 309
rect 41750 309 41760 314
rect 41942 309 41952 314
rect 41570 258 41580 263
rect 41750 263 41761 309
rect 41941 263 41952 309
rect 42122 309 42132 314
rect 41750 258 41760 263
rect 41942 258 41952 263
rect 42122 263 42133 309
rect 42122 258 42132 263
rect 42194 226 42252 340
rect 42314 309 42324 314
rect 42313 263 42324 309
rect 42494 309 42504 314
rect 42686 309 42696 314
rect 42314 258 42324 263
rect 42494 263 42505 309
rect 42685 263 42696 309
rect 42866 309 42876 314
rect 42494 258 42504 263
rect 42686 258 42696 263
rect 42866 263 42877 309
rect 42866 258 42876 263
rect 42938 226 42996 340
rect 43058 309 43068 314
rect 43057 304 43068 309
rect 43056 258 43068 304
rect 43238 309 43248 314
rect 43238 304 43249 309
rect 43304 304 43374 341
rect 43676 340 43746 341
rect 44048 340 44118 341
rect 44420 340 44490 341
rect 44792 340 44862 341
rect 45164 340 45234 341
rect 45536 340 45606 341
rect 45908 340 45978 341
rect 46280 340 46350 341
rect 46652 340 46722 341
rect 47024 340 47094 341
rect 47396 340 47466 341
rect 47768 340 47838 341
rect 48140 340 48210 341
rect 48512 340 48582 341
rect 48884 340 48954 341
rect 49256 340 49326 341
rect 43430 309 43440 314
rect 43429 304 43440 309
rect 43238 258 43440 304
rect 43610 309 43620 314
rect 43610 304 43621 309
rect 43610 258 43622 304
rect 43056 246 43622 258
rect 43682 226 43740 340
rect 43802 309 43812 314
rect 43801 263 43812 309
rect 43982 309 43992 314
rect 44174 309 44184 314
rect 43802 258 43812 263
rect 43982 263 43993 309
rect 44173 263 44184 309
rect 44354 309 44364 314
rect 43982 258 43992 263
rect 44174 258 44184 263
rect 44354 263 44365 309
rect 44354 258 44364 263
rect 44426 226 44484 340
rect 44546 309 44556 314
rect 44545 263 44556 309
rect 44726 309 44736 314
rect 44918 309 44928 314
rect 44546 258 44556 263
rect 44726 263 44737 309
rect 44917 263 44928 309
rect 45098 309 45108 314
rect 44726 258 44736 263
rect 44918 258 44928 263
rect 45098 263 45109 309
rect 45098 258 45108 263
rect 45170 226 45228 340
rect 45290 309 45300 314
rect 45289 263 45300 309
rect 45470 309 45480 314
rect 45662 309 45672 314
rect 45290 258 45300 263
rect 45470 263 45481 309
rect 45661 263 45672 309
rect 45842 309 45852 314
rect 45470 258 45480 263
rect 45662 258 45672 263
rect 45842 263 45853 309
rect 45842 258 45852 263
rect 45914 226 45972 340
rect 46034 309 46044 314
rect 46033 263 46044 309
rect 46214 309 46224 314
rect 46406 309 46416 314
rect 46034 258 46044 263
rect 46214 263 46225 309
rect 46405 263 46416 309
rect 46586 309 46596 314
rect 46214 258 46224 263
rect 46406 258 46416 263
rect 46586 263 46597 309
rect 46586 258 46596 263
rect 46658 226 46716 340
rect 46778 309 46788 314
rect 46777 263 46788 309
rect 46958 309 46968 314
rect 47150 309 47160 314
rect 46778 258 46788 263
rect 46958 263 46969 309
rect 47149 263 47160 309
rect 47330 309 47340 314
rect 46958 258 46968 263
rect 47150 258 47160 263
rect 47330 263 47341 309
rect 47330 258 47340 263
rect 47402 226 47460 340
rect 47522 309 47532 314
rect 47521 263 47532 309
rect 47702 309 47712 314
rect 47894 309 47904 314
rect 47522 258 47532 263
rect 47702 263 47713 309
rect 47893 263 47904 309
rect 48074 309 48084 314
rect 47702 258 47712 263
rect 47894 258 47904 263
rect 48074 263 48085 309
rect 48074 258 48084 263
rect 48146 226 48204 340
rect 48266 309 48276 314
rect 48265 263 48276 309
rect 48446 309 48456 314
rect 48638 309 48648 314
rect 48266 258 48276 263
rect 48446 263 48457 309
rect 48637 263 48648 309
rect 48818 309 48828 314
rect 48446 258 48456 263
rect 48638 258 48648 263
rect 48818 263 48829 309
rect 48818 258 48828 263
rect 48890 226 48948 340
rect 49010 309 49020 314
rect 49009 263 49020 309
rect 49190 309 49200 314
rect 49382 309 49392 314
rect 49010 258 49020 263
rect 49190 263 49201 309
rect 49381 263 49392 309
rect 49562 309 49572 314
rect 49190 258 49200 263
rect 49382 258 49392 263
rect 49562 263 49573 309
rect 49562 258 49572 263
rect 41432 220 41526 226
rect 40720 212 40858 218
rect 40720 142 40776 212
rect 40846 142 40858 212
rect 41432 150 41444 220
rect 41514 150 41526 220
rect 41432 144 41526 150
rect 42176 220 42270 226
rect 42176 150 42188 220
rect 42258 150 42270 220
rect 42176 144 42270 150
rect 42920 220 43014 226
rect 42920 150 42932 220
rect 43002 150 43014 220
rect 42920 144 43014 150
rect 43664 220 43758 226
rect 43664 150 43676 220
rect 43746 150 43758 220
rect 43664 144 43758 150
rect 44408 220 44502 226
rect 44408 150 44420 220
rect 44490 150 44502 220
rect 44408 144 44502 150
rect 45152 220 45246 226
rect 45152 150 45164 220
rect 45234 150 45246 220
rect 45152 144 45246 150
rect 45896 220 45990 226
rect 45896 150 45908 220
rect 45978 150 45990 220
rect 45896 144 45990 150
rect 46640 220 46734 226
rect 46640 150 46652 220
rect 46722 150 46734 220
rect 46640 144 46734 150
rect 47384 220 47478 226
rect 47384 150 47396 220
rect 47466 150 47478 220
rect 47384 144 47478 150
rect 48128 220 48222 226
rect 48128 150 48140 220
rect 48210 150 48222 220
rect 48128 144 48222 150
rect 48872 220 48966 226
rect 49604 222 49678 341
rect 48872 150 48884 220
rect 48954 150 48966 220
rect 48872 144 48966 150
rect 49534 216 49678 222
rect 49534 146 49546 216
rect 49616 146 49678 216
rect 40720 136 40858 142
rect 40720 104 40794 136
rect 41450 104 41508 144
rect 42194 104 42252 144
rect 42938 104 42996 144
rect 43682 104 43740 144
rect 44426 104 44484 144
rect 45170 104 45228 144
rect 45914 104 45972 144
rect 46658 104 46716 144
rect 47402 104 47460 144
rect 48146 104 48204 144
rect 48890 104 48948 144
rect 49534 140 49678 146
rect 49604 116 49678 140
rect 49604 104 49692 116
rect 40646 -96 40656 104
rect 40856 -96 40866 104
rect 41370 -96 41380 104
rect 41580 -96 41590 104
rect 42114 -96 42124 104
rect 42324 -96 42334 104
rect 42858 -96 42868 104
rect 43068 -96 43078 104
rect 43602 -96 43612 104
rect 43812 -96 43822 104
rect 44346 -96 44356 104
rect 44556 -96 44566 104
rect 45090 -96 45100 104
rect 45300 -96 45310 104
rect 45834 -96 45844 104
rect 46044 -96 46054 104
rect 46578 -96 46588 104
rect 46788 -96 46798 104
rect 47322 -96 47332 104
rect 47532 -96 47542 104
rect 48066 -96 48076 104
rect 48276 -96 48286 104
rect 48810 -96 48820 104
rect 49020 -96 49030 104
rect 49554 -96 49564 104
rect 49764 -96 49774 104
<< via1 >>
rect 40656 19761 40856 19961
rect 41380 19761 41580 19961
rect 42124 19761 42324 19961
rect 42868 19761 43068 19961
rect 43612 19761 43812 19961
rect 44356 19761 44556 19961
rect 45100 19761 45300 19961
rect 45844 19761 46044 19961
rect 46588 19761 46788 19961
rect 47332 19761 47532 19961
rect 48076 19761 48276 19961
rect 48820 19761 49020 19961
rect 49564 19761 49764 19961
rect 40836 19596 41006 19607
rect 40836 19562 40837 19596
rect 40837 19562 41005 19596
rect 41005 19562 41006 19596
rect 40836 19551 41006 19562
rect 41208 19596 41378 19607
rect 41208 19562 41209 19596
rect 41209 19562 41377 19596
rect 41377 19562 41378 19596
rect 41208 19551 41378 19562
rect 41580 19596 41750 19607
rect 41580 19562 41581 19596
rect 41581 19562 41749 19596
rect 41749 19562 41750 19596
rect 41580 19551 41750 19562
rect 41952 19596 42122 19607
rect 41952 19562 41953 19596
rect 41953 19562 42121 19596
rect 42121 19562 42122 19596
rect 41952 19551 42122 19562
rect 42324 19596 42494 19607
rect 42324 19562 42325 19596
rect 42325 19562 42493 19596
rect 42493 19562 42494 19596
rect 42324 19551 42494 19562
rect 42696 19596 42866 19607
rect 42696 19562 42697 19596
rect 42697 19562 42865 19596
rect 42865 19562 42866 19596
rect 42696 19551 42866 19562
rect 43068 19596 43238 19607
rect 43068 19562 43069 19596
rect 43069 19562 43237 19596
rect 43237 19562 43238 19596
rect 43068 19551 43238 19562
rect 43440 19596 43610 19607
rect 43440 19562 43441 19596
rect 43441 19562 43609 19596
rect 43609 19562 43610 19596
rect 43440 19551 43610 19562
rect 43812 19596 43982 19607
rect 43812 19562 43813 19596
rect 43813 19562 43981 19596
rect 43981 19562 43982 19596
rect 43812 19551 43982 19562
rect 44184 19596 44354 19607
rect 44184 19562 44185 19596
rect 44185 19562 44353 19596
rect 44353 19562 44354 19596
rect 44184 19551 44354 19562
rect 44556 19596 44726 19607
rect 44556 19562 44557 19596
rect 44557 19562 44725 19596
rect 44725 19562 44726 19596
rect 44556 19551 44726 19562
rect 44928 19596 45098 19607
rect 44928 19562 44929 19596
rect 44929 19562 45097 19596
rect 45097 19562 45098 19596
rect 44928 19551 45098 19562
rect 45300 19596 45470 19607
rect 45300 19562 45301 19596
rect 45301 19562 45469 19596
rect 45469 19562 45470 19596
rect 45300 19551 45470 19562
rect 45672 19596 45842 19607
rect 45672 19562 45673 19596
rect 45673 19562 45841 19596
rect 45841 19562 45842 19596
rect 45672 19551 45842 19562
rect 46044 19596 46214 19607
rect 46044 19562 46045 19596
rect 46045 19562 46213 19596
rect 46213 19562 46214 19596
rect 46044 19551 46214 19562
rect 46416 19596 46586 19607
rect 46416 19562 46417 19596
rect 46417 19562 46585 19596
rect 46585 19562 46586 19596
rect 46416 19551 46586 19562
rect 46788 19596 46958 19607
rect 46788 19562 46789 19596
rect 46789 19562 46957 19596
rect 46957 19562 46958 19596
rect 46788 19551 46958 19562
rect 47160 19596 47330 19607
rect 47160 19562 47161 19596
rect 47161 19562 47329 19596
rect 47329 19562 47330 19596
rect 47160 19551 47330 19562
rect 47532 19596 47702 19607
rect 47532 19562 47533 19596
rect 47533 19562 47701 19596
rect 47701 19562 47702 19596
rect 47532 19551 47702 19562
rect 47904 19596 48074 19607
rect 47904 19562 47905 19596
rect 47905 19562 48073 19596
rect 48073 19562 48074 19596
rect 47904 19551 48074 19562
rect 48276 19596 48446 19607
rect 48276 19562 48277 19596
rect 48277 19562 48445 19596
rect 48445 19562 48446 19596
rect 48276 19551 48446 19562
rect 48648 19596 48818 19607
rect 48648 19562 48649 19596
rect 48649 19562 48817 19596
rect 48817 19562 48818 19596
rect 48648 19551 48818 19562
rect 49020 19596 49190 19607
rect 49020 19562 49021 19596
rect 49021 19562 49189 19596
rect 49189 19562 49190 19596
rect 49020 19551 49190 19562
rect 49392 19596 49562 19607
rect 49392 19562 49393 19596
rect 49393 19562 49561 19596
rect 49561 19562 49562 19596
rect 49392 19551 49562 19562
rect 40836 19286 41006 19287
rect 40836 19252 40837 19286
rect 40837 19252 41005 19286
rect 41005 19252 41006 19286
rect 40836 19178 41006 19252
rect 40836 19144 40837 19178
rect 40837 19144 41005 19178
rect 41005 19144 41006 19178
rect 40836 19143 41006 19144
rect 41208 19286 41378 19287
rect 41208 19252 41209 19286
rect 41209 19252 41377 19286
rect 41377 19252 41378 19286
rect 41208 19178 41378 19252
rect 41208 19144 41209 19178
rect 41209 19144 41377 19178
rect 41377 19144 41378 19178
rect 41208 19143 41378 19144
rect 41580 19286 41750 19287
rect 41580 19252 41581 19286
rect 41581 19252 41749 19286
rect 41749 19252 41750 19286
rect 41580 19178 41750 19252
rect 41580 19144 41581 19178
rect 41581 19144 41749 19178
rect 41749 19144 41750 19178
rect 41580 19143 41750 19144
rect 41952 19286 42122 19287
rect 41952 19252 41953 19286
rect 41953 19252 42121 19286
rect 42121 19252 42122 19286
rect 41952 19178 42122 19252
rect 41952 19144 41953 19178
rect 41953 19144 42121 19178
rect 42121 19144 42122 19178
rect 41952 19143 42122 19144
rect 42324 19286 42494 19287
rect 42324 19252 42325 19286
rect 42325 19252 42493 19286
rect 42493 19252 42494 19286
rect 42324 19178 42494 19252
rect 42324 19144 42325 19178
rect 42325 19144 42493 19178
rect 42493 19144 42494 19178
rect 42324 19143 42494 19144
rect 42696 19286 42866 19287
rect 42696 19252 42697 19286
rect 42697 19252 42865 19286
rect 42865 19252 42866 19286
rect 42696 19178 42866 19252
rect 42696 19144 42697 19178
rect 42697 19144 42865 19178
rect 42865 19144 42866 19178
rect 42696 19143 42866 19144
rect 43068 19286 43238 19287
rect 43068 19252 43069 19286
rect 43069 19252 43237 19286
rect 43237 19252 43238 19286
rect 43068 19178 43238 19252
rect 43068 19144 43069 19178
rect 43069 19144 43237 19178
rect 43237 19144 43238 19178
rect 43068 19143 43238 19144
rect 43440 19286 43610 19287
rect 43440 19252 43441 19286
rect 43441 19252 43609 19286
rect 43609 19252 43610 19286
rect 43440 19178 43610 19252
rect 43440 19144 43441 19178
rect 43441 19144 43609 19178
rect 43609 19144 43610 19178
rect 43440 19143 43610 19144
rect 43812 19286 43982 19287
rect 43812 19252 43813 19286
rect 43813 19252 43981 19286
rect 43981 19252 43982 19286
rect 43812 19178 43982 19252
rect 43812 19144 43813 19178
rect 43813 19144 43981 19178
rect 43981 19144 43982 19178
rect 43812 19143 43982 19144
rect 44184 19286 44354 19287
rect 44184 19252 44185 19286
rect 44185 19252 44353 19286
rect 44353 19252 44354 19286
rect 44184 19178 44354 19252
rect 44184 19144 44185 19178
rect 44185 19144 44353 19178
rect 44353 19144 44354 19178
rect 44184 19143 44354 19144
rect 44556 19286 44726 19287
rect 44556 19252 44557 19286
rect 44557 19252 44725 19286
rect 44725 19252 44726 19286
rect 44556 19178 44726 19252
rect 44556 19144 44557 19178
rect 44557 19144 44725 19178
rect 44725 19144 44726 19178
rect 44556 19143 44726 19144
rect 44928 19286 45098 19287
rect 44928 19252 44929 19286
rect 44929 19252 45097 19286
rect 45097 19252 45098 19286
rect 44928 19178 45098 19252
rect 44928 19144 44929 19178
rect 44929 19144 45097 19178
rect 45097 19144 45098 19178
rect 44928 19143 45098 19144
rect 45300 19286 45470 19287
rect 45300 19252 45301 19286
rect 45301 19252 45469 19286
rect 45469 19252 45470 19286
rect 45300 19178 45470 19252
rect 45300 19144 45301 19178
rect 45301 19144 45469 19178
rect 45469 19144 45470 19178
rect 45300 19143 45470 19144
rect 45672 19286 45842 19287
rect 45672 19252 45673 19286
rect 45673 19252 45841 19286
rect 45841 19252 45842 19286
rect 45672 19178 45842 19252
rect 45672 19144 45673 19178
rect 45673 19144 45841 19178
rect 45841 19144 45842 19178
rect 45672 19143 45842 19144
rect 46044 19286 46214 19287
rect 46044 19252 46045 19286
rect 46045 19252 46213 19286
rect 46213 19252 46214 19286
rect 46044 19178 46214 19252
rect 46044 19144 46045 19178
rect 46045 19144 46213 19178
rect 46213 19144 46214 19178
rect 46044 19143 46214 19144
rect 46416 19286 46586 19287
rect 46416 19252 46417 19286
rect 46417 19252 46585 19286
rect 46585 19252 46586 19286
rect 46416 19178 46586 19252
rect 46416 19144 46417 19178
rect 46417 19144 46585 19178
rect 46585 19144 46586 19178
rect 46416 19143 46586 19144
rect 46788 19286 46958 19287
rect 46788 19252 46789 19286
rect 46789 19252 46957 19286
rect 46957 19252 46958 19286
rect 46788 19178 46958 19252
rect 46788 19144 46789 19178
rect 46789 19144 46957 19178
rect 46957 19144 46958 19178
rect 46788 19143 46958 19144
rect 47160 19286 47330 19287
rect 47160 19252 47161 19286
rect 47161 19252 47329 19286
rect 47329 19252 47330 19286
rect 47160 19178 47330 19252
rect 47160 19144 47161 19178
rect 47161 19144 47329 19178
rect 47329 19144 47330 19178
rect 47160 19143 47330 19144
rect 47532 19286 47702 19287
rect 47532 19252 47533 19286
rect 47533 19252 47701 19286
rect 47701 19252 47702 19286
rect 47532 19178 47702 19252
rect 47532 19144 47533 19178
rect 47533 19144 47701 19178
rect 47701 19144 47702 19178
rect 47532 19143 47702 19144
rect 47904 19286 48074 19287
rect 47904 19252 47905 19286
rect 47905 19252 48073 19286
rect 48073 19252 48074 19286
rect 47904 19178 48074 19252
rect 47904 19144 47905 19178
rect 47905 19144 48073 19178
rect 48073 19144 48074 19178
rect 47904 19143 48074 19144
rect 48276 19286 48446 19287
rect 48276 19252 48277 19286
rect 48277 19252 48445 19286
rect 48445 19252 48446 19286
rect 48276 19178 48446 19252
rect 48276 19144 48277 19178
rect 48277 19144 48445 19178
rect 48445 19144 48446 19178
rect 48276 19143 48446 19144
rect 48648 19286 48818 19287
rect 48648 19252 48649 19286
rect 48649 19252 48817 19286
rect 48817 19252 48818 19286
rect 48648 19178 48818 19252
rect 48648 19144 48649 19178
rect 48649 19144 48817 19178
rect 48817 19144 48818 19178
rect 48648 19143 48818 19144
rect 49020 19286 49190 19287
rect 49020 19252 49021 19286
rect 49021 19252 49189 19286
rect 49189 19252 49190 19286
rect 49020 19178 49190 19252
rect 49020 19144 49021 19178
rect 49021 19144 49189 19178
rect 49189 19144 49190 19178
rect 49020 19143 49190 19144
rect 49392 19286 49562 19287
rect 49392 19252 49393 19286
rect 49393 19252 49561 19286
rect 49561 19252 49562 19286
rect 49392 19178 49562 19252
rect 49392 19144 49393 19178
rect 49393 19144 49561 19178
rect 49561 19144 49562 19178
rect 49392 19143 49562 19144
rect 40836 18868 41006 18869
rect 40836 18834 40837 18868
rect 40837 18834 41005 18868
rect 41005 18834 41006 18868
rect 40836 18760 41006 18834
rect 40836 18726 40837 18760
rect 40837 18726 41005 18760
rect 41005 18726 41006 18760
rect 40836 18725 41006 18726
rect 41208 18868 41378 18869
rect 41208 18834 41209 18868
rect 41209 18834 41377 18868
rect 41377 18834 41378 18868
rect 41208 18760 41378 18834
rect 41208 18726 41209 18760
rect 41209 18726 41377 18760
rect 41377 18726 41378 18760
rect 41208 18725 41378 18726
rect 41580 18868 41750 18869
rect 41580 18834 41581 18868
rect 41581 18834 41749 18868
rect 41749 18834 41750 18868
rect 41580 18760 41750 18834
rect 41580 18726 41581 18760
rect 41581 18726 41749 18760
rect 41749 18726 41750 18760
rect 41580 18725 41750 18726
rect 41952 18868 42122 18869
rect 41952 18834 41953 18868
rect 41953 18834 42121 18868
rect 42121 18834 42122 18868
rect 41952 18760 42122 18834
rect 41952 18726 41953 18760
rect 41953 18726 42121 18760
rect 42121 18726 42122 18760
rect 41952 18725 42122 18726
rect 42324 18868 42494 18869
rect 42324 18834 42325 18868
rect 42325 18834 42493 18868
rect 42493 18834 42494 18868
rect 42324 18760 42494 18834
rect 42324 18726 42325 18760
rect 42325 18726 42493 18760
rect 42493 18726 42494 18760
rect 42324 18725 42494 18726
rect 42696 18868 42866 18869
rect 42696 18834 42697 18868
rect 42697 18834 42865 18868
rect 42865 18834 42866 18868
rect 42696 18760 42866 18834
rect 42696 18726 42697 18760
rect 42697 18726 42865 18760
rect 42865 18726 42866 18760
rect 42696 18725 42866 18726
rect 43068 18868 43238 18869
rect 43068 18834 43069 18868
rect 43069 18834 43237 18868
rect 43237 18834 43238 18868
rect 43068 18760 43238 18834
rect 43068 18726 43069 18760
rect 43069 18726 43237 18760
rect 43237 18726 43238 18760
rect 43068 18725 43238 18726
rect 43440 18868 43610 18869
rect 43440 18834 43441 18868
rect 43441 18834 43609 18868
rect 43609 18834 43610 18868
rect 43440 18760 43610 18834
rect 43440 18726 43441 18760
rect 43441 18726 43609 18760
rect 43609 18726 43610 18760
rect 43440 18725 43610 18726
rect 43812 18868 43982 18869
rect 43812 18834 43813 18868
rect 43813 18834 43981 18868
rect 43981 18834 43982 18868
rect 43812 18760 43982 18834
rect 43812 18726 43813 18760
rect 43813 18726 43981 18760
rect 43981 18726 43982 18760
rect 43812 18725 43982 18726
rect 44184 18868 44354 18869
rect 44184 18834 44185 18868
rect 44185 18834 44353 18868
rect 44353 18834 44354 18868
rect 44184 18760 44354 18834
rect 44184 18726 44185 18760
rect 44185 18726 44353 18760
rect 44353 18726 44354 18760
rect 44184 18725 44354 18726
rect 44556 18868 44726 18869
rect 44556 18834 44557 18868
rect 44557 18834 44725 18868
rect 44725 18834 44726 18868
rect 44556 18760 44726 18834
rect 44556 18726 44557 18760
rect 44557 18726 44725 18760
rect 44725 18726 44726 18760
rect 44556 18725 44726 18726
rect 44928 18868 45098 18869
rect 44928 18834 44929 18868
rect 44929 18834 45097 18868
rect 45097 18834 45098 18868
rect 44928 18760 45098 18834
rect 44928 18726 44929 18760
rect 44929 18726 45097 18760
rect 45097 18726 45098 18760
rect 44928 18725 45098 18726
rect 45300 18868 45470 18869
rect 45300 18834 45301 18868
rect 45301 18834 45469 18868
rect 45469 18834 45470 18868
rect 45300 18760 45470 18834
rect 45300 18726 45301 18760
rect 45301 18726 45469 18760
rect 45469 18726 45470 18760
rect 45300 18725 45470 18726
rect 45672 18868 45842 18869
rect 45672 18834 45673 18868
rect 45673 18834 45841 18868
rect 45841 18834 45842 18868
rect 45672 18760 45842 18834
rect 45672 18726 45673 18760
rect 45673 18726 45841 18760
rect 45841 18726 45842 18760
rect 45672 18725 45842 18726
rect 46044 18868 46214 18869
rect 46044 18834 46045 18868
rect 46045 18834 46213 18868
rect 46213 18834 46214 18868
rect 46044 18760 46214 18834
rect 46044 18726 46045 18760
rect 46045 18726 46213 18760
rect 46213 18726 46214 18760
rect 46044 18725 46214 18726
rect 46416 18868 46586 18869
rect 46416 18834 46417 18868
rect 46417 18834 46585 18868
rect 46585 18834 46586 18868
rect 46416 18760 46586 18834
rect 46416 18726 46417 18760
rect 46417 18726 46585 18760
rect 46585 18726 46586 18760
rect 46416 18725 46586 18726
rect 46788 18868 46958 18869
rect 46788 18834 46789 18868
rect 46789 18834 46957 18868
rect 46957 18834 46958 18868
rect 46788 18760 46958 18834
rect 46788 18726 46789 18760
rect 46789 18726 46957 18760
rect 46957 18726 46958 18760
rect 46788 18725 46958 18726
rect 47160 18868 47330 18869
rect 47160 18834 47161 18868
rect 47161 18834 47329 18868
rect 47329 18834 47330 18868
rect 47160 18760 47330 18834
rect 47160 18726 47161 18760
rect 47161 18726 47329 18760
rect 47329 18726 47330 18760
rect 47160 18725 47330 18726
rect 47532 18868 47702 18869
rect 47532 18834 47533 18868
rect 47533 18834 47701 18868
rect 47701 18834 47702 18868
rect 47532 18760 47702 18834
rect 47532 18726 47533 18760
rect 47533 18726 47701 18760
rect 47701 18726 47702 18760
rect 47532 18725 47702 18726
rect 47904 18868 48074 18869
rect 47904 18834 47905 18868
rect 47905 18834 48073 18868
rect 48073 18834 48074 18868
rect 47904 18760 48074 18834
rect 47904 18726 47905 18760
rect 47905 18726 48073 18760
rect 48073 18726 48074 18760
rect 47904 18725 48074 18726
rect 48276 18868 48446 18869
rect 48276 18834 48277 18868
rect 48277 18834 48445 18868
rect 48445 18834 48446 18868
rect 48276 18760 48446 18834
rect 48276 18726 48277 18760
rect 48277 18726 48445 18760
rect 48445 18726 48446 18760
rect 48276 18725 48446 18726
rect 48648 18868 48818 18869
rect 48648 18834 48649 18868
rect 48649 18834 48817 18868
rect 48817 18834 48818 18868
rect 48648 18760 48818 18834
rect 48648 18726 48649 18760
rect 48649 18726 48817 18760
rect 48817 18726 48818 18760
rect 48648 18725 48818 18726
rect 49020 18868 49190 18869
rect 49020 18834 49021 18868
rect 49021 18834 49189 18868
rect 49189 18834 49190 18868
rect 49020 18760 49190 18834
rect 49020 18726 49021 18760
rect 49021 18726 49189 18760
rect 49189 18726 49190 18760
rect 49020 18725 49190 18726
rect 49392 18868 49562 18869
rect 49392 18834 49393 18868
rect 49393 18834 49561 18868
rect 49561 18834 49562 18868
rect 49392 18760 49562 18834
rect 49392 18726 49393 18760
rect 49393 18726 49561 18760
rect 49561 18726 49562 18760
rect 49392 18725 49562 18726
rect 40836 18450 41006 18451
rect 40836 18416 40837 18450
rect 40837 18416 41005 18450
rect 41005 18416 41006 18450
rect 40836 18342 41006 18416
rect 40836 18308 40837 18342
rect 40837 18308 41005 18342
rect 41005 18308 41006 18342
rect 40836 18307 41006 18308
rect 41208 18450 41378 18451
rect 41208 18416 41209 18450
rect 41209 18416 41377 18450
rect 41377 18416 41378 18450
rect 41208 18342 41378 18416
rect 41208 18308 41209 18342
rect 41209 18308 41377 18342
rect 41377 18308 41378 18342
rect 41208 18307 41378 18308
rect 41580 18450 41750 18451
rect 41580 18416 41581 18450
rect 41581 18416 41749 18450
rect 41749 18416 41750 18450
rect 41580 18342 41750 18416
rect 41580 18308 41581 18342
rect 41581 18308 41749 18342
rect 41749 18308 41750 18342
rect 41580 18307 41750 18308
rect 41952 18450 42122 18451
rect 41952 18416 41953 18450
rect 41953 18416 42121 18450
rect 42121 18416 42122 18450
rect 41952 18342 42122 18416
rect 41952 18308 41953 18342
rect 41953 18308 42121 18342
rect 42121 18308 42122 18342
rect 41952 18307 42122 18308
rect 42324 18450 42494 18451
rect 42324 18416 42325 18450
rect 42325 18416 42493 18450
rect 42493 18416 42494 18450
rect 42324 18342 42494 18416
rect 42324 18308 42325 18342
rect 42325 18308 42493 18342
rect 42493 18308 42494 18342
rect 42324 18307 42494 18308
rect 42696 18450 42866 18451
rect 42696 18416 42697 18450
rect 42697 18416 42865 18450
rect 42865 18416 42866 18450
rect 42696 18342 42866 18416
rect 42696 18308 42697 18342
rect 42697 18308 42865 18342
rect 42865 18308 42866 18342
rect 42696 18307 42866 18308
rect 43068 18450 43238 18451
rect 43068 18416 43069 18450
rect 43069 18416 43237 18450
rect 43237 18416 43238 18450
rect 43068 18342 43238 18416
rect 43068 18308 43069 18342
rect 43069 18308 43237 18342
rect 43237 18308 43238 18342
rect 43068 18307 43238 18308
rect 43440 18450 43610 18451
rect 43440 18416 43441 18450
rect 43441 18416 43609 18450
rect 43609 18416 43610 18450
rect 43440 18342 43610 18416
rect 43440 18308 43441 18342
rect 43441 18308 43609 18342
rect 43609 18308 43610 18342
rect 43440 18307 43610 18308
rect 43812 18450 43982 18451
rect 43812 18416 43813 18450
rect 43813 18416 43981 18450
rect 43981 18416 43982 18450
rect 43812 18342 43982 18416
rect 43812 18308 43813 18342
rect 43813 18308 43981 18342
rect 43981 18308 43982 18342
rect 43812 18307 43982 18308
rect 44184 18450 44354 18451
rect 44184 18416 44185 18450
rect 44185 18416 44353 18450
rect 44353 18416 44354 18450
rect 44184 18342 44354 18416
rect 44184 18308 44185 18342
rect 44185 18308 44353 18342
rect 44353 18308 44354 18342
rect 44184 18307 44354 18308
rect 44556 18450 44726 18451
rect 44556 18416 44557 18450
rect 44557 18416 44725 18450
rect 44725 18416 44726 18450
rect 44556 18342 44726 18416
rect 44556 18308 44557 18342
rect 44557 18308 44725 18342
rect 44725 18308 44726 18342
rect 44556 18307 44726 18308
rect 44928 18450 45098 18451
rect 44928 18416 44929 18450
rect 44929 18416 45097 18450
rect 45097 18416 45098 18450
rect 44928 18342 45098 18416
rect 44928 18308 44929 18342
rect 44929 18308 45097 18342
rect 45097 18308 45098 18342
rect 44928 18307 45098 18308
rect 45300 18450 45470 18451
rect 45300 18416 45301 18450
rect 45301 18416 45469 18450
rect 45469 18416 45470 18450
rect 45300 18342 45470 18416
rect 45300 18308 45301 18342
rect 45301 18308 45469 18342
rect 45469 18308 45470 18342
rect 45300 18307 45470 18308
rect 45672 18450 45842 18451
rect 45672 18416 45673 18450
rect 45673 18416 45841 18450
rect 45841 18416 45842 18450
rect 45672 18342 45842 18416
rect 45672 18308 45673 18342
rect 45673 18308 45841 18342
rect 45841 18308 45842 18342
rect 45672 18307 45842 18308
rect 46044 18450 46214 18451
rect 46044 18416 46045 18450
rect 46045 18416 46213 18450
rect 46213 18416 46214 18450
rect 46044 18342 46214 18416
rect 46044 18308 46045 18342
rect 46045 18308 46213 18342
rect 46213 18308 46214 18342
rect 46044 18307 46214 18308
rect 46416 18450 46586 18451
rect 46416 18416 46417 18450
rect 46417 18416 46585 18450
rect 46585 18416 46586 18450
rect 46416 18342 46586 18416
rect 46416 18308 46417 18342
rect 46417 18308 46585 18342
rect 46585 18308 46586 18342
rect 46416 18307 46586 18308
rect 46788 18450 46958 18451
rect 46788 18416 46789 18450
rect 46789 18416 46957 18450
rect 46957 18416 46958 18450
rect 46788 18342 46958 18416
rect 46788 18308 46789 18342
rect 46789 18308 46957 18342
rect 46957 18308 46958 18342
rect 46788 18307 46958 18308
rect 47160 18450 47330 18451
rect 47160 18416 47161 18450
rect 47161 18416 47329 18450
rect 47329 18416 47330 18450
rect 47160 18342 47330 18416
rect 47160 18308 47161 18342
rect 47161 18308 47329 18342
rect 47329 18308 47330 18342
rect 47160 18307 47330 18308
rect 47532 18450 47702 18451
rect 47532 18416 47533 18450
rect 47533 18416 47701 18450
rect 47701 18416 47702 18450
rect 47532 18342 47702 18416
rect 47532 18308 47533 18342
rect 47533 18308 47701 18342
rect 47701 18308 47702 18342
rect 47532 18307 47702 18308
rect 47904 18450 48074 18451
rect 47904 18416 47905 18450
rect 47905 18416 48073 18450
rect 48073 18416 48074 18450
rect 47904 18342 48074 18416
rect 47904 18308 47905 18342
rect 47905 18308 48073 18342
rect 48073 18308 48074 18342
rect 47904 18307 48074 18308
rect 48276 18450 48446 18451
rect 48276 18416 48277 18450
rect 48277 18416 48445 18450
rect 48445 18416 48446 18450
rect 48276 18342 48446 18416
rect 48276 18308 48277 18342
rect 48277 18308 48445 18342
rect 48445 18308 48446 18342
rect 48276 18307 48446 18308
rect 48648 18450 48818 18451
rect 48648 18416 48649 18450
rect 48649 18416 48817 18450
rect 48817 18416 48818 18450
rect 48648 18342 48818 18416
rect 48648 18308 48649 18342
rect 48649 18308 48817 18342
rect 48817 18308 48818 18342
rect 48648 18307 48818 18308
rect 49020 18450 49190 18451
rect 49020 18416 49021 18450
rect 49021 18416 49189 18450
rect 49189 18416 49190 18450
rect 49020 18342 49190 18416
rect 49020 18308 49021 18342
rect 49021 18308 49189 18342
rect 49189 18308 49190 18342
rect 49020 18307 49190 18308
rect 49392 18450 49562 18451
rect 49392 18416 49393 18450
rect 49393 18416 49561 18450
rect 49561 18416 49562 18450
rect 49392 18342 49562 18416
rect 49392 18308 49393 18342
rect 49393 18308 49561 18342
rect 49561 18308 49562 18342
rect 49392 18307 49562 18308
rect 40836 18032 41006 18043
rect 40836 17998 40837 18032
rect 40837 17998 41005 18032
rect 41005 17998 41006 18032
rect 40836 17987 41006 17998
rect 41208 18032 41378 18043
rect 41208 17998 41209 18032
rect 41209 17998 41377 18032
rect 41377 17998 41378 18032
rect 41208 17987 41378 17998
rect 41580 18032 41750 18043
rect 41580 17998 41581 18032
rect 41581 17998 41749 18032
rect 41749 17998 41750 18032
rect 41580 17987 41750 17998
rect 38314 17108 38800 17616
rect 40836 17374 41006 17383
rect 40836 17340 40837 17374
rect 40837 17340 41005 17374
rect 41005 17340 41006 17374
rect 40836 17329 41006 17340
rect 41952 18032 42122 18043
rect 41952 17998 41953 18032
rect 41953 17998 42121 18032
rect 42121 17998 42122 18032
rect 41952 17987 42122 17998
rect 42324 18032 42494 18043
rect 42324 17998 42325 18032
rect 42325 17998 42493 18032
rect 42493 17998 42494 18032
rect 42324 17987 42494 17998
rect 42696 18032 42866 18043
rect 42696 17998 42697 18032
rect 42697 17998 42865 18032
rect 42865 17998 42866 18032
rect 42696 17987 42866 17998
rect 43068 18032 43238 18043
rect 43068 17998 43069 18032
rect 43069 17998 43237 18032
rect 43237 17998 43238 18032
rect 43068 17987 43238 17998
rect 43440 18032 43610 18043
rect 43440 17998 43441 18032
rect 43441 17998 43609 18032
rect 43609 17998 43610 18032
rect 43440 17987 43610 17998
rect 43812 18032 43982 18043
rect 43812 17998 43813 18032
rect 43813 17998 43981 18032
rect 43981 17998 43982 18032
rect 43812 17987 43982 17998
rect 41816 17669 42630 17849
rect 41208 17374 41378 17383
rect 41208 17340 41209 17374
rect 41209 17340 41377 17374
rect 41377 17340 41378 17374
rect 41208 17329 41378 17340
rect 41580 17374 41750 17383
rect 41580 17340 41581 17374
rect 41581 17340 41749 17374
rect 41749 17340 41750 17374
rect 41580 17329 41750 17340
rect 41952 17374 42122 17383
rect 41952 17340 41953 17374
rect 41953 17340 42121 17374
rect 42121 17340 42122 17374
rect 41952 17329 42122 17340
rect 42324 17374 42494 17383
rect 42324 17340 42325 17374
rect 42325 17340 42493 17374
rect 42493 17340 42494 17374
rect 42324 17329 42494 17340
rect 42696 17374 42866 17383
rect 42696 17340 42697 17374
rect 42697 17340 42865 17374
rect 42865 17340 42866 17374
rect 42696 17329 42866 17340
rect 43068 17374 43238 17383
rect 43068 17340 43069 17374
rect 43069 17340 43237 17374
rect 43237 17340 43238 17374
rect 43068 17329 43238 17340
rect 44184 18032 44354 18043
rect 44184 17998 44185 18032
rect 44185 17998 44353 18032
rect 44353 17998 44354 18032
rect 44184 17987 44354 17998
rect 44556 18032 44726 18043
rect 44556 17998 44557 18032
rect 44557 17998 44725 18032
rect 44725 17998 44726 18032
rect 44556 17987 44726 17998
rect 44928 18032 45098 18043
rect 44928 17998 44929 18032
rect 44929 17998 45097 18032
rect 45097 17998 45098 18032
rect 44928 17987 45098 17998
rect 45300 18032 45470 18043
rect 45300 17998 45301 18032
rect 45301 17998 45469 18032
rect 45469 17998 45470 18032
rect 45300 17987 45470 17998
rect 45672 18032 45842 18043
rect 45672 17998 45673 18032
rect 45673 17998 45841 18032
rect 45841 17998 45842 18032
rect 45672 17987 45842 17998
rect 46044 18032 46214 18043
rect 46044 17998 46045 18032
rect 46045 17998 46213 18032
rect 46213 17998 46214 18032
rect 46044 17987 46214 17998
rect 45826 17541 46104 17815
rect 43440 17374 43610 17383
rect 43440 17340 43441 17374
rect 43441 17340 43609 17374
rect 43609 17340 43610 17374
rect 43440 17329 43610 17340
rect 43942 17253 44224 17525
rect 44686 17253 44968 17525
rect 45430 17253 45712 17525
rect 46416 18032 46586 18043
rect 46416 17998 46417 18032
rect 46417 17998 46585 18032
rect 46585 17998 46586 18032
rect 46416 17987 46586 17998
rect 46788 18032 46958 18043
rect 46788 17998 46789 18032
rect 46789 17998 46957 18032
rect 46957 17998 46958 18032
rect 46788 17987 46958 17998
rect 47160 18032 47330 18043
rect 47160 17998 47161 18032
rect 47161 17998 47329 18032
rect 47329 17998 47330 18032
rect 47160 17987 47330 17998
rect 47532 18032 47702 18043
rect 47532 17998 47533 18032
rect 47533 17998 47701 18032
rect 47701 17998 47702 18032
rect 47532 17987 47702 17998
rect 47904 18032 48074 18043
rect 47904 17998 47905 18032
rect 47905 17998 48073 18032
rect 48073 17998 48074 18032
rect 47904 17987 48074 17998
rect 48276 18032 48446 18043
rect 48276 17998 48277 18032
rect 48277 17998 48445 18032
rect 48445 17998 48446 18032
rect 48276 17987 48446 17998
rect 48648 18032 48818 18043
rect 48648 17998 48649 18032
rect 48649 17998 48817 18032
rect 48817 17998 48818 18032
rect 48648 17987 48818 17998
rect 49020 18032 49190 18043
rect 49020 17998 49021 18032
rect 49021 17998 49189 18032
rect 49189 17998 49190 18032
rect 49020 17987 49190 17998
rect 49392 18032 49562 18043
rect 49392 17998 49393 18032
rect 49393 17998 49561 18032
rect 49561 17998 49562 18032
rect 49392 17987 49562 17998
rect 40836 16446 41006 16447
rect 40836 16412 40837 16446
rect 40837 16412 41005 16446
rect 41005 16412 41006 16446
rect 40836 16338 41006 16412
rect 40836 16304 40837 16338
rect 40837 16304 41005 16338
rect 41005 16304 41006 16338
rect 40836 16303 41006 16304
rect 41208 16446 41378 16447
rect 41208 16412 41209 16446
rect 41209 16412 41377 16446
rect 41377 16412 41378 16446
rect 41208 16338 41378 16412
rect 41208 16304 41209 16338
rect 41209 16304 41377 16338
rect 41377 16304 41378 16338
rect 41208 16303 41378 16304
rect 41580 16446 41750 16447
rect 41580 16412 41581 16446
rect 41581 16412 41749 16446
rect 41749 16412 41750 16446
rect 41580 16338 41750 16412
rect 41580 16304 41581 16338
rect 41581 16304 41749 16338
rect 41749 16304 41750 16338
rect 41580 16303 41750 16304
rect 41952 16446 42122 16447
rect 41952 16412 41953 16446
rect 41953 16412 42121 16446
rect 42121 16412 42122 16446
rect 41952 16338 42122 16412
rect 41952 16304 41953 16338
rect 41953 16304 42121 16338
rect 42121 16304 42122 16338
rect 41952 16303 42122 16304
rect 42324 16446 42494 16447
rect 42324 16412 42325 16446
rect 42325 16412 42493 16446
rect 42493 16412 42494 16446
rect 42324 16338 42494 16412
rect 42324 16304 42325 16338
rect 42325 16304 42493 16338
rect 42493 16304 42494 16338
rect 42324 16303 42494 16304
rect 42696 16446 42866 16447
rect 42696 16412 42697 16446
rect 42697 16412 42865 16446
rect 42865 16412 42866 16446
rect 42696 16338 42866 16412
rect 42696 16304 42697 16338
rect 42697 16304 42865 16338
rect 42865 16304 42866 16338
rect 42696 16303 42866 16304
rect 43068 16446 43238 16447
rect 43068 16412 43069 16446
rect 43069 16412 43237 16446
rect 43237 16412 43238 16446
rect 43068 16338 43238 16412
rect 43068 16304 43069 16338
rect 43069 16304 43237 16338
rect 43237 16304 43238 16338
rect 43068 16303 43238 16304
rect 43440 16446 43610 16447
rect 43440 16412 43441 16446
rect 43441 16412 43609 16446
rect 43609 16412 43610 16446
rect 43440 16338 43610 16412
rect 43440 16304 43441 16338
rect 43441 16304 43609 16338
rect 43609 16304 43610 16338
rect 43440 16303 43610 16304
rect 45566 16304 45734 16470
rect 46174 17253 46456 17525
rect 46918 17253 47200 17525
rect 47662 17253 47944 17525
rect 48406 17253 48688 17525
rect 49150 17253 49432 17525
rect 45566 15904 45734 16070
rect 45566 15504 45734 15670
rect 40836 15410 41006 15411
rect 40836 15376 40837 15410
rect 40837 15376 41005 15410
rect 41005 15376 41006 15410
rect 40836 15302 41006 15376
rect 40836 15268 40837 15302
rect 40837 15268 41005 15302
rect 41005 15268 41006 15302
rect 40836 15267 41006 15268
rect 41208 15410 41378 15411
rect 41208 15376 41209 15410
rect 41209 15376 41377 15410
rect 41377 15376 41378 15410
rect 41208 15302 41378 15376
rect 41208 15268 41209 15302
rect 41209 15268 41377 15302
rect 41377 15268 41378 15302
rect 41208 15267 41378 15268
rect 41580 15410 41750 15411
rect 41580 15376 41581 15410
rect 41581 15376 41749 15410
rect 41749 15376 41750 15410
rect 41580 15302 41750 15376
rect 41580 15268 41581 15302
rect 41581 15268 41749 15302
rect 41749 15268 41750 15302
rect 41580 15267 41750 15268
rect 41952 15410 42122 15411
rect 41952 15376 41953 15410
rect 41953 15376 42121 15410
rect 42121 15376 42122 15410
rect 41952 15302 42122 15376
rect 41952 15268 41953 15302
rect 41953 15268 42121 15302
rect 42121 15268 42122 15302
rect 41952 15267 42122 15268
rect 42324 15410 42494 15411
rect 42324 15376 42325 15410
rect 42325 15376 42493 15410
rect 42493 15376 42494 15410
rect 42324 15302 42494 15376
rect 42324 15268 42325 15302
rect 42325 15268 42493 15302
rect 42493 15268 42494 15302
rect 42324 15267 42494 15268
rect 42696 15410 42866 15411
rect 42696 15376 42697 15410
rect 42697 15376 42865 15410
rect 42865 15376 42866 15410
rect 42696 15302 42866 15376
rect 42696 15268 42697 15302
rect 42697 15268 42865 15302
rect 42865 15268 42866 15302
rect 42696 15267 42866 15268
rect 43068 15410 43238 15411
rect 43068 15376 43069 15410
rect 43069 15376 43237 15410
rect 43237 15376 43238 15410
rect 43068 15302 43238 15376
rect 43068 15268 43069 15302
rect 43069 15268 43237 15302
rect 43237 15268 43238 15302
rect 43068 15267 43238 15268
rect 43440 15410 43610 15411
rect 43440 15376 43441 15410
rect 43441 15376 43609 15410
rect 43609 15376 43610 15410
rect 43440 15302 43610 15376
rect 43440 15268 43441 15302
rect 43441 15268 43609 15302
rect 43609 15268 43610 15302
rect 43440 15267 43610 15268
rect 45852 14845 46134 15117
rect 40836 14374 41006 14375
rect 40836 14340 40837 14374
rect 40837 14340 41005 14374
rect 41005 14340 41006 14374
rect 40836 14266 41006 14340
rect 40836 14232 40837 14266
rect 40837 14232 41005 14266
rect 41005 14232 41006 14266
rect 40836 14231 41006 14232
rect 41208 14374 41378 14375
rect 41208 14340 41209 14374
rect 41209 14340 41377 14374
rect 41377 14340 41378 14374
rect 41208 14266 41378 14340
rect 41208 14232 41209 14266
rect 41209 14232 41377 14266
rect 41377 14232 41378 14266
rect 41208 14231 41378 14232
rect 41580 14374 41750 14375
rect 41580 14340 41581 14374
rect 41581 14340 41749 14374
rect 41749 14340 41750 14374
rect 41580 14266 41750 14340
rect 41580 14232 41581 14266
rect 41581 14232 41749 14266
rect 41749 14232 41750 14266
rect 41580 14231 41750 14232
rect 41952 14374 42122 14375
rect 41952 14340 41953 14374
rect 41953 14340 42121 14374
rect 42121 14340 42122 14374
rect 41952 14266 42122 14340
rect 41952 14232 41953 14266
rect 41953 14232 42121 14266
rect 42121 14232 42122 14266
rect 41952 14231 42122 14232
rect 42324 14374 42494 14375
rect 42324 14340 42325 14374
rect 42325 14340 42493 14374
rect 42493 14340 42494 14374
rect 42324 14266 42494 14340
rect 42324 14232 42325 14266
rect 42325 14232 42493 14266
rect 42493 14232 42494 14266
rect 42324 14231 42494 14232
rect 42696 14374 42866 14375
rect 42696 14340 42697 14374
rect 42697 14340 42865 14374
rect 42865 14340 42866 14374
rect 42696 14266 42866 14340
rect 42696 14232 42697 14266
rect 42697 14232 42865 14266
rect 42865 14232 42866 14266
rect 42696 14231 42866 14232
rect 43068 14374 43238 14375
rect 43068 14340 43069 14374
rect 43069 14340 43237 14374
rect 43237 14340 43238 14374
rect 43068 14266 43238 14340
rect 43068 14232 43069 14266
rect 43069 14232 43237 14266
rect 43237 14232 43238 14266
rect 43068 14231 43238 14232
rect 43440 14374 43610 14375
rect 43440 14340 43441 14374
rect 43441 14340 43609 14374
rect 43609 14340 43610 14374
rect 43440 14266 43610 14340
rect 43440 14232 43441 14266
rect 43441 14232 43609 14266
rect 43609 14232 43610 14266
rect 43440 14231 43610 14232
rect 40836 13338 41006 13353
rect 40836 13304 40837 13338
rect 40837 13304 41005 13338
rect 41005 13304 41006 13338
rect 40836 13289 41006 13304
rect 41208 13338 41378 13353
rect 41208 13304 41209 13338
rect 41209 13304 41377 13338
rect 41377 13304 41378 13338
rect 41208 13289 41378 13304
rect 41580 13338 41750 13353
rect 41580 13304 41581 13338
rect 41581 13304 41749 13338
rect 41749 13304 41750 13338
rect 41580 13289 41750 13304
rect 41952 13338 42122 13353
rect 41952 13304 41953 13338
rect 41953 13304 42121 13338
rect 42121 13304 42122 13338
rect 41952 13289 42122 13304
rect 42324 13338 42494 13353
rect 42324 13304 42325 13338
rect 42325 13304 42493 13338
rect 42493 13304 42494 13338
rect 42324 13289 42494 13304
rect 42696 13338 42866 13353
rect 42696 13304 42697 13338
rect 42697 13304 42865 13338
rect 42865 13304 42866 13338
rect 42696 13289 42866 13304
rect 43068 13338 43238 13353
rect 43068 13304 43069 13338
rect 43069 13304 43237 13338
rect 43237 13304 43238 13338
rect 43068 13289 43238 13304
rect 43440 13338 43610 13353
rect 43440 13304 43441 13338
rect 43441 13304 43609 13338
rect 43609 13304 43610 13338
rect 43440 13289 43610 13304
rect 45432 13071 45714 13343
rect 46176 13071 46458 13343
rect 46920 13071 47202 13343
rect 47664 13071 47946 13343
rect 48408 13071 48690 13343
rect 49152 13071 49434 13343
rect 49896 13071 50178 13343
rect 50640 13071 50922 13343
rect 39348 12750 39518 12763
rect 39348 12716 39349 12750
rect 39349 12716 39517 12750
rect 39517 12716 39518 12750
rect 39348 12703 39518 12716
rect 39720 12750 39890 12763
rect 39720 12716 39721 12750
rect 39721 12716 39889 12750
rect 39889 12716 39890 12750
rect 39720 12703 39890 12716
rect 40092 12750 40262 12763
rect 40092 12716 40093 12750
rect 40093 12716 40261 12750
rect 40261 12716 40262 12750
rect 40092 12703 40262 12716
rect 40464 12750 40634 12763
rect 40464 12716 40465 12750
rect 40465 12716 40633 12750
rect 40633 12716 40634 12750
rect 40464 12703 40634 12716
rect 40836 12750 41006 12763
rect 40836 12716 40837 12750
rect 40837 12716 41005 12750
rect 41005 12716 41006 12750
rect 40836 12703 41006 12716
rect 41208 12750 41378 12763
rect 41208 12716 41209 12750
rect 41209 12716 41377 12750
rect 41377 12716 41378 12750
rect 41208 12703 41378 12716
rect 41580 12750 41750 12763
rect 41580 12716 41581 12750
rect 41581 12716 41749 12750
rect 41749 12716 41750 12750
rect 41580 12703 41750 12716
rect 41952 12750 42122 12763
rect 41952 12716 41953 12750
rect 41953 12716 42121 12750
rect 42121 12716 42122 12750
rect 41952 12703 42122 12716
rect 42324 12750 42494 12763
rect 42324 12716 42325 12750
rect 42325 12716 42493 12750
rect 42493 12716 42494 12750
rect 42324 12703 42494 12716
rect 42696 12750 42866 12763
rect 42696 12716 42697 12750
rect 42697 12716 42865 12750
rect 42865 12716 42866 12750
rect 42696 12703 42866 12716
rect 43068 12750 43238 12763
rect 43068 12716 43069 12750
rect 43069 12716 43237 12750
rect 43237 12716 43238 12750
rect 43068 12703 43238 12716
rect 43440 12750 43610 12763
rect 43440 12716 43441 12750
rect 43441 12716 43609 12750
rect 43609 12716 43610 12750
rect 43440 12703 43610 12716
rect 43812 12750 43982 12763
rect 43812 12716 43813 12750
rect 43813 12716 43981 12750
rect 43981 12716 43982 12750
rect 43812 12703 43982 12716
rect 44184 12750 44354 12763
rect 44184 12716 44185 12750
rect 44185 12716 44353 12750
rect 44353 12716 44354 12750
rect 44184 12703 44354 12716
rect 44556 12750 44726 12763
rect 44556 12716 44557 12750
rect 44557 12716 44725 12750
rect 44725 12716 44726 12750
rect 44556 12703 44726 12716
rect 44928 12750 45098 12763
rect 44928 12716 44929 12750
rect 44929 12716 45097 12750
rect 45097 12716 45098 12750
rect 44928 12703 45098 12716
rect 45300 12750 45470 12763
rect 45300 12716 45301 12750
rect 45301 12716 45469 12750
rect 45469 12716 45470 12750
rect 45300 12703 45470 12716
rect 45672 12750 45842 12763
rect 45672 12716 45673 12750
rect 45673 12716 45841 12750
rect 45841 12716 45842 12750
rect 45672 12703 45842 12716
rect 46044 12750 46214 12763
rect 46044 12716 46045 12750
rect 46045 12716 46213 12750
rect 46213 12716 46214 12750
rect 46044 12703 46214 12716
rect 46416 12750 46586 12763
rect 46416 12716 46417 12750
rect 46417 12716 46585 12750
rect 46585 12716 46586 12750
rect 46416 12703 46586 12716
rect 46788 12750 46958 12763
rect 46788 12716 46789 12750
rect 46789 12716 46957 12750
rect 46957 12716 46958 12750
rect 46788 12703 46958 12716
rect 47160 12750 47330 12763
rect 47160 12716 47161 12750
rect 47161 12716 47329 12750
rect 47329 12716 47330 12750
rect 47160 12703 47330 12716
rect 47532 12750 47702 12763
rect 47532 12716 47533 12750
rect 47533 12716 47701 12750
rect 47701 12716 47702 12750
rect 47532 12703 47702 12716
rect 47904 12750 48074 12763
rect 47904 12716 47905 12750
rect 47905 12716 48073 12750
rect 48073 12716 48074 12750
rect 47904 12703 48074 12716
rect 48276 12750 48446 12763
rect 48276 12716 48277 12750
rect 48277 12716 48445 12750
rect 48445 12716 48446 12750
rect 48276 12703 48446 12716
rect 48648 12750 48818 12763
rect 48648 12716 48649 12750
rect 48649 12716 48817 12750
rect 48817 12716 48818 12750
rect 48648 12703 48818 12716
rect 49020 12750 49190 12763
rect 49020 12716 49021 12750
rect 49021 12716 49189 12750
rect 49189 12716 49190 12750
rect 49020 12703 49190 12716
rect 49392 12750 49562 12763
rect 49392 12716 49393 12750
rect 49393 12716 49561 12750
rect 49561 12716 49562 12750
rect 49392 12703 49562 12716
rect 49764 12750 49934 12763
rect 49764 12716 49765 12750
rect 49765 12716 49933 12750
rect 49933 12716 49934 12750
rect 49764 12703 49934 12716
rect 50136 12750 50306 12763
rect 50136 12716 50137 12750
rect 50137 12716 50305 12750
rect 50305 12716 50306 12750
rect 50136 12703 50306 12716
rect 50508 12750 50678 12763
rect 50508 12716 50509 12750
rect 50509 12716 50677 12750
rect 50677 12716 50678 12750
rect 50508 12703 50678 12716
rect 50880 12750 51050 12763
rect 50880 12716 50881 12750
rect 50881 12716 51049 12750
rect 51049 12716 51050 12750
rect 50880 12703 51050 12716
rect 39348 12222 39518 12223
rect 39348 12188 39349 12222
rect 39349 12188 39517 12222
rect 39517 12188 39518 12222
rect 39348 12114 39518 12188
rect 39348 12080 39349 12114
rect 39349 12080 39517 12114
rect 39517 12080 39518 12114
rect 39348 12079 39518 12080
rect 39720 12222 39890 12223
rect 39720 12188 39721 12222
rect 39721 12188 39889 12222
rect 39889 12188 39890 12222
rect 39720 12114 39890 12188
rect 39720 12080 39721 12114
rect 39721 12080 39889 12114
rect 39889 12080 39890 12114
rect 39720 12079 39890 12080
rect 40092 12222 40262 12223
rect 40092 12188 40093 12222
rect 40093 12188 40261 12222
rect 40261 12188 40262 12222
rect 40092 12114 40262 12188
rect 40092 12080 40093 12114
rect 40093 12080 40261 12114
rect 40261 12080 40262 12114
rect 40092 12079 40262 12080
rect 40464 12222 40634 12223
rect 40464 12188 40465 12222
rect 40465 12188 40633 12222
rect 40633 12188 40634 12222
rect 40464 12114 40634 12188
rect 40464 12080 40465 12114
rect 40465 12080 40633 12114
rect 40633 12080 40634 12114
rect 40464 12079 40634 12080
rect 40836 12222 41006 12223
rect 40836 12188 40837 12222
rect 40837 12188 41005 12222
rect 41005 12188 41006 12222
rect 40836 12114 41006 12188
rect 40836 12080 40837 12114
rect 40837 12080 41005 12114
rect 41005 12080 41006 12114
rect 40836 12079 41006 12080
rect 41208 12222 41378 12223
rect 41208 12188 41209 12222
rect 41209 12188 41377 12222
rect 41377 12188 41378 12222
rect 41208 12114 41378 12188
rect 41208 12080 41209 12114
rect 41209 12080 41377 12114
rect 41377 12080 41378 12114
rect 41208 12079 41378 12080
rect 41580 12222 41750 12223
rect 41580 12188 41581 12222
rect 41581 12188 41749 12222
rect 41749 12188 41750 12222
rect 41580 12114 41750 12188
rect 41580 12080 41581 12114
rect 41581 12080 41749 12114
rect 41749 12080 41750 12114
rect 41580 12079 41750 12080
rect 41952 12222 42122 12223
rect 41952 12188 41953 12222
rect 41953 12188 42121 12222
rect 42121 12188 42122 12222
rect 41952 12114 42122 12188
rect 41952 12080 41953 12114
rect 41953 12080 42121 12114
rect 42121 12080 42122 12114
rect 41952 12079 42122 12080
rect 42324 12222 42494 12223
rect 42324 12188 42325 12222
rect 42325 12188 42493 12222
rect 42493 12188 42494 12222
rect 42324 12114 42494 12188
rect 42324 12080 42325 12114
rect 42325 12080 42493 12114
rect 42493 12080 42494 12114
rect 42324 12079 42494 12080
rect 42696 12222 42866 12223
rect 42696 12188 42697 12222
rect 42697 12188 42865 12222
rect 42865 12188 42866 12222
rect 42696 12114 42866 12188
rect 42696 12080 42697 12114
rect 42697 12080 42865 12114
rect 42865 12080 42866 12114
rect 42696 12079 42866 12080
rect 43068 12222 43238 12223
rect 43068 12188 43069 12222
rect 43069 12188 43237 12222
rect 43237 12188 43238 12222
rect 43068 12114 43238 12188
rect 43068 12080 43069 12114
rect 43069 12080 43237 12114
rect 43237 12080 43238 12114
rect 43068 12079 43238 12080
rect 43440 12222 43610 12223
rect 43440 12188 43441 12222
rect 43441 12188 43609 12222
rect 43609 12188 43610 12222
rect 43440 12114 43610 12188
rect 43440 12080 43441 12114
rect 43441 12080 43609 12114
rect 43609 12080 43610 12114
rect 43440 12079 43610 12080
rect 43812 12222 43982 12223
rect 43812 12188 43813 12222
rect 43813 12188 43981 12222
rect 43981 12188 43982 12222
rect 43812 12114 43982 12188
rect 43812 12080 43813 12114
rect 43813 12080 43981 12114
rect 43981 12080 43982 12114
rect 43812 12079 43982 12080
rect 44184 12222 44354 12223
rect 44184 12188 44185 12222
rect 44185 12188 44353 12222
rect 44353 12188 44354 12222
rect 44184 12114 44354 12188
rect 44184 12080 44185 12114
rect 44185 12080 44353 12114
rect 44353 12080 44354 12114
rect 44184 12079 44354 12080
rect 44556 12222 44726 12223
rect 44556 12188 44557 12222
rect 44557 12188 44725 12222
rect 44725 12188 44726 12222
rect 44556 12114 44726 12188
rect 44556 12080 44557 12114
rect 44557 12080 44725 12114
rect 44725 12080 44726 12114
rect 44556 12079 44726 12080
rect 44928 12222 45098 12223
rect 44928 12188 44929 12222
rect 44929 12188 45097 12222
rect 45097 12188 45098 12222
rect 44928 12114 45098 12188
rect 44928 12080 44929 12114
rect 44929 12080 45097 12114
rect 45097 12080 45098 12114
rect 44928 12079 45098 12080
rect 39348 11586 39518 11587
rect 39348 11552 39349 11586
rect 39349 11552 39517 11586
rect 39517 11552 39518 11586
rect 39348 11478 39518 11552
rect 39348 11444 39349 11478
rect 39349 11444 39517 11478
rect 39517 11444 39518 11478
rect 39348 11443 39518 11444
rect 39720 11586 39890 11587
rect 39720 11552 39721 11586
rect 39721 11552 39889 11586
rect 39889 11552 39890 11586
rect 39720 11478 39890 11552
rect 39720 11444 39721 11478
rect 39721 11444 39889 11478
rect 39889 11444 39890 11478
rect 39720 11443 39890 11444
rect 40092 11586 40262 11587
rect 40092 11552 40093 11586
rect 40093 11552 40261 11586
rect 40261 11552 40262 11586
rect 40092 11478 40262 11552
rect 40092 11444 40093 11478
rect 40093 11444 40261 11478
rect 40261 11444 40262 11478
rect 40092 11443 40262 11444
rect 40464 11586 40634 11587
rect 40464 11552 40465 11586
rect 40465 11552 40633 11586
rect 40633 11552 40634 11586
rect 40464 11478 40634 11552
rect 40464 11444 40465 11478
rect 40465 11444 40633 11478
rect 40633 11444 40634 11478
rect 40464 11443 40634 11444
rect 40836 11586 41006 11587
rect 40836 11552 40837 11586
rect 40837 11552 41005 11586
rect 41005 11552 41006 11586
rect 40836 11478 41006 11552
rect 40836 11444 40837 11478
rect 40837 11444 41005 11478
rect 41005 11444 41006 11478
rect 40836 11443 41006 11444
rect 41208 11586 41378 11587
rect 41208 11552 41209 11586
rect 41209 11552 41377 11586
rect 41377 11552 41378 11586
rect 41208 11478 41378 11552
rect 41208 11444 41209 11478
rect 41209 11444 41377 11478
rect 41377 11444 41378 11478
rect 41208 11443 41378 11444
rect 41580 11586 41750 11587
rect 41580 11552 41581 11586
rect 41581 11552 41749 11586
rect 41749 11552 41750 11586
rect 41580 11478 41750 11552
rect 41580 11444 41581 11478
rect 41581 11444 41749 11478
rect 41749 11444 41750 11478
rect 41580 11443 41750 11444
rect 41952 11586 42122 11587
rect 41952 11552 41953 11586
rect 41953 11552 42121 11586
rect 42121 11552 42122 11586
rect 41952 11478 42122 11552
rect 41952 11444 41953 11478
rect 41953 11444 42121 11478
rect 42121 11444 42122 11478
rect 41952 11443 42122 11444
rect 42324 11586 42494 11587
rect 42324 11552 42325 11586
rect 42325 11552 42493 11586
rect 42493 11552 42494 11586
rect 42324 11478 42494 11552
rect 42324 11444 42325 11478
rect 42325 11444 42493 11478
rect 42493 11444 42494 11478
rect 42324 11443 42494 11444
rect 42696 11586 42866 11587
rect 42696 11552 42697 11586
rect 42697 11552 42865 11586
rect 42865 11552 42866 11586
rect 42696 11478 42866 11552
rect 42696 11444 42697 11478
rect 42697 11444 42865 11478
rect 42865 11444 42866 11478
rect 42696 11443 42866 11444
rect 43068 11586 43238 11587
rect 43068 11552 43069 11586
rect 43069 11552 43237 11586
rect 43237 11552 43238 11586
rect 43068 11478 43238 11552
rect 43068 11444 43069 11478
rect 43069 11444 43237 11478
rect 43237 11444 43238 11478
rect 43068 11443 43238 11444
rect 43440 11586 43610 11587
rect 43440 11552 43441 11586
rect 43441 11552 43609 11586
rect 43609 11552 43610 11586
rect 43440 11478 43610 11552
rect 43440 11444 43441 11478
rect 43441 11444 43609 11478
rect 43609 11444 43610 11478
rect 43440 11443 43610 11444
rect 43812 11586 43982 11587
rect 43812 11552 43813 11586
rect 43813 11552 43981 11586
rect 43981 11552 43982 11586
rect 43812 11478 43982 11552
rect 43812 11444 43813 11478
rect 43813 11444 43981 11478
rect 43981 11444 43982 11478
rect 43812 11443 43982 11444
rect 44184 11586 44354 11587
rect 44184 11552 44185 11586
rect 44185 11552 44353 11586
rect 44353 11552 44354 11586
rect 44184 11478 44354 11552
rect 44184 11444 44185 11478
rect 44185 11444 44353 11478
rect 44353 11444 44354 11478
rect 44184 11443 44354 11444
rect 44556 11586 44726 11587
rect 44556 11552 44557 11586
rect 44557 11552 44725 11586
rect 44725 11552 44726 11586
rect 44556 11478 44726 11552
rect 44556 11444 44557 11478
rect 44557 11444 44725 11478
rect 44725 11444 44726 11478
rect 44556 11443 44726 11444
rect 44928 11586 45098 11587
rect 44928 11552 44929 11586
rect 44929 11552 45097 11586
rect 45097 11552 45098 11586
rect 44928 11478 45098 11552
rect 44928 11444 44929 11478
rect 44929 11444 45097 11478
rect 45097 11444 45098 11478
rect 44928 11443 45098 11444
rect 39348 10950 39518 10963
rect 39348 10916 39349 10950
rect 39349 10916 39517 10950
rect 39517 10916 39518 10950
rect 39348 10903 39518 10916
rect 39720 10950 39890 10963
rect 39720 10916 39721 10950
rect 39721 10916 39889 10950
rect 39889 10916 39890 10950
rect 39720 10903 39890 10916
rect 40092 10950 40262 10963
rect 40092 10916 40093 10950
rect 40093 10916 40261 10950
rect 40261 10916 40262 10950
rect 40092 10903 40262 10916
rect 40464 10950 40634 10963
rect 40464 10916 40465 10950
rect 40465 10916 40633 10950
rect 40633 10916 40634 10950
rect 40464 10903 40634 10916
rect 40836 10950 41006 10963
rect 40836 10916 40837 10950
rect 40837 10916 41005 10950
rect 41005 10916 41006 10950
rect 40836 10903 41006 10916
rect 41208 10950 41378 10963
rect 41208 10916 41209 10950
rect 41209 10916 41377 10950
rect 41377 10916 41378 10950
rect 41208 10903 41378 10916
rect 41580 10950 41750 10963
rect 41580 10916 41581 10950
rect 41581 10916 41749 10950
rect 41749 10916 41750 10950
rect 41580 10903 41750 10916
rect 41952 10950 42122 10963
rect 41952 10916 41953 10950
rect 41953 10916 42121 10950
rect 42121 10916 42122 10950
rect 41952 10903 42122 10916
rect 42324 10950 42494 10963
rect 42324 10916 42325 10950
rect 42325 10916 42493 10950
rect 42493 10916 42494 10950
rect 42324 10903 42494 10916
rect 42696 10950 42866 10963
rect 42696 10916 42697 10950
rect 42697 10916 42865 10950
rect 42865 10916 42866 10950
rect 42696 10903 42866 10916
rect 43068 10950 43238 10963
rect 43068 10916 43069 10950
rect 43069 10916 43237 10950
rect 43237 10916 43238 10950
rect 43068 10903 43238 10916
rect 43440 10950 43610 10963
rect 43440 10916 43441 10950
rect 43441 10916 43609 10950
rect 43609 10916 43610 10950
rect 43440 10903 43610 10916
rect 43812 10950 43982 10963
rect 43812 10916 43813 10950
rect 43813 10916 43981 10950
rect 43981 10916 43982 10950
rect 43812 10903 43982 10916
rect 44184 10950 44354 10963
rect 44184 10916 44185 10950
rect 44185 10916 44353 10950
rect 44353 10916 44354 10950
rect 44184 10903 44354 10916
rect 44556 10950 44726 10963
rect 44556 10916 44557 10950
rect 44557 10916 44725 10950
rect 44725 10916 44726 10950
rect 44556 10903 44726 10916
rect 44928 10950 45098 10963
rect 44928 10916 44929 10950
rect 44929 10916 45097 10950
rect 45097 10916 45098 10950
rect 44928 10903 45098 10916
rect 45300 12222 45470 12223
rect 45300 12188 45301 12222
rect 45301 12188 45469 12222
rect 45469 12188 45470 12222
rect 45300 12114 45470 12188
rect 45300 12080 45301 12114
rect 45301 12080 45469 12114
rect 45469 12080 45470 12114
rect 45300 12079 45470 12080
rect 45672 12222 45842 12223
rect 45672 12188 45673 12222
rect 45673 12188 45841 12222
rect 45841 12188 45842 12222
rect 45672 12114 45842 12188
rect 45672 12080 45673 12114
rect 45673 12080 45841 12114
rect 45841 12080 45842 12114
rect 45672 12079 45842 12080
rect 46044 12222 46214 12223
rect 46044 12188 46045 12222
rect 46045 12188 46213 12222
rect 46213 12188 46214 12222
rect 46044 12114 46214 12188
rect 46044 12080 46045 12114
rect 46045 12080 46213 12114
rect 46213 12080 46214 12114
rect 46044 12079 46214 12080
rect 46416 12222 46586 12223
rect 46416 12188 46417 12222
rect 46417 12188 46585 12222
rect 46585 12188 46586 12222
rect 46416 12114 46586 12188
rect 46416 12080 46417 12114
rect 46417 12080 46585 12114
rect 46585 12080 46586 12114
rect 46416 12079 46586 12080
rect 46788 12222 46958 12223
rect 46788 12188 46789 12222
rect 46789 12188 46957 12222
rect 46957 12188 46958 12222
rect 46788 12114 46958 12188
rect 46788 12080 46789 12114
rect 46789 12080 46957 12114
rect 46957 12080 46958 12114
rect 46788 12079 46958 12080
rect 47160 12222 47330 12223
rect 47160 12188 47161 12222
rect 47161 12188 47329 12222
rect 47329 12188 47330 12222
rect 47160 12114 47330 12188
rect 47160 12080 47161 12114
rect 47161 12080 47329 12114
rect 47329 12080 47330 12114
rect 47160 12079 47330 12080
rect 47532 12222 47702 12223
rect 47532 12188 47533 12222
rect 47533 12188 47701 12222
rect 47701 12188 47702 12222
rect 47532 12114 47702 12188
rect 47532 12080 47533 12114
rect 47533 12080 47701 12114
rect 47701 12080 47702 12114
rect 47532 12079 47702 12080
rect 47904 12222 48074 12223
rect 47904 12188 47905 12222
rect 47905 12188 48073 12222
rect 48073 12188 48074 12222
rect 47904 12114 48074 12188
rect 47904 12080 47905 12114
rect 47905 12080 48073 12114
rect 48073 12080 48074 12114
rect 47904 12079 48074 12080
rect 48276 12222 48446 12223
rect 48276 12188 48277 12222
rect 48277 12188 48445 12222
rect 48445 12188 48446 12222
rect 48276 12114 48446 12188
rect 48276 12080 48277 12114
rect 48277 12080 48445 12114
rect 48445 12080 48446 12114
rect 48276 12079 48446 12080
rect 48648 12222 48818 12223
rect 48648 12188 48649 12222
rect 48649 12188 48817 12222
rect 48817 12188 48818 12222
rect 48648 12114 48818 12188
rect 48648 12080 48649 12114
rect 48649 12080 48817 12114
rect 48817 12080 48818 12114
rect 48648 12079 48818 12080
rect 49020 12222 49190 12223
rect 49020 12188 49021 12222
rect 49021 12188 49189 12222
rect 49189 12188 49190 12222
rect 49020 12114 49190 12188
rect 49020 12080 49021 12114
rect 49021 12080 49189 12114
rect 49189 12080 49190 12114
rect 49020 12079 49190 12080
rect 49392 12222 49562 12223
rect 49392 12188 49393 12222
rect 49393 12188 49561 12222
rect 49561 12188 49562 12222
rect 49392 12114 49562 12188
rect 49392 12080 49393 12114
rect 49393 12080 49561 12114
rect 49561 12080 49562 12114
rect 49392 12079 49562 12080
rect 49764 12222 49934 12223
rect 49764 12188 49765 12222
rect 49765 12188 49933 12222
rect 49933 12188 49934 12222
rect 49764 12114 49934 12188
rect 49764 12080 49765 12114
rect 49765 12080 49933 12114
rect 49933 12080 49934 12114
rect 49764 12079 49934 12080
rect 50136 12222 50306 12223
rect 50136 12188 50137 12222
rect 50137 12188 50305 12222
rect 50305 12188 50306 12222
rect 50136 12114 50306 12188
rect 50136 12080 50137 12114
rect 50137 12080 50305 12114
rect 50305 12080 50306 12114
rect 50136 12079 50306 12080
rect 50508 12222 50678 12223
rect 50508 12188 50509 12222
rect 50509 12188 50677 12222
rect 50677 12188 50678 12222
rect 50508 12114 50678 12188
rect 50508 12080 50509 12114
rect 50509 12080 50677 12114
rect 50677 12080 50678 12114
rect 50508 12079 50678 12080
rect 50880 12222 51050 12223
rect 50880 12188 50881 12222
rect 50881 12188 51049 12222
rect 51049 12188 51050 12222
rect 50880 12114 51050 12188
rect 50880 12080 50881 12114
rect 50881 12080 51049 12114
rect 51049 12080 51050 12114
rect 50880 12079 51050 12080
rect 45300 11586 45470 11587
rect 45300 11552 45301 11586
rect 45301 11552 45469 11586
rect 45469 11552 45470 11586
rect 45300 11478 45470 11552
rect 45300 11444 45301 11478
rect 45301 11444 45469 11478
rect 45469 11444 45470 11478
rect 45300 11443 45470 11444
rect 45672 11586 45842 11587
rect 45672 11552 45673 11586
rect 45673 11552 45841 11586
rect 45841 11552 45842 11586
rect 45672 11478 45842 11552
rect 45672 11444 45673 11478
rect 45673 11444 45841 11478
rect 45841 11444 45842 11478
rect 45672 11443 45842 11444
rect 46044 11586 46214 11587
rect 46044 11552 46045 11586
rect 46045 11552 46213 11586
rect 46213 11552 46214 11586
rect 46044 11478 46214 11552
rect 46044 11444 46045 11478
rect 46045 11444 46213 11478
rect 46213 11444 46214 11478
rect 46044 11443 46214 11444
rect 46416 11586 46586 11587
rect 46416 11552 46417 11586
rect 46417 11552 46585 11586
rect 46585 11552 46586 11586
rect 46416 11478 46586 11552
rect 46416 11444 46417 11478
rect 46417 11444 46585 11478
rect 46585 11444 46586 11478
rect 46416 11443 46586 11444
rect 46788 11586 46958 11587
rect 46788 11552 46789 11586
rect 46789 11552 46957 11586
rect 46957 11552 46958 11586
rect 46788 11478 46958 11552
rect 46788 11444 46789 11478
rect 46789 11444 46957 11478
rect 46957 11444 46958 11478
rect 46788 11443 46958 11444
rect 47160 11586 47330 11587
rect 47160 11552 47161 11586
rect 47161 11552 47329 11586
rect 47329 11552 47330 11586
rect 47160 11478 47330 11552
rect 47160 11444 47161 11478
rect 47161 11444 47329 11478
rect 47329 11444 47330 11478
rect 47160 11443 47330 11444
rect 47532 11586 47702 11587
rect 47532 11552 47533 11586
rect 47533 11552 47701 11586
rect 47701 11552 47702 11586
rect 47532 11478 47702 11552
rect 47532 11444 47533 11478
rect 47533 11444 47701 11478
rect 47701 11444 47702 11478
rect 47532 11443 47702 11444
rect 47904 11586 48074 11587
rect 47904 11552 47905 11586
rect 47905 11552 48073 11586
rect 48073 11552 48074 11586
rect 47904 11478 48074 11552
rect 47904 11444 47905 11478
rect 47905 11444 48073 11478
rect 48073 11444 48074 11478
rect 47904 11443 48074 11444
rect 48276 11586 48446 11587
rect 48276 11552 48277 11586
rect 48277 11552 48445 11586
rect 48445 11552 48446 11586
rect 48276 11478 48446 11552
rect 48276 11444 48277 11478
rect 48277 11444 48445 11478
rect 48445 11444 48446 11478
rect 48276 11443 48446 11444
rect 48648 11586 48818 11587
rect 48648 11552 48649 11586
rect 48649 11552 48817 11586
rect 48817 11552 48818 11586
rect 48648 11478 48818 11552
rect 48648 11444 48649 11478
rect 48649 11444 48817 11478
rect 48817 11444 48818 11478
rect 48648 11443 48818 11444
rect 49020 11586 49190 11587
rect 49020 11552 49021 11586
rect 49021 11552 49189 11586
rect 49189 11552 49190 11586
rect 49020 11478 49190 11552
rect 49020 11444 49021 11478
rect 49021 11444 49189 11478
rect 49189 11444 49190 11478
rect 49020 11443 49190 11444
rect 49392 11586 49562 11587
rect 49392 11552 49393 11586
rect 49393 11552 49561 11586
rect 49561 11552 49562 11586
rect 49392 11478 49562 11552
rect 49392 11444 49393 11478
rect 49393 11444 49561 11478
rect 49561 11444 49562 11478
rect 49392 11443 49562 11444
rect 49764 11586 49934 11587
rect 49764 11552 49765 11586
rect 49765 11552 49933 11586
rect 49933 11552 49934 11586
rect 49764 11478 49934 11552
rect 49764 11444 49765 11478
rect 49765 11444 49933 11478
rect 49933 11444 49934 11478
rect 49764 11443 49934 11444
rect 50136 11586 50306 11587
rect 50136 11552 50137 11586
rect 50137 11552 50305 11586
rect 50305 11552 50306 11586
rect 50136 11478 50306 11552
rect 50136 11444 50137 11478
rect 50137 11444 50305 11478
rect 50305 11444 50306 11478
rect 50136 11443 50306 11444
rect 50508 11586 50678 11587
rect 50508 11552 50509 11586
rect 50509 11552 50677 11586
rect 50677 11552 50678 11586
rect 50508 11478 50678 11552
rect 50508 11444 50509 11478
rect 50509 11444 50677 11478
rect 50677 11444 50678 11478
rect 50508 11443 50678 11444
rect 50880 11586 51050 11587
rect 50880 11552 50881 11586
rect 50881 11552 51049 11586
rect 51049 11552 51050 11586
rect 50880 11478 51050 11552
rect 50880 11444 50881 11478
rect 50881 11444 51049 11478
rect 51049 11444 51050 11478
rect 50880 11443 51050 11444
rect 45300 10950 45470 10963
rect 45300 10916 45301 10950
rect 45301 10916 45469 10950
rect 45469 10916 45470 10950
rect 45300 10903 45470 10916
rect 45672 10950 45842 10963
rect 45672 10916 45673 10950
rect 45673 10916 45841 10950
rect 45841 10916 45842 10950
rect 45672 10903 45842 10916
rect 46044 10950 46214 10963
rect 46044 10916 46045 10950
rect 46045 10916 46213 10950
rect 46213 10916 46214 10950
rect 46044 10903 46214 10916
rect 46416 10950 46586 10963
rect 46416 10916 46417 10950
rect 46417 10916 46585 10950
rect 46585 10916 46586 10950
rect 46416 10903 46586 10916
rect 46788 10950 46958 10963
rect 46788 10916 46789 10950
rect 46789 10916 46957 10950
rect 46957 10916 46958 10950
rect 46788 10903 46958 10916
rect 47160 10950 47330 10963
rect 47160 10916 47161 10950
rect 47161 10916 47329 10950
rect 47329 10916 47330 10950
rect 47160 10903 47330 10916
rect 47532 10950 47702 10963
rect 47532 10916 47533 10950
rect 47533 10916 47701 10950
rect 47701 10916 47702 10950
rect 47532 10903 47702 10916
rect 47904 10950 48074 10963
rect 47904 10916 47905 10950
rect 47905 10916 48073 10950
rect 48073 10916 48074 10950
rect 47904 10903 48074 10916
rect 48276 10950 48446 10963
rect 48276 10916 48277 10950
rect 48277 10916 48445 10950
rect 48445 10916 48446 10950
rect 48276 10903 48446 10916
rect 48648 10950 48818 10963
rect 48648 10916 48649 10950
rect 48649 10916 48817 10950
rect 48817 10916 48818 10950
rect 48648 10903 48818 10916
rect 49020 10950 49190 10963
rect 49020 10916 49021 10950
rect 49021 10916 49189 10950
rect 49189 10916 49190 10950
rect 49020 10903 49190 10916
rect 49392 10950 49562 10963
rect 49392 10916 49393 10950
rect 49393 10916 49561 10950
rect 49561 10916 49562 10950
rect 49392 10903 49562 10916
rect 49764 10950 49934 10963
rect 49764 10916 49765 10950
rect 49765 10916 49933 10950
rect 49933 10916 49934 10950
rect 49764 10903 49934 10916
rect 50136 10950 50306 10963
rect 50136 10916 50137 10950
rect 50137 10916 50305 10950
rect 50305 10916 50306 10950
rect 50136 10903 50306 10916
rect 50508 10950 50678 10963
rect 50508 10916 50509 10950
rect 50509 10916 50677 10950
rect 50677 10916 50678 10950
rect 50508 10903 50678 10916
rect 50880 10950 51050 10963
rect 50880 10916 50881 10950
rect 50881 10916 51049 10950
rect 51049 10916 51050 10950
rect 50880 10903 51050 10916
rect 39518 10515 39718 10715
rect 40262 10515 40462 10715
rect 41006 10515 41206 10715
rect 41750 10515 41950 10715
rect 42494 10515 42694 10715
rect 43238 10515 43438 10715
rect 43982 10515 44182 10715
rect 44726 10515 44926 10715
rect 45098 10515 45298 10715
rect 45842 10515 46042 10715
rect 46586 10515 46786 10715
rect 47330 10515 47530 10715
rect 48074 10515 48274 10715
rect 48818 10515 49018 10715
rect 49562 10515 49762 10715
rect 50306 10515 50506 10715
rect 51050 10515 51250 10715
rect 39518 9150 39718 9350
rect 40262 9150 40462 9350
rect 41006 9150 41206 9350
rect 41750 9150 41950 9350
rect 42494 9150 42694 9350
rect 43238 9150 43438 9350
rect 43982 9150 44182 9350
rect 44726 9150 44926 9350
rect 45098 9150 45298 9350
rect 45842 9150 46042 9350
rect 46586 9150 46786 9350
rect 47330 9150 47530 9350
rect 48074 9150 48274 9350
rect 48818 9150 49018 9350
rect 49562 9150 49762 9350
rect 50306 9150 50506 9350
rect 51050 9150 51250 9350
rect 39348 8949 39518 8962
rect 39348 8915 39349 8949
rect 39349 8915 39517 8949
rect 39517 8915 39518 8949
rect 39348 8902 39518 8915
rect 39720 8949 39890 8962
rect 39720 8915 39721 8949
rect 39721 8915 39889 8949
rect 39889 8915 39890 8949
rect 39720 8902 39890 8915
rect 40092 8949 40262 8962
rect 40092 8915 40093 8949
rect 40093 8915 40261 8949
rect 40261 8915 40262 8949
rect 40092 8902 40262 8915
rect 40464 8949 40634 8962
rect 40464 8915 40465 8949
rect 40465 8915 40633 8949
rect 40633 8915 40634 8949
rect 40464 8902 40634 8915
rect 40836 8949 41006 8962
rect 40836 8915 40837 8949
rect 40837 8915 41005 8949
rect 41005 8915 41006 8949
rect 40836 8902 41006 8915
rect 41208 8949 41378 8962
rect 41208 8915 41209 8949
rect 41209 8915 41377 8949
rect 41377 8915 41378 8949
rect 41208 8902 41378 8915
rect 41580 8949 41750 8962
rect 41580 8915 41581 8949
rect 41581 8915 41749 8949
rect 41749 8915 41750 8949
rect 41580 8902 41750 8915
rect 41952 8949 42122 8962
rect 41952 8915 41953 8949
rect 41953 8915 42121 8949
rect 42121 8915 42122 8949
rect 41952 8902 42122 8915
rect 42324 8949 42494 8962
rect 42324 8915 42325 8949
rect 42325 8915 42493 8949
rect 42493 8915 42494 8949
rect 42324 8902 42494 8915
rect 42696 8949 42866 8962
rect 42696 8915 42697 8949
rect 42697 8915 42865 8949
rect 42865 8915 42866 8949
rect 42696 8902 42866 8915
rect 43068 8949 43238 8962
rect 43068 8915 43069 8949
rect 43069 8915 43237 8949
rect 43237 8915 43238 8949
rect 43068 8902 43238 8915
rect 43440 8949 43610 8962
rect 43440 8915 43441 8949
rect 43441 8915 43609 8949
rect 43609 8915 43610 8949
rect 43440 8902 43610 8915
rect 43812 8949 43982 8962
rect 43812 8915 43813 8949
rect 43813 8915 43981 8949
rect 43981 8915 43982 8949
rect 43812 8902 43982 8915
rect 44184 8949 44354 8962
rect 44184 8915 44185 8949
rect 44185 8915 44353 8949
rect 44353 8915 44354 8949
rect 44184 8902 44354 8915
rect 44556 8949 44726 8962
rect 44556 8915 44557 8949
rect 44557 8915 44725 8949
rect 44725 8915 44726 8949
rect 44556 8902 44726 8915
rect 44928 8949 45098 8962
rect 44928 8915 44929 8949
rect 44929 8915 45097 8949
rect 45097 8915 45098 8949
rect 44928 8902 45098 8915
rect 39348 8421 39518 8422
rect 39348 8387 39349 8421
rect 39349 8387 39517 8421
rect 39517 8387 39518 8421
rect 39348 8313 39518 8387
rect 39348 8279 39349 8313
rect 39349 8279 39517 8313
rect 39517 8279 39518 8313
rect 39348 8278 39518 8279
rect 39720 8421 39890 8422
rect 39720 8387 39721 8421
rect 39721 8387 39889 8421
rect 39889 8387 39890 8421
rect 39720 8313 39890 8387
rect 39720 8279 39721 8313
rect 39721 8279 39889 8313
rect 39889 8279 39890 8313
rect 39720 8278 39890 8279
rect 40092 8421 40262 8422
rect 40092 8387 40093 8421
rect 40093 8387 40261 8421
rect 40261 8387 40262 8421
rect 40092 8313 40262 8387
rect 40092 8279 40093 8313
rect 40093 8279 40261 8313
rect 40261 8279 40262 8313
rect 40092 8278 40262 8279
rect 40464 8421 40634 8422
rect 40464 8387 40465 8421
rect 40465 8387 40633 8421
rect 40633 8387 40634 8421
rect 40464 8313 40634 8387
rect 40464 8279 40465 8313
rect 40465 8279 40633 8313
rect 40633 8279 40634 8313
rect 40464 8278 40634 8279
rect 40836 8421 41006 8422
rect 40836 8387 40837 8421
rect 40837 8387 41005 8421
rect 41005 8387 41006 8421
rect 40836 8313 41006 8387
rect 40836 8279 40837 8313
rect 40837 8279 41005 8313
rect 41005 8279 41006 8313
rect 40836 8278 41006 8279
rect 41208 8421 41378 8422
rect 41208 8387 41209 8421
rect 41209 8387 41377 8421
rect 41377 8387 41378 8421
rect 41208 8313 41378 8387
rect 41208 8279 41209 8313
rect 41209 8279 41377 8313
rect 41377 8279 41378 8313
rect 41208 8278 41378 8279
rect 41580 8421 41750 8422
rect 41580 8387 41581 8421
rect 41581 8387 41749 8421
rect 41749 8387 41750 8421
rect 41580 8313 41750 8387
rect 41580 8279 41581 8313
rect 41581 8279 41749 8313
rect 41749 8279 41750 8313
rect 41580 8278 41750 8279
rect 41952 8421 42122 8422
rect 41952 8387 41953 8421
rect 41953 8387 42121 8421
rect 42121 8387 42122 8421
rect 41952 8313 42122 8387
rect 41952 8279 41953 8313
rect 41953 8279 42121 8313
rect 42121 8279 42122 8313
rect 41952 8278 42122 8279
rect 42324 8421 42494 8422
rect 42324 8387 42325 8421
rect 42325 8387 42493 8421
rect 42493 8387 42494 8421
rect 42324 8313 42494 8387
rect 42324 8279 42325 8313
rect 42325 8279 42493 8313
rect 42493 8279 42494 8313
rect 42324 8278 42494 8279
rect 42696 8421 42866 8422
rect 42696 8387 42697 8421
rect 42697 8387 42865 8421
rect 42865 8387 42866 8421
rect 42696 8313 42866 8387
rect 42696 8279 42697 8313
rect 42697 8279 42865 8313
rect 42865 8279 42866 8313
rect 42696 8278 42866 8279
rect 43068 8421 43238 8422
rect 43068 8387 43069 8421
rect 43069 8387 43237 8421
rect 43237 8387 43238 8421
rect 43068 8313 43238 8387
rect 43068 8279 43069 8313
rect 43069 8279 43237 8313
rect 43237 8279 43238 8313
rect 43068 8278 43238 8279
rect 43440 8421 43610 8422
rect 43440 8387 43441 8421
rect 43441 8387 43609 8421
rect 43609 8387 43610 8421
rect 43440 8313 43610 8387
rect 43440 8279 43441 8313
rect 43441 8279 43609 8313
rect 43609 8279 43610 8313
rect 43440 8278 43610 8279
rect 43812 8421 43982 8422
rect 43812 8387 43813 8421
rect 43813 8387 43981 8421
rect 43981 8387 43982 8421
rect 43812 8313 43982 8387
rect 43812 8279 43813 8313
rect 43813 8279 43981 8313
rect 43981 8279 43982 8313
rect 43812 8278 43982 8279
rect 44184 8421 44354 8422
rect 44184 8387 44185 8421
rect 44185 8387 44353 8421
rect 44353 8387 44354 8421
rect 44184 8313 44354 8387
rect 44184 8279 44185 8313
rect 44185 8279 44353 8313
rect 44353 8279 44354 8313
rect 44184 8278 44354 8279
rect 44556 8421 44726 8422
rect 44556 8387 44557 8421
rect 44557 8387 44725 8421
rect 44725 8387 44726 8421
rect 44556 8313 44726 8387
rect 44556 8279 44557 8313
rect 44557 8279 44725 8313
rect 44725 8279 44726 8313
rect 44556 8278 44726 8279
rect 44928 8421 45098 8422
rect 44928 8387 44929 8421
rect 44929 8387 45097 8421
rect 45097 8387 45098 8421
rect 44928 8313 45098 8387
rect 44928 8279 44929 8313
rect 44929 8279 45097 8313
rect 45097 8279 45098 8313
rect 44928 8278 45098 8279
rect 39348 7785 39518 7786
rect 39348 7751 39349 7785
rect 39349 7751 39517 7785
rect 39517 7751 39518 7785
rect 39348 7677 39518 7751
rect 39348 7643 39349 7677
rect 39349 7643 39517 7677
rect 39517 7643 39518 7677
rect 39348 7642 39518 7643
rect 39720 7785 39890 7786
rect 39720 7751 39721 7785
rect 39721 7751 39889 7785
rect 39889 7751 39890 7785
rect 39720 7677 39890 7751
rect 39720 7643 39721 7677
rect 39721 7643 39889 7677
rect 39889 7643 39890 7677
rect 39720 7642 39890 7643
rect 40092 7785 40262 7786
rect 40092 7751 40093 7785
rect 40093 7751 40261 7785
rect 40261 7751 40262 7785
rect 40092 7677 40262 7751
rect 40092 7643 40093 7677
rect 40093 7643 40261 7677
rect 40261 7643 40262 7677
rect 40092 7642 40262 7643
rect 40464 7785 40634 7786
rect 40464 7751 40465 7785
rect 40465 7751 40633 7785
rect 40633 7751 40634 7785
rect 40464 7677 40634 7751
rect 40464 7643 40465 7677
rect 40465 7643 40633 7677
rect 40633 7643 40634 7677
rect 40464 7642 40634 7643
rect 40836 7785 41006 7786
rect 40836 7751 40837 7785
rect 40837 7751 41005 7785
rect 41005 7751 41006 7785
rect 40836 7677 41006 7751
rect 40836 7643 40837 7677
rect 40837 7643 41005 7677
rect 41005 7643 41006 7677
rect 40836 7642 41006 7643
rect 41208 7785 41378 7786
rect 41208 7751 41209 7785
rect 41209 7751 41377 7785
rect 41377 7751 41378 7785
rect 41208 7677 41378 7751
rect 41208 7643 41209 7677
rect 41209 7643 41377 7677
rect 41377 7643 41378 7677
rect 41208 7642 41378 7643
rect 41580 7785 41750 7786
rect 41580 7751 41581 7785
rect 41581 7751 41749 7785
rect 41749 7751 41750 7785
rect 41580 7677 41750 7751
rect 41580 7643 41581 7677
rect 41581 7643 41749 7677
rect 41749 7643 41750 7677
rect 41580 7642 41750 7643
rect 41952 7785 42122 7786
rect 41952 7751 41953 7785
rect 41953 7751 42121 7785
rect 42121 7751 42122 7785
rect 41952 7677 42122 7751
rect 41952 7643 41953 7677
rect 41953 7643 42121 7677
rect 42121 7643 42122 7677
rect 41952 7642 42122 7643
rect 42324 7785 42494 7786
rect 42324 7751 42325 7785
rect 42325 7751 42493 7785
rect 42493 7751 42494 7785
rect 42324 7677 42494 7751
rect 42324 7643 42325 7677
rect 42325 7643 42493 7677
rect 42493 7643 42494 7677
rect 42324 7642 42494 7643
rect 42696 7785 42866 7786
rect 42696 7751 42697 7785
rect 42697 7751 42865 7785
rect 42865 7751 42866 7785
rect 42696 7677 42866 7751
rect 42696 7643 42697 7677
rect 42697 7643 42865 7677
rect 42865 7643 42866 7677
rect 42696 7642 42866 7643
rect 43068 7785 43238 7786
rect 43068 7751 43069 7785
rect 43069 7751 43237 7785
rect 43237 7751 43238 7785
rect 43068 7677 43238 7751
rect 43068 7643 43069 7677
rect 43069 7643 43237 7677
rect 43237 7643 43238 7677
rect 43068 7642 43238 7643
rect 43440 7785 43610 7786
rect 43440 7751 43441 7785
rect 43441 7751 43609 7785
rect 43609 7751 43610 7785
rect 43440 7677 43610 7751
rect 43440 7643 43441 7677
rect 43441 7643 43609 7677
rect 43609 7643 43610 7677
rect 43440 7642 43610 7643
rect 43812 7785 43982 7786
rect 43812 7751 43813 7785
rect 43813 7751 43981 7785
rect 43981 7751 43982 7785
rect 43812 7677 43982 7751
rect 43812 7643 43813 7677
rect 43813 7643 43981 7677
rect 43981 7643 43982 7677
rect 43812 7642 43982 7643
rect 44184 7785 44354 7786
rect 44184 7751 44185 7785
rect 44185 7751 44353 7785
rect 44353 7751 44354 7785
rect 44184 7677 44354 7751
rect 44184 7643 44185 7677
rect 44185 7643 44353 7677
rect 44353 7643 44354 7677
rect 44184 7642 44354 7643
rect 44556 7785 44726 7786
rect 44556 7751 44557 7785
rect 44557 7751 44725 7785
rect 44725 7751 44726 7785
rect 44556 7677 44726 7751
rect 44556 7643 44557 7677
rect 44557 7643 44725 7677
rect 44725 7643 44726 7677
rect 44556 7642 44726 7643
rect 44928 7785 45098 7786
rect 44928 7751 44929 7785
rect 44929 7751 45097 7785
rect 45097 7751 45098 7785
rect 44928 7677 45098 7751
rect 44928 7643 44929 7677
rect 44929 7643 45097 7677
rect 45097 7643 45098 7677
rect 44928 7642 45098 7643
rect 39348 7149 39518 7162
rect 39348 7115 39349 7149
rect 39349 7115 39517 7149
rect 39517 7115 39518 7149
rect 39348 7102 39518 7115
rect 39720 7149 39890 7162
rect 39720 7115 39721 7149
rect 39721 7115 39889 7149
rect 39889 7115 39890 7149
rect 39720 7102 39890 7115
rect 40092 7149 40262 7162
rect 40092 7115 40093 7149
rect 40093 7115 40261 7149
rect 40261 7115 40262 7149
rect 40092 7102 40262 7115
rect 40464 7149 40634 7162
rect 40464 7115 40465 7149
rect 40465 7115 40633 7149
rect 40633 7115 40634 7149
rect 40464 7102 40634 7115
rect 40836 7149 41006 7162
rect 40836 7115 40837 7149
rect 40837 7115 41005 7149
rect 41005 7115 41006 7149
rect 40836 7102 41006 7115
rect 41208 7149 41378 7162
rect 41208 7115 41209 7149
rect 41209 7115 41377 7149
rect 41377 7115 41378 7149
rect 41208 7102 41378 7115
rect 41580 7149 41750 7162
rect 41580 7115 41581 7149
rect 41581 7115 41749 7149
rect 41749 7115 41750 7149
rect 41580 7102 41750 7115
rect 41952 7149 42122 7162
rect 41952 7115 41953 7149
rect 41953 7115 42121 7149
rect 42121 7115 42122 7149
rect 41952 7102 42122 7115
rect 42324 7149 42494 7162
rect 42324 7115 42325 7149
rect 42325 7115 42493 7149
rect 42493 7115 42494 7149
rect 42324 7102 42494 7115
rect 42696 7149 42866 7162
rect 42696 7115 42697 7149
rect 42697 7115 42865 7149
rect 42865 7115 42866 7149
rect 42696 7102 42866 7115
rect 43068 7149 43238 7162
rect 43068 7115 43069 7149
rect 43069 7115 43237 7149
rect 43237 7115 43238 7149
rect 43068 7102 43238 7115
rect 43440 7149 43610 7162
rect 43440 7115 43441 7149
rect 43441 7115 43609 7149
rect 43609 7115 43610 7149
rect 43440 7102 43610 7115
rect 43812 7149 43982 7162
rect 43812 7115 43813 7149
rect 43813 7115 43981 7149
rect 43981 7115 43982 7149
rect 43812 7102 43982 7115
rect 44184 7149 44354 7162
rect 44184 7115 44185 7149
rect 44185 7115 44353 7149
rect 44353 7115 44354 7149
rect 44184 7102 44354 7115
rect 45300 8949 45470 8962
rect 45300 8915 45301 8949
rect 45301 8915 45469 8949
rect 45469 8915 45470 8949
rect 45300 8902 45470 8915
rect 45672 8949 45842 8962
rect 45672 8915 45673 8949
rect 45673 8915 45841 8949
rect 45841 8915 45842 8949
rect 45672 8902 45842 8915
rect 46044 8949 46214 8962
rect 46044 8915 46045 8949
rect 46045 8915 46213 8949
rect 46213 8915 46214 8949
rect 46044 8902 46214 8915
rect 46416 8949 46586 8962
rect 46416 8915 46417 8949
rect 46417 8915 46585 8949
rect 46585 8915 46586 8949
rect 46416 8902 46586 8915
rect 46788 8949 46958 8962
rect 46788 8915 46789 8949
rect 46789 8915 46957 8949
rect 46957 8915 46958 8949
rect 46788 8902 46958 8915
rect 47160 8949 47330 8962
rect 47160 8915 47161 8949
rect 47161 8915 47329 8949
rect 47329 8915 47330 8949
rect 47160 8902 47330 8915
rect 47532 8949 47702 8962
rect 47532 8915 47533 8949
rect 47533 8915 47701 8949
rect 47701 8915 47702 8949
rect 47532 8902 47702 8915
rect 47904 8949 48074 8962
rect 47904 8915 47905 8949
rect 47905 8915 48073 8949
rect 48073 8915 48074 8949
rect 47904 8902 48074 8915
rect 48276 8949 48446 8962
rect 48276 8915 48277 8949
rect 48277 8915 48445 8949
rect 48445 8915 48446 8949
rect 48276 8902 48446 8915
rect 48648 8949 48818 8962
rect 48648 8915 48649 8949
rect 48649 8915 48817 8949
rect 48817 8915 48818 8949
rect 48648 8902 48818 8915
rect 49020 8949 49190 8962
rect 49020 8915 49021 8949
rect 49021 8915 49189 8949
rect 49189 8915 49190 8949
rect 49020 8902 49190 8915
rect 49392 8949 49562 8962
rect 49392 8915 49393 8949
rect 49393 8915 49561 8949
rect 49561 8915 49562 8949
rect 49392 8902 49562 8915
rect 49764 8949 49934 8962
rect 49764 8915 49765 8949
rect 49765 8915 49933 8949
rect 49933 8915 49934 8949
rect 49764 8902 49934 8915
rect 50136 8949 50306 8962
rect 50136 8915 50137 8949
rect 50137 8915 50305 8949
rect 50305 8915 50306 8949
rect 50136 8902 50306 8915
rect 50508 8949 50678 8962
rect 50508 8915 50509 8949
rect 50509 8915 50677 8949
rect 50677 8915 50678 8949
rect 50508 8902 50678 8915
rect 50880 8949 51050 8962
rect 50880 8915 50881 8949
rect 50881 8915 51049 8949
rect 51049 8915 51050 8949
rect 50880 8902 51050 8915
rect 45300 8421 45470 8422
rect 45300 8387 45301 8421
rect 45301 8387 45469 8421
rect 45469 8387 45470 8421
rect 45300 8313 45470 8387
rect 45300 8279 45301 8313
rect 45301 8279 45469 8313
rect 45469 8279 45470 8313
rect 45300 8278 45470 8279
rect 45672 8421 45842 8422
rect 45672 8387 45673 8421
rect 45673 8387 45841 8421
rect 45841 8387 45842 8421
rect 45672 8313 45842 8387
rect 45672 8279 45673 8313
rect 45673 8279 45841 8313
rect 45841 8279 45842 8313
rect 45672 8278 45842 8279
rect 46044 8421 46214 8422
rect 46044 8387 46045 8421
rect 46045 8387 46213 8421
rect 46213 8387 46214 8421
rect 46044 8313 46214 8387
rect 46044 8279 46045 8313
rect 46045 8279 46213 8313
rect 46213 8279 46214 8313
rect 46044 8278 46214 8279
rect 46416 8421 46586 8422
rect 46416 8387 46417 8421
rect 46417 8387 46585 8421
rect 46585 8387 46586 8421
rect 46416 8313 46586 8387
rect 46416 8279 46417 8313
rect 46417 8279 46585 8313
rect 46585 8279 46586 8313
rect 46416 8278 46586 8279
rect 46788 8421 46958 8422
rect 46788 8387 46789 8421
rect 46789 8387 46957 8421
rect 46957 8387 46958 8421
rect 46788 8313 46958 8387
rect 46788 8279 46789 8313
rect 46789 8279 46957 8313
rect 46957 8279 46958 8313
rect 46788 8278 46958 8279
rect 47160 8421 47330 8422
rect 47160 8387 47161 8421
rect 47161 8387 47329 8421
rect 47329 8387 47330 8421
rect 47160 8313 47330 8387
rect 47160 8279 47161 8313
rect 47161 8279 47329 8313
rect 47329 8279 47330 8313
rect 47160 8278 47330 8279
rect 47532 8421 47702 8422
rect 47532 8387 47533 8421
rect 47533 8387 47701 8421
rect 47701 8387 47702 8421
rect 47532 8313 47702 8387
rect 47532 8279 47533 8313
rect 47533 8279 47701 8313
rect 47701 8279 47702 8313
rect 47532 8278 47702 8279
rect 47904 8421 48074 8422
rect 47904 8387 47905 8421
rect 47905 8387 48073 8421
rect 48073 8387 48074 8421
rect 47904 8313 48074 8387
rect 47904 8279 47905 8313
rect 47905 8279 48073 8313
rect 48073 8279 48074 8313
rect 47904 8278 48074 8279
rect 48276 8421 48446 8422
rect 48276 8387 48277 8421
rect 48277 8387 48445 8421
rect 48445 8387 48446 8421
rect 48276 8313 48446 8387
rect 48276 8279 48277 8313
rect 48277 8279 48445 8313
rect 48445 8279 48446 8313
rect 48276 8278 48446 8279
rect 48648 8421 48818 8422
rect 48648 8387 48649 8421
rect 48649 8387 48817 8421
rect 48817 8387 48818 8421
rect 48648 8313 48818 8387
rect 48648 8279 48649 8313
rect 48649 8279 48817 8313
rect 48817 8279 48818 8313
rect 48648 8278 48818 8279
rect 49020 8421 49190 8422
rect 49020 8387 49021 8421
rect 49021 8387 49189 8421
rect 49189 8387 49190 8421
rect 49020 8313 49190 8387
rect 49020 8279 49021 8313
rect 49021 8279 49189 8313
rect 49189 8279 49190 8313
rect 49020 8278 49190 8279
rect 49392 8421 49562 8422
rect 49392 8387 49393 8421
rect 49393 8387 49561 8421
rect 49561 8387 49562 8421
rect 49392 8313 49562 8387
rect 49392 8279 49393 8313
rect 49393 8279 49561 8313
rect 49561 8279 49562 8313
rect 49392 8278 49562 8279
rect 49764 8421 49934 8422
rect 49764 8387 49765 8421
rect 49765 8387 49933 8421
rect 49933 8387 49934 8421
rect 49764 8313 49934 8387
rect 49764 8279 49765 8313
rect 49765 8279 49933 8313
rect 49933 8279 49934 8313
rect 49764 8278 49934 8279
rect 50136 8421 50306 8422
rect 50136 8387 50137 8421
rect 50137 8387 50305 8421
rect 50305 8387 50306 8421
rect 50136 8313 50306 8387
rect 50136 8279 50137 8313
rect 50137 8279 50305 8313
rect 50305 8279 50306 8313
rect 50136 8278 50306 8279
rect 50508 8421 50678 8422
rect 50508 8387 50509 8421
rect 50509 8387 50677 8421
rect 50677 8387 50678 8421
rect 50508 8313 50678 8387
rect 50508 8279 50509 8313
rect 50509 8279 50677 8313
rect 50677 8279 50678 8313
rect 50508 8278 50678 8279
rect 50880 8421 51050 8422
rect 50880 8387 50881 8421
rect 50881 8387 51049 8421
rect 51049 8387 51050 8421
rect 50880 8313 51050 8387
rect 50880 8279 50881 8313
rect 50881 8279 51049 8313
rect 51049 8279 51050 8313
rect 50880 8278 51050 8279
rect 45300 7785 45470 7786
rect 45300 7751 45301 7785
rect 45301 7751 45469 7785
rect 45469 7751 45470 7785
rect 45300 7677 45470 7751
rect 45300 7643 45301 7677
rect 45301 7643 45469 7677
rect 45469 7643 45470 7677
rect 45300 7642 45470 7643
rect 45672 7785 45842 7786
rect 45672 7751 45673 7785
rect 45673 7751 45841 7785
rect 45841 7751 45842 7785
rect 45672 7677 45842 7751
rect 45672 7643 45673 7677
rect 45673 7643 45841 7677
rect 45841 7643 45842 7677
rect 45672 7642 45842 7643
rect 46044 7785 46214 7786
rect 46044 7751 46045 7785
rect 46045 7751 46213 7785
rect 46213 7751 46214 7785
rect 46044 7677 46214 7751
rect 46044 7643 46045 7677
rect 46045 7643 46213 7677
rect 46213 7643 46214 7677
rect 46044 7642 46214 7643
rect 46416 7785 46586 7786
rect 46416 7751 46417 7785
rect 46417 7751 46585 7785
rect 46585 7751 46586 7785
rect 46416 7677 46586 7751
rect 46416 7643 46417 7677
rect 46417 7643 46585 7677
rect 46585 7643 46586 7677
rect 46416 7642 46586 7643
rect 46788 7785 46958 7786
rect 46788 7751 46789 7785
rect 46789 7751 46957 7785
rect 46957 7751 46958 7785
rect 46788 7677 46958 7751
rect 46788 7643 46789 7677
rect 46789 7643 46957 7677
rect 46957 7643 46958 7677
rect 46788 7642 46958 7643
rect 47160 7785 47330 7786
rect 47160 7751 47161 7785
rect 47161 7751 47329 7785
rect 47329 7751 47330 7785
rect 47160 7677 47330 7751
rect 47160 7643 47161 7677
rect 47161 7643 47329 7677
rect 47329 7643 47330 7677
rect 47160 7642 47330 7643
rect 47532 7785 47702 7786
rect 47532 7751 47533 7785
rect 47533 7751 47701 7785
rect 47701 7751 47702 7785
rect 47532 7677 47702 7751
rect 47532 7643 47533 7677
rect 47533 7643 47701 7677
rect 47701 7643 47702 7677
rect 47532 7642 47702 7643
rect 47904 7785 48074 7786
rect 47904 7751 47905 7785
rect 47905 7751 48073 7785
rect 48073 7751 48074 7785
rect 47904 7677 48074 7751
rect 47904 7643 47905 7677
rect 47905 7643 48073 7677
rect 48073 7643 48074 7677
rect 47904 7642 48074 7643
rect 48276 7785 48446 7786
rect 48276 7751 48277 7785
rect 48277 7751 48445 7785
rect 48445 7751 48446 7785
rect 48276 7677 48446 7751
rect 48276 7643 48277 7677
rect 48277 7643 48445 7677
rect 48445 7643 48446 7677
rect 48276 7642 48446 7643
rect 48648 7785 48818 7786
rect 48648 7751 48649 7785
rect 48649 7751 48817 7785
rect 48817 7751 48818 7785
rect 48648 7677 48818 7751
rect 48648 7643 48649 7677
rect 48649 7643 48817 7677
rect 48817 7643 48818 7677
rect 48648 7642 48818 7643
rect 49020 7785 49190 7786
rect 49020 7751 49021 7785
rect 49021 7751 49189 7785
rect 49189 7751 49190 7785
rect 49020 7677 49190 7751
rect 49020 7643 49021 7677
rect 49021 7643 49189 7677
rect 49189 7643 49190 7677
rect 49020 7642 49190 7643
rect 49392 7785 49562 7786
rect 49392 7751 49393 7785
rect 49393 7751 49561 7785
rect 49561 7751 49562 7785
rect 49392 7677 49562 7751
rect 49392 7643 49393 7677
rect 49393 7643 49561 7677
rect 49561 7643 49562 7677
rect 49392 7642 49562 7643
rect 49764 7785 49934 7786
rect 49764 7751 49765 7785
rect 49765 7751 49933 7785
rect 49933 7751 49934 7785
rect 49764 7677 49934 7751
rect 49764 7643 49765 7677
rect 49765 7643 49933 7677
rect 49933 7643 49934 7677
rect 49764 7642 49934 7643
rect 50136 7785 50306 7786
rect 50136 7751 50137 7785
rect 50137 7751 50305 7785
rect 50305 7751 50306 7785
rect 50136 7677 50306 7751
rect 50136 7643 50137 7677
rect 50137 7643 50305 7677
rect 50305 7643 50306 7677
rect 50136 7642 50306 7643
rect 50508 7785 50678 7786
rect 50508 7751 50509 7785
rect 50509 7751 50677 7785
rect 50677 7751 50678 7785
rect 50508 7677 50678 7751
rect 50508 7643 50509 7677
rect 50509 7643 50677 7677
rect 50677 7643 50678 7677
rect 50508 7642 50678 7643
rect 50880 7785 51050 7786
rect 50880 7751 50881 7785
rect 50881 7751 51049 7785
rect 51049 7751 51050 7785
rect 50880 7677 51050 7751
rect 50880 7643 50881 7677
rect 50881 7643 51049 7677
rect 51049 7643 51050 7677
rect 50880 7642 51050 7643
rect 44556 7149 44726 7162
rect 44556 7115 44557 7149
rect 44557 7115 44725 7149
rect 44725 7115 44726 7149
rect 44556 7102 44726 7115
rect 44928 7149 45098 7162
rect 44928 7115 44929 7149
rect 44929 7115 45097 7149
rect 45097 7115 45098 7149
rect 44928 7102 45098 7115
rect 45300 7149 45470 7162
rect 45300 7115 45301 7149
rect 45301 7115 45469 7149
rect 45469 7115 45470 7149
rect 45300 7102 45470 7115
rect 40122 6401 40404 6675
rect 40836 6561 41006 6576
rect 40836 6527 40837 6561
rect 40837 6527 41005 6561
rect 41005 6527 41006 6561
rect 40836 6512 41006 6527
rect 41208 6561 41378 6576
rect 41208 6527 41209 6561
rect 41209 6527 41377 6561
rect 41377 6527 41378 6561
rect 41208 6512 41378 6527
rect 41580 6561 41750 6576
rect 41580 6527 41581 6561
rect 41581 6527 41749 6561
rect 41749 6527 41750 6561
rect 41580 6512 41750 6527
rect 41952 6561 42122 6576
rect 41952 6527 41953 6561
rect 41953 6527 42121 6561
rect 42121 6527 42122 6561
rect 41952 6512 42122 6527
rect 42324 6561 42494 6576
rect 42324 6527 42325 6561
rect 42325 6527 42493 6561
rect 42493 6527 42494 6561
rect 42324 6512 42494 6527
rect 42696 6561 42866 6576
rect 42696 6527 42697 6561
rect 42697 6527 42865 6561
rect 42865 6527 42866 6561
rect 42696 6512 42866 6527
rect 43068 6561 43238 6576
rect 43068 6527 43069 6561
rect 43069 6527 43237 6561
rect 43237 6527 43238 6561
rect 43068 6512 43238 6527
rect 43440 6561 43610 6576
rect 43440 6527 43441 6561
rect 43441 6527 43609 6561
rect 43609 6527 43610 6561
rect 43440 6512 43610 6527
rect 44616 6557 44898 6831
rect 45672 7149 45842 7162
rect 45672 7115 45673 7149
rect 45673 7115 45841 7149
rect 45841 7115 45842 7149
rect 45672 7102 45842 7115
rect 46044 7149 46214 7162
rect 46044 7115 46045 7149
rect 46045 7115 46213 7149
rect 46213 7115 46214 7149
rect 46044 7102 46214 7115
rect 46416 7149 46586 7162
rect 46416 7115 46417 7149
rect 46417 7115 46585 7149
rect 46585 7115 46586 7149
rect 46416 7102 46586 7115
rect 46788 7149 46958 7162
rect 46788 7115 46789 7149
rect 46789 7115 46957 7149
rect 46957 7115 46958 7149
rect 46788 7102 46958 7115
rect 47160 7149 47330 7162
rect 47160 7115 47161 7149
rect 47161 7115 47329 7149
rect 47329 7115 47330 7149
rect 47160 7102 47330 7115
rect 47532 7149 47702 7162
rect 47532 7115 47533 7149
rect 47533 7115 47701 7149
rect 47701 7115 47702 7149
rect 47532 7102 47702 7115
rect 47904 7149 48074 7162
rect 47904 7115 47905 7149
rect 47905 7115 48073 7149
rect 48073 7115 48074 7149
rect 47904 7102 48074 7115
rect 48276 7149 48446 7162
rect 48276 7115 48277 7149
rect 48277 7115 48445 7149
rect 48445 7115 48446 7149
rect 48276 7102 48446 7115
rect 48648 7149 48818 7162
rect 48648 7115 48649 7149
rect 48649 7115 48817 7149
rect 48817 7115 48818 7149
rect 48648 7102 48818 7115
rect 49020 7149 49190 7162
rect 49020 7115 49021 7149
rect 49021 7115 49189 7149
rect 49189 7115 49190 7149
rect 49020 7102 49190 7115
rect 49392 7149 49562 7162
rect 49392 7115 49393 7149
rect 49393 7115 49561 7149
rect 49561 7115 49562 7149
rect 49392 7102 49562 7115
rect 49764 7149 49934 7162
rect 49764 7115 49765 7149
rect 49765 7115 49933 7149
rect 49933 7115 49934 7149
rect 49764 7102 49934 7115
rect 50136 7149 50306 7162
rect 50136 7115 50137 7149
rect 50137 7115 50305 7149
rect 50305 7115 50306 7149
rect 50136 7102 50306 7115
rect 50508 7149 50678 7162
rect 50508 7115 50509 7149
rect 50509 7115 50677 7149
rect 50677 7115 50678 7149
rect 50508 7102 50678 7115
rect 50880 7149 51050 7162
rect 50880 7115 50881 7149
rect 50881 7115 51049 7149
rect 51049 7115 51050 7149
rect 50880 7102 51050 7115
rect 40246 6109 40392 6259
rect 40246 5709 40392 5859
rect 45432 6522 45714 6794
rect 46176 6522 46458 6794
rect 46920 6522 47202 6794
rect 47664 6522 47946 6794
rect 48408 6522 48690 6794
rect 49152 6522 49434 6794
rect 49896 6522 50178 6794
rect 50640 6522 50922 6794
rect 40246 5309 40392 5459
rect 40836 5633 41006 5634
rect 40836 5599 40837 5633
rect 40837 5599 41005 5633
rect 41005 5599 41006 5633
rect 40836 5525 41006 5599
rect 40836 5491 40837 5525
rect 40837 5491 41005 5525
rect 41005 5491 41006 5525
rect 40836 5490 41006 5491
rect 41208 5633 41378 5634
rect 41208 5599 41209 5633
rect 41209 5599 41377 5633
rect 41377 5599 41378 5633
rect 41208 5525 41378 5599
rect 41208 5491 41209 5525
rect 41209 5491 41377 5525
rect 41377 5491 41378 5525
rect 41208 5490 41378 5491
rect 41580 5633 41750 5634
rect 41580 5599 41581 5633
rect 41581 5599 41749 5633
rect 41749 5599 41750 5633
rect 41580 5525 41750 5599
rect 41580 5491 41581 5525
rect 41581 5491 41749 5525
rect 41749 5491 41750 5525
rect 41580 5490 41750 5491
rect 41952 5633 42122 5634
rect 41952 5599 41953 5633
rect 41953 5599 42121 5633
rect 42121 5599 42122 5633
rect 41952 5525 42122 5599
rect 41952 5491 41953 5525
rect 41953 5491 42121 5525
rect 42121 5491 42122 5525
rect 41952 5490 42122 5491
rect 42324 5633 42494 5634
rect 42324 5599 42325 5633
rect 42325 5599 42493 5633
rect 42493 5599 42494 5633
rect 42324 5525 42494 5599
rect 42324 5491 42325 5525
rect 42325 5491 42493 5525
rect 42493 5491 42494 5525
rect 42324 5490 42494 5491
rect 42696 5633 42866 5634
rect 42696 5599 42697 5633
rect 42697 5599 42865 5633
rect 42865 5599 42866 5633
rect 42696 5525 42866 5599
rect 42696 5491 42697 5525
rect 42697 5491 42865 5525
rect 42865 5491 42866 5525
rect 42696 5490 42866 5491
rect 43068 5633 43238 5634
rect 43068 5599 43069 5633
rect 43069 5599 43237 5633
rect 43237 5599 43238 5633
rect 43068 5525 43238 5599
rect 43068 5491 43069 5525
rect 43069 5491 43237 5525
rect 43237 5491 43238 5525
rect 43068 5490 43238 5491
rect 43440 5633 43610 5634
rect 43440 5599 43441 5633
rect 43441 5599 43609 5633
rect 43609 5599 43610 5633
rect 43440 5525 43610 5599
rect 43440 5491 43441 5525
rect 43441 5491 43609 5525
rect 43609 5491 43610 5525
rect 43440 5490 43610 5491
rect 44162 5569 44308 5719
rect 45638 5635 46122 6135
rect 40246 4909 40392 5059
rect 44162 5169 44308 5319
rect 44162 4769 44308 4919
rect 45852 4748 46134 5020
rect 40836 4597 41006 4598
rect 40836 4563 40837 4597
rect 40837 4563 41005 4597
rect 41005 4563 41006 4597
rect 40836 4489 41006 4563
rect 40836 4455 40837 4489
rect 40837 4455 41005 4489
rect 41005 4455 41006 4489
rect 40836 4454 41006 4455
rect 41208 4597 41378 4598
rect 41208 4563 41209 4597
rect 41209 4563 41377 4597
rect 41377 4563 41378 4597
rect 41208 4489 41378 4563
rect 41208 4455 41209 4489
rect 41209 4455 41377 4489
rect 41377 4455 41378 4489
rect 41208 4454 41378 4455
rect 41580 4597 41750 4598
rect 41580 4563 41581 4597
rect 41581 4563 41749 4597
rect 41749 4563 41750 4597
rect 41580 4489 41750 4563
rect 41580 4455 41581 4489
rect 41581 4455 41749 4489
rect 41749 4455 41750 4489
rect 41580 4454 41750 4455
rect 41952 4597 42122 4598
rect 41952 4563 41953 4597
rect 41953 4563 42121 4597
rect 42121 4563 42122 4597
rect 41952 4489 42122 4563
rect 41952 4455 41953 4489
rect 41953 4455 42121 4489
rect 42121 4455 42122 4489
rect 41952 4454 42122 4455
rect 42324 4597 42494 4598
rect 42324 4563 42325 4597
rect 42325 4563 42493 4597
rect 42493 4563 42494 4597
rect 42324 4489 42494 4563
rect 42324 4455 42325 4489
rect 42325 4455 42493 4489
rect 42493 4455 42494 4489
rect 42324 4454 42494 4455
rect 42696 4597 42866 4598
rect 42696 4563 42697 4597
rect 42697 4563 42865 4597
rect 42865 4563 42866 4597
rect 42696 4489 42866 4563
rect 42696 4455 42697 4489
rect 42697 4455 42865 4489
rect 42865 4455 42866 4489
rect 42696 4454 42866 4455
rect 43068 4597 43238 4598
rect 43068 4563 43069 4597
rect 43069 4563 43237 4597
rect 43237 4563 43238 4597
rect 43068 4489 43238 4563
rect 43068 4455 43069 4489
rect 43069 4455 43237 4489
rect 43237 4455 43238 4489
rect 43068 4454 43238 4455
rect 43440 4597 43610 4598
rect 43440 4563 43441 4597
rect 43441 4563 43609 4597
rect 43609 4563 43610 4597
rect 43440 4489 43610 4563
rect 43440 4455 43441 4489
rect 43441 4455 43609 4489
rect 43609 4455 43610 4489
rect 43440 4454 43610 4455
rect 44162 4369 44308 4519
rect 45556 4132 45730 4306
rect 45556 3732 45730 3906
rect 40836 3561 41006 3562
rect 40836 3527 40837 3561
rect 40837 3527 41005 3561
rect 41005 3527 41006 3561
rect 40836 3453 41006 3527
rect 40836 3419 40837 3453
rect 40837 3419 41005 3453
rect 41005 3419 41006 3453
rect 40836 3418 41006 3419
rect 41208 3561 41378 3562
rect 41208 3527 41209 3561
rect 41209 3527 41377 3561
rect 41377 3527 41378 3561
rect 41208 3453 41378 3527
rect 41208 3419 41209 3453
rect 41209 3419 41377 3453
rect 41377 3419 41378 3453
rect 41208 3418 41378 3419
rect 41580 3561 41750 3562
rect 41580 3527 41581 3561
rect 41581 3527 41749 3561
rect 41749 3527 41750 3561
rect 41580 3453 41750 3527
rect 41580 3419 41581 3453
rect 41581 3419 41749 3453
rect 41749 3419 41750 3453
rect 41580 3418 41750 3419
rect 41952 3561 42122 3562
rect 41952 3527 41953 3561
rect 41953 3527 42121 3561
rect 42121 3527 42122 3561
rect 41952 3453 42122 3527
rect 41952 3419 41953 3453
rect 41953 3419 42121 3453
rect 42121 3419 42122 3453
rect 41952 3418 42122 3419
rect 42324 3561 42494 3562
rect 42324 3527 42325 3561
rect 42325 3527 42493 3561
rect 42493 3527 42494 3561
rect 42324 3453 42494 3527
rect 42324 3419 42325 3453
rect 42325 3419 42493 3453
rect 42493 3419 42494 3453
rect 42324 3418 42494 3419
rect 42696 3561 42866 3562
rect 42696 3527 42697 3561
rect 42697 3527 42865 3561
rect 42865 3527 42866 3561
rect 42696 3453 42866 3527
rect 42696 3419 42697 3453
rect 42697 3419 42865 3453
rect 42865 3419 42866 3453
rect 42696 3418 42866 3419
rect 43068 3561 43238 3562
rect 43068 3527 43069 3561
rect 43069 3527 43237 3561
rect 43237 3527 43238 3561
rect 43068 3453 43238 3527
rect 43068 3419 43069 3453
rect 43069 3419 43237 3453
rect 43237 3419 43238 3453
rect 43068 3418 43238 3419
rect 43440 3561 43610 3562
rect 43440 3527 43441 3561
rect 43441 3527 43609 3561
rect 43609 3527 43610 3561
rect 43440 3453 43610 3527
rect 43440 3419 43441 3453
rect 43441 3419 43609 3453
rect 43609 3419 43610 3453
rect 43440 3418 43610 3419
rect 45556 3332 45730 3506
rect 40836 2525 41006 2536
rect 40836 2491 40837 2525
rect 40837 2491 41005 2525
rect 41005 2491 41006 2525
rect 40836 2482 41006 2491
rect 41208 2525 41378 2536
rect 41208 2491 41209 2525
rect 41209 2491 41377 2525
rect 41377 2491 41378 2525
rect 41208 2482 41378 2491
rect 41580 2525 41750 2536
rect 41580 2491 41581 2525
rect 41581 2491 41749 2525
rect 41749 2491 41750 2525
rect 41580 2482 41750 2491
rect 41952 2525 42122 2536
rect 41952 2491 41953 2525
rect 41953 2491 42121 2525
rect 42121 2491 42122 2525
rect 41952 2482 42122 2491
rect 42324 2525 42494 2536
rect 42324 2491 42325 2525
rect 42325 2491 42493 2525
rect 42493 2491 42494 2525
rect 42324 2482 42494 2491
rect 42696 2525 42866 2536
rect 42696 2491 42697 2525
rect 42697 2491 42865 2525
rect 42865 2491 42866 2525
rect 42696 2482 42866 2491
rect 43068 2525 43238 2536
rect 43068 2491 43069 2525
rect 43069 2491 43237 2525
rect 43237 2491 43238 2525
rect 43068 2482 43238 2491
rect 41816 2016 42630 2196
rect 40836 1867 41006 1878
rect 40836 1833 40837 1867
rect 40837 1833 41005 1867
rect 41005 1833 41006 1867
rect 40836 1822 41006 1833
rect 41208 1867 41378 1878
rect 41208 1833 41209 1867
rect 41209 1833 41377 1867
rect 41377 1833 41378 1867
rect 41208 1822 41378 1833
rect 41580 1867 41750 1878
rect 41580 1833 41581 1867
rect 41581 1833 41749 1867
rect 41749 1833 41750 1867
rect 41580 1822 41750 1833
rect 41952 1867 42122 1878
rect 41952 1833 41953 1867
rect 41953 1833 42121 1867
rect 42121 1833 42122 1867
rect 41952 1822 42122 1833
rect 42324 1867 42494 1878
rect 42324 1833 42325 1867
rect 42325 1833 42493 1867
rect 42493 1833 42494 1867
rect 42324 1822 42494 1833
rect 43440 2525 43610 2536
rect 43440 2491 43441 2525
rect 43441 2491 43609 2525
rect 43609 2491 43610 2525
rect 43440 2482 43610 2491
rect 43942 2340 44224 2612
rect 44686 2340 44968 2612
rect 45430 2340 45712 2612
rect 42696 1867 42866 1878
rect 42696 1833 42697 1867
rect 42697 1833 42865 1867
rect 42865 1833 42866 1867
rect 42696 1822 42866 1833
rect 43068 1867 43238 1878
rect 43068 1833 43069 1867
rect 43069 1833 43237 1867
rect 43237 1833 43238 1867
rect 43068 1822 43238 1833
rect 43440 1867 43610 1878
rect 43440 1833 43441 1867
rect 43441 1833 43609 1867
rect 43609 1833 43610 1867
rect 43440 1822 43610 1833
rect 43812 1867 43982 1878
rect 43812 1833 43813 1867
rect 43813 1833 43981 1867
rect 43981 1833 43982 1867
rect 43812 1822 43982 1833
rect 44184 1867 44354 1878
rect 44184 1833 44185 1867
rect 44185 1833 44353 1867
rect 44353 1833 44354 1867
rect 44184 1822 44354 1833
rect 44556 1867 44726 1878
rect 44556 1833 44557 1867
rect 44557 1833 44725 1867
rect 44725 1833 44726 1867
rect 44556 1822 44726 1833
rect 44928 1867 45098 1878
rect 44928 1833 44929 1867
rect 44929 1833 45097 1867
rect 45097 1833 45098 1867
rect 44928 1822 45098 1833
rect 45300 1867 45470 1878
rect 45300 1833 45301 1867
rect 45301 1833 45469 1867
rect 45469 1833 45470 1867
rect 45300 1822 45470 1833
rect 46174 2340 46456 2612
rect 46918 2340 47200 2612
rect 47662 2340 47944 2612
rect 48406 2340 48688 2612
rect 49150 2340 49432 2612
rect 45826 2050 46104 2324
rect 45672 1867 45842 1878
rect 45672 1833 45673 1867
rect 45673 1833 45841 1867
rect 45841 1833 45842 1867
rect 45672 1822 45842 1833
rect 46044 1867 46214 1878
rect 46044 1833 46045 1867
rect 46045 1833 46213 1867
rect 46213 1833 46214 1867
rect 46044 1822 46214 1833
rect 46416 1867 46586 1878
rect 46416 1833 46417 1867
rect 46417 1833 46585 1867
rect 46585 1833 46586 1867
rect 46416 1822 46586 1833
rect 46788 1867 46958 1878
rect 46788 1833 46789 1867
rect 46789 1833 46957 1867
rect 46957 1833 46958 1867
rect 46788 1822 46958 1833
rect 47160 1867 47330 1878
rect 47160 1833 47161 1867
rect 47161 1833 47329 1867
rect 47329 1833 47330 1867
rect 47160 1822 47330 1833
rect 47532 1867 47702 1878
rect 47532 1833 47533 1867
rect 47533 1833 47701 1867
rect 47701 1833 47702 1867
rect 47532 1822 47702 1833
rect 47904 1867 48074 1878
rect 47904 1833 47905 1867
rect 47905 1833 48073 1867
rect 48073 1833 48074 1867
rect 47904 1822 48074 1833
rect 48276 1867 48446 1878
rect 48276 1833 48277 1867
rect 48277 1833 48445 1867
rect 48445 1833 48446 1867
rect 48276 1822 48446 1833
rect 48648 1867 48818 1878
rect 48648 1833 48649 1867
rect 48649 1833 48817 1867
rect 48817 1833 48818 1867
rect 48648 1822 48818 1833
rect 49020 1867 49190 1878
rect 49020 1833 49021 1867
rect 49021 1833 49189 1867
rect 49189 1833 49190 1867
rect 49020 1822 49190 1833
rect 49392 1867 49562 1878
rect 49392 1833 49393 1867
rect 49393 1833 49561 1867
rect 49561 1833 49562 1867
rect 49392 1822 49562 1833
rect 40836 1557 41006 1558
rect 40836 1523 40837 1557
rect 40837 1523 41005 1557
rect 41005 1523 41006 1557
rect 40836 1449 41006 1523
rect 40836 1415 40837 1449
rect 40837 1415 41005 1449
rect 41005 1415 41006 1449
rect 40836 1414 41006 1415
rect 41208 1557 41378 1558
rect 41208 1523 41209 1557
rect 41209 1523 41377 1557
rect 41377 1523 41378 1557
rect 41208 1449 41378 1523
rect 41208 1415 41209 1449
rect 41209 1415 41377 1449
rect 41377 1415 41378 1449
rect 41208 1414 41378 1415
rect 41580 1557 41750 1558
rect 41580 1523 41581 1557
rect 41581 1523 41749 1557
rect 41749 1523 41750 1557
rect 41580 1449 41750 1523
rect 41580 1415 41581 1449
rect 41581 1415 41749 1449
rect 41749 1415 41750 1449
rect 41580 1414 41750 1415
rect 41952 1557 42122 1558
rect 41952 1523 41953 1557
rect 41953 1523 42121 1557
rect 42121 1523 42122 1557
rect 41952 1449 42122 1523
rect 41952 1415 41953 1449
rect 41953 1415 42121 1449
rect 42121 1415 42122 1449
rect 41952 1414 42122 1415
rect 42324 1557 42494 1558
rect 42324 1523 42325 1557
rect 42325 1523 42493 1557
rect 42493 1523 42494 1557
rect 42324 1449 42494 1523
rect 42324 1415 42325 1449
rect 42325 1415 42493 1449
rect 42493 1415 42494 1449
rect 42324 1414 42494 1415
rect 42696 1557 42866 1558
rect 42696 1523 42697 1557
rect 42697 1523 42865 1557
rect 42865 1523 42866 1557
rect 42696 1449 42866 1523
rect 42696 1415 42697 1449
rect 42697 1415 42865 1449
rect 42865 1415 42866 1449
rect 42696 1414 42866 1415
rect 43068 1557 43238 1558
rect 43068 1523 43069 1557
rect 43069 1523 43237 1557
rect 43237 1523 43238 1557
rect 43068 1449 43238 1523
rect 43068 1415 43069 1449
rect 43069 1415 43237 1449
rect 43237 1415 43238 1449
rect 43068 1414 43238 1415
rect 43440 1557 43610 1558
rect 43440 1523 43441 1557
rect 43441 1523 43609 1557
rect 43609 1523 43610 1557
rect 43440 1449 43610 1523
rect 43440 1415 43441 1449
rect 43441 1415 43609 1449
rect 43609 1415 43610 1449
rect 43440 1414 43610 1415
rect 43812 1557 43982 1558
rect 43812 1523 43813 1557
rect 43813 1523 43981 1557
rect 43981 1523 43982 1557
rect 43812 1449 43982 1523
rect 43812 1415 43813 1449
rect 43813 1415 43981 1449
rect 43981 1415 43982 1449
rect 43812 1414 43982 1415
rect 44184 1557 44354 1558
rect 44184 1523 44185 1557
rect 44185 1523 44353 1557
rect 44353 1523 44354 1557
rect 44184 1449 44354 1523
rect 44184 1415 44185 1449
rect 44185 1415 44353 1449
rect 44353 1415 44354 1449
rect 44184 1414 44354 1415
rect 44556 1557 44726 1558
rect 44556 1523 44557 1557
rect 44557 1523 44725 1557
rect 44725 1523 44726 1557
rect 44556 1449 44726 1523
rect 44556 1415 44557 1449
rect 44557 1415 44725 1449
rect 44725 1415 44726 1449
rect 44556 1414 44726 1415
rect 44928 1557 45098 1558
rect 44928 1523 44929 1557
rect 44929 1523 45097 1557
rect 45097 1523 45098 1557
rect 44928 1449 45098 1523
rect 44928 1415 44929 1449
rect 44929 1415 45097 1449
rect 45097 1415 45098 1449
rect 44928 1414 45098 1415
rect 45300 1557 45470 1558
rect 45300 1523 45301 1557
rect 45301 1523 45469 1557
rect 45469 1523 45470 1557
rect 45300 1449 45470 1523
rect 45300 1415 45301 1449
rect 45301 1415 45469 1449
rect 45469 1415 45470 1449
rect 45300 1414 45470 1415
rect 45672 1557 45842 1558
rect 45672 1523 45673 1557
rect 45673 1523 45841 1557
rect 45841 1523 45842 1557
rect 45672 1449 45842 1523
rect 45672 1415 45673 1449
rect 45673 1415 45841 1449
rect 45841 1415 45842 1449
rect 45672 1414 45842 1415
rect 46044 1557 46214 1558
rect 46044 1523 46045 1557
rect 46045 1523 46213 1557
rect 46213 1523 46214 1557
rect 46044 1449 46214 1523
rect 46044 1415 46045 1449
rect 46045 1415 46213 1449
rect 46213 1415 46214 1449
rect 46044 1414 46214 1415
rect 46416 1557 46586 1558
rect 46416 1523 46417 1557
rect 46417 1523 46585 1557
rect 46585 1523 46586 1557
rect 46416 1449 46586 1523
rect 46416 1415 46417 1449
rect 46417 1415 46585 1449
rect 46585 1415 46586 1449
rect 46416 1414 46586 1415
rect 46788 1557 46958 1558
rect 46788 1523 46789 1557
rect 46789 1523 46957 1557
rect 46957 1523 46958 1557
rect 46788 1449 46958 1523
rect 46788 1415 46789 1449
rect 46789 1415 46957 1449
rect 46957 1415 46958 1449
rect 46788 1414 46958 1415
rect 47160 1557 47330 1558
rect 47160 1523 47161 1557
rect 47161 1523 47329 1557
rect 47329 1523 47330 1557
rect 47160 1449 47330 1523
rect 47160 1415 47161 1449
rect 47161 1415 47329 1449
rect 47329 1415 47330 1449
rect 47160 1414 47330 1415
rect 47532 1557 47702 1558
rect 47532 1523 47533 1557
rect 47533 1523 47701 1557
rect 47701 1523 47702 1557
rect 47532 1449 47702 1523
rect 47532 1415 47533 1449
rect 47533 1415 47701 1449
rect 47701 1415 47702 1449
rect 47532 1414 47702 1415
rect 47904 1557 48074 1558
rect 47904 1523 47905 1557
rect 47905 1523 48073 1557
rect 48073 1523 48074 1557
rect 47904 1449 48074 1523
rect 47904 1415 47905 1449
rect 47905 1415 48073 1449
rect 48073 1415 48074 1449
rect 47904 1414 48074 1415
rect 48276 1557 48446 1558
rect 48276 1523 48277 1557
rect 48277 1523 48445 1557
rect 48445 1523 48446 1557
rect 48276 1449 48446 1523
rect 48276 1415 48277 1449
rect 48277 1415 48445 1449
rect 48445 1415 48446 1449
rect 48276 1414 48446 1415
rect 48648 1557 48818 1558
rect 48648 1523 48649 1557
rect 48649 1523 48817 1557
rect 48817 1523 48818 1557
rect 48648 1449 48818 1523
rect 48648 1415 48649 1449
rect 48649 1415 48817 1449
rect 48817 1415 48818 1449
rect 48648 1414 48818 1415
rect 49020 1557 49190 1558
rect 49020 1523 49021 1557
rect 49021 1523 49189 1557
rect 49189 1523 49190 1557
rect 49020 1449 49190 1523
rect 49020 1415 49021 1449
rect 49021 1415 49189 1449
rect 49189 1415 49190 1449
rect 49020 1414 49190 1415
rect 49392 1557 49562 1558
rect 49392 1523 49393 1557
rect 49393 1523 49561 1557
rect 49561 1523 49562 1557
rect 49392 1449 49562 1523
rect 49392 1415 49393 1449
rect 49393 1415 49561 1449
rect 49561 1415 49562 1449
rect 49392 1414 49562 1415
rect 40836 1139 41006 1140
rect 40836 1105 40837 1139
rect 40837 1105 41005 1139
rect 41005 1105 41006 1139
rect 40836 1031 41006 1105
rect 40836 997 40837 1031
rect 40837 997 41005 1031
rect 41005 997 41006 1031
rect 40836 996 41006 997
rect 41208 1139 41378 1140
rect 41208 1105 41209 1139
rect 41209 1105 41377 1139
rect 41377 1105 41378 1139
rect 41208 1031 41378 1105
rect 41208 997 41209 1031
rect 41209 997 41377 1031
rect 41377 997 41378 1031
rect 41208 996 41378 997
rect 41580 1139 41750 1140
rect 41580 1105 41581 1139
rect 41581 1105 41749 1139
rect 41749 1105 41750 1139
rect 41580 1031 41750 1105
rect 41580 997 41581 1031
rect 41581 997 41749 1031
rect 41749 997 41750 1031
rect 41580 996 41750 997
rect 41952 1139 42122 1140
rect 41952 1105 41953 1139
rect 41953 1105 42121 1139
rect 42121 1105 42122 1139
rect 41952 1031 42122 1105
rect 41952 997 41953 1031
rect 41953 997 42121 1031
rect 42121 997 42122 1031
rect 41952 996 42122 997
rect 42324 1139 42494 1140
rect 42324 1105 42325 1139
rect 42325 1105 42493 1139
rect 42493 1105 42494 1139
rect 42324 1031 42494 1105
rect 42324 997 42325 1031
rect 42325 997 42493 1031
rect 42493 997 42494 1031
rect 42324 996 42494 997
rect 42696 1139 42866 1140
rect 42696 1105 42697 1139
rect 42697 1105 42865 1139
rect 42865 1105 42866 1139
rect 42696 1031 42866 1105
rect 42696 997 42697 1031
rect 42697 997 42865 1031
rect 42865 997 42866 1031
rect 42696 996 42866 997
rect 43068 1139 43238 1140
rect 43068 1105 43069 1139
rect 43069 1105 43237 1139
rect 43237 1105 43238 1139
rect 43068 1031 43238 1105
rect 43068 997 43069 1031
rect 43069 997 43237 1031
rect 43237 997 43238 1031
rect 43068 996 43238 997
rect 43440 1139 43610 1140
rect 43440 1105 43441 1139
rect 43441 1105 43609 1139
rect 43609 1105 43610 1139
rect 43440 1031 43610 1105
rect 43440 997 43441 1031
rect 43441 997 43609 1031
rect 43609 997 43610 1031
rect 43440 996 43610 997
rect 43812 1139 43982 1140
rect 43812 1105 43813 1139
rect 43813 1105 43981 1139
rect 43981 1105 43982 1139
rect 43812 1031 43982 1105
rect 43812 997 43813 1031
rect 43813 997 43981 1031
rect 43981 997 43982 1031
rect 43812 996 43982 997
rect 44184 1139 44354 1140
rect 44184 1105 44185 1139
rect 44185 1105 44353 1139
rect 44353 1105 44354 1139
rect 44184 1031 44354 1105
rect 44184 997 44185 1031
rect 44185 997 44353 1031
rect 44353 997 44354 1031
rect 44184 996 44354 997
rect 44556 1139 44726 1140
rect 44556 1105 44557 1139
rect 44557 1105 44725 1139
rect 44725 1105 44726 1139
rect 44556 1031 44726 1105
rect 44556 997 44557 1031
rect 44557 997 44725 1031
rect 44725 997 44726 1031
rect 44556 996 44726 997
rect 44928 1139 45098 1140
rect 44928 1105 44929 1139
rect 44929 1105 45097 1139
rect 45097 1105 45098 1139
rect 44928 1031 45098 1105
rect 44928 997 44929 1031
rect 44929 997 45097 1031
rect 45097 997 45098 1031
rect 44928 996 45098 997
rect 45300 1139 45470 1140
rect 45300 1105 45301 1139
rect 45301 1105 45469 1139
rect 45469 1105 45470 1139
rect 45300 1031 45470 1105
rect 45300 997 45301 1031
rect 45301 997 45469 1031
rect 45469 997 45470 1031
rect 45300 996 45470 997
rect 45672 1139 45842 1140
rect 45672 1105 45673 1139
rect 45673 1105 45841 1139
rect 45841 1105 45842 1139
rect 45672 1031 45842 1105
rect 45672 997 45673 1031
rect 45673 997 45841 1031
rect 45841 997 45842 1031
rect 45672 996 45842 997
rect 46044 1139 46214 1140
rect 46044 1105 46045 1139
rect 46045 1105 46213 1139
rect 46213 1105 46214 1139
rect 46044 1031 46214 1105
rect 46044 997 46045 1031
rect 46045 997 46213 1031
rect 46213 997 46214 1031
rect 46044 996 46214 997
rect 46416 1139 46586 1140
rect 46416 1105 46417 1139
rect 46417 1105 46585 1139
rect 46585 1105 46586 1139
rect 46416 1031 46586 1105
rect 46416 997 46417 1031
rect 46417 997 46585 1031
rect 46585 997 46586 1031
rect 46416 996 46586 997
rect 46788 1139 46958 1140
rect 46788 1105 46789 1139
rect 46789 1105 46957 1139
rect 46957 1105 46958 1139
rect 46788 1031 46958 1105
rect 46788 997 46789 1031
rect 46789 997 46957 1031
rect 46957 997 46958 1031
rect 46788 996 46958 997
rect 47160 1139 47330 1140
rect 47160 1105 47161 1139
rect 47161 1105 47329 1139
rect 47329 1105 47330 1139
rect 47160 1031 47330 1105
rect 47160 997 47161 1031
rect 47161 997 47329 1031
rect 47329 997 47330 1031
rect 47160 996 47330 997
rect 47532 1139 47702 1140
rect 47532 1105 47533 1139
rect 47533 1105 47701 1139
rect 47701 1105 47702 1139
rect 47532 1031 47702 1105
rect 47532 997 47533 1031
rect 47533 997 47701 1031
rect 47701 997 47702 1031
rect 47532 996 47702 997
rect 47904 1139 48074 1140
rect 47904 1105 47905 1139
rect 47905 1105 48073 1139
rect 48073 1105 48074 1139
rect 47904 1031 48074 1105
rect 47904 997 47905 1031
rect 47905 997 48073 1031
rect 48073 997 48074 1031
rect 47904 996 48074 997
rect 48276 1139 48446 1140
rect 48276 1105 48277 1139
rect 48277 1105 48445 1139
rect 48445 1105 48446 1139
rect 48276 1031 48446 1105
rect 48276 997 48277 1031
rect 48277 997 48445 1031
rect 48445 997 48446 1031
rect 48276 996 48446 997
rect 48648 1139 48818 1140
rect 48648 1105 48649 1139
rect 48649 1105 48817 1139
rect 48817 1105 48818 1139
rect 48648 1031 48818 1105
rect 48648 997 48649 1031
rect 48649 997 48817 1031
rect 48817 997 48818 1031
rect 48648 996 48818 997
rect 49020 1139 49190 1140
rect 49020 1105 49021 1139
rect 49021 1105 49189 1139
rect 49189 1105 49190 1139
rect 49020 1031 49190 1105
rect 49020 997 49021 1031
rect 49021 997 49189 1031
rect 49189 997 49190 1031
rect 49020 996 49190 997
rect 49392 1139 49562 1140
rect 49392 1105 49393 1139
rect 49393 1105 49561 1139
rect 49561 1105 49562 1139
rect 49392 1031 49562 1105
rect 49392 997 49393 1031
rect 49393 997 49561 1031
rect 49561 997 49562 1031
rect 49392 996 49562 997
rect 40836 721 41006 722
rect 40836 687 40837 721
rect 40837 687 41005 721
rect 41005 687 41006 721
rect 40836 613 41006 687
rect 40836 579 40837 613
rect 40837 579 41005 613
rect 41005 579 41006 613
rect 40836 578 41006 579
rect 41208 721 41378 722
rect 41208 687 41209 721
rect 41209 687 41377 721
rect 41377 687 41378 721
rect 41208 613 41378 687
rect 41208 579 41209 613
rect 41209 579 41377 613
rect 41377 579 41378 613
rect 41208 578 41378 579
rect 41580 721 41750 722
rect 41580 687 41581 721
rect 41581 687 41749 721
rect 41749 687 41750 721
rect 41580 613 41750 687
rect 41580 579 41581 613
rect 41581 579 41749 613
rect 41749 579 41750 613
rect 41580 578 41750 579
rect 41952 721 42122 722
rect 41952 687 41953 721
rect 41953 687 42121 721
rect 42121 687 42122 721
rect 41952 613 42122 687
rect 41952 579 41953 613
rect 41953 579 42121 613
rect 42121 579 42122 613
rect 41952 578 42122 579
rect 42324 721 42494 722
rect 42324 687 42325 721
rect 42325 687 42493 721
rect 42493 687 42494 721
rect 42324 613 42494 687
rect 42324 579 42325 613
rect 42325 579 42493 613
rect 42493 579 42494 613
rect 42324 578 42494 579
rect 42696 721 42866 722
rect 42696 687 42697 721
rect 42697 687 42865 721
rect 42865 687 42866 721
rect 42696 613 42866 687
rect 42696 579 42697 613
rect 42697 579 42865 613
rect 42865 579 42866 613
rect 42696 578 42866 579
rect 43068 721 43238 722
rect 43068 687 43069 721
rect 43069 687 43237 721
rect 43237 687 43238 721
rect 43068 613 43238 687
rect 43068 579 43069 613
rect 43069 579 43237 613
rect 43237 579 43238 613
rect 43068 578 43238 579
rect 43440 721 43610 722
rect 43440 687 43441 721
rect 43441 687 43609 721
rect 43609 687 43610 721
rect 43440 613 43610 687
rect 43440 579 43441 613
rect 43441 579 43609 613
rect 43609 579 43610 613
rect 43440 578 43610 579
rect 43812 721 43982 722
rect 43812 687 43813 721
rect 43813 687 43981 721
rect 43981 687 43982 721
rect 43812 613 43982 687
rect 43812 579 43813 613
rect 43813 579 43981 613
rect 43981 579 43982 613
rect 43812 578 43982 579
rect 44184 721 44354 722
rect 44184 687 44185 721
rect 44185 687 44353 721
rect 44353 687 44354 721
rect 44184 613 44354 687
rect 44184 579 44185 613
rect 44185 579 44353 613
rect 44353 579 44354 613
rect 44184 578 44354 579
rect 44556 721 44726 722
rect 44556 687 44557 721
rect 44557 687 44725 721
rect 44725 687 44726 721
rect 44556 613 44726 687
rect 44556 579 44557 613
rect 44557 579 44725 613
rect 44725 579 44726 613
rect 44556 578 44726 579
rect 44928 721 45098 722
rect 44928 687 44929 721
rect 44929 687 45097 721
rect 45097 687 45098 721
rect 44928 613 45098 687
rect 44928 579 44929 613
rect 44929 579 45097 613
rect 45097 579 45098 613
rect 44928 578 45098 579
rect 45300 721 45470 722
rect 45300 687 45301 721
rect 45301 687 45469 721
rect 45469 687 45470 721
rect 45300 613 45470 687
rect 45300 579 45301 613
rect 45301 579 45469 613
rect 45469 579 45470 613
rect 45300 578 45470 579
rect 45672 721 45842 722
rect 45672 687 45673 721
rect 45673 687 45841 721
rect 45841 687 45842 721
rect 45672 613 45842 687
rect 45672 579 45673 613
rect 45673 579 45841 613
rect 45841 579 45842 613
rect 45672 578 45842 579
rect 46044 721 46214 722
rect 46044 687 46045 721
rect 46045 687 46213 721
rect 46213 687 46214 721
rect 46044 613 46214 687
rect 46044 579 46045 613
rect 46045 579 46213 613
rect 46213 579 46214 613
rect 46044 578 46214 579
rect 46416 721 46586 722
rect 46416 687 46417 721
rect 46417 687 46585 721
rect 46585 687 46586 721
rect 46416 613 46586 687
rect 46416 579 46417 613
rect 46417 579 46585 613
rect 46585 579 46586 613
rect 46416 578 46586 579
rect 46788 721 46958 722
rect 46788 687 46789 721
rect 46789 687 46957 721
rect 46957 687 46958 721
rect 46788 613 46958 687
rect 46788 579 46789 613
rect 46789 579 46957 613
rect 46957 579 46958 613
rect 46788 578 46958 579
rect 47160 721 47330 722
rect 47160 687 47161 721
rect 47161 687 47329 721
rect 47329 687 47330 721
rect 47160 613 47330 687
rect 47160 579 47161 613
rect 47161 579 47329 613
rect 47329 579 47330 613
rect 47160 578 47330 579
rect 47532 721 47702 722
rect 47532 687 47533 721
rect 47533 687 47701 721
rect 47701 687 47702 721
rect 47532 613 47702 687
rect 47532 579 47533 613
rect 47533 579 47701 613
rect 47701 579 47702 613
rect 47532 578 47702 579
rect 47904 721 48074 722
rect 47904 687 47905 721
rect 47905 687 48073 721
rect 48073 687 48074 721
rect 47904 613 48074 687
rect 47904 579 47905 613
rect 47905 579 48073 613
rect 48073 579 48074 613
rect 47904 578 48074 579
rect 48276 721 48446 722
rect 48276 687 48277 721
rect 48277 687 48445 721
rect 48445 687 48446 721
rect 48276 613 48446 687
rect 48276 579 48277 613
rect 48277 579 48445 613
rect 48445 579 48446 613
rect 48276 578 48446 579
rect 48648 721 48818 722
rect 48648 687 48649 721
rect 48649 687 48817 721
rect 48817 687 48818 721
rect 48648 613 48818 687
rect 48648 579 48649 613
rect 48649 579 48817 613
rect 48817 579 48818 613
rect 48648 578 48818 579
rect 49020 721 49190 722
rect 49020 687 49021 721
rect 49021 687 49189 721
rect 49189 687 49190 721
rect 49020 613 49190 687
rect 49020 579 49021 613
rect 49021 579 49189 613
rect 49189 579 49190 613
rect 49020 578 49190 579
rect 49392 721 49562 722
rect 49392 687 49393 721
rect 49393 687 49561 721
rect 49561 687 49562 721
rect 49392 613 49562 687
rect 49392 579 49393 613
rect 49393 579 49561 613
rect 49561 579 49562 613
rect 49392 578 49562 579
rect 40836 303 41006 314
rect 40836 269 40837 303
rect 40837 269 41005 303
rect 41005 269 41006 303
rect 40836 258 41006 269
rect 41208 303 41378 314
rect 41208 269 41209 303
rect 41209 269 41377 303
rect 41377 269 41378 303
rect 41208 258 41378 269
rect 41580 303 41750 314
rect 41580 269 41581 303
rect 41581 269 41749 303
rect 41749 269 41750 303
rect 41580 258 41750 269
rect 41952 303 42122 314
rect 41952 269 41953 303
rect 41953 269 42121 303
rect 42121 269 42122 303
rect 41952 258 42122 269
rect 42324 303 42494 314
rect 42324 269 42325 303
rect 42325 269 42493 303
rect 42493 269 42494 303
rect 42324 258 42494 269
rect 42696 303 42866 314
rect 42696 269 42697 303
rect 42697 269 42865 303
rect 42865 269 42866 303
rect 42696 258 42866 269
rect 43068 303 43238 314
rect 43068 269 43069 303
rect 43069 269 43237 303
rect 43237 269 43238 303
rect 43068 258 43238 269
rect 43440 303 43610 314
rect 43440 269 43441 303
rect 43441 269 43609 303
rect 43609 269 43610 303
rect 43440 258 43610 269
rect 43812 303 43982 314
rect 43812 269 43813 303
rect 43813 269 43981 303
rect 43981 269 43982 303
rect 43812 258 43982 269
rect 44184 303 44354 314
rect 44184 269 44185 303
rect 44185 269 44353 303
rect 44353 269 44354 303
rect 44184 258 44354 269
rect 44556 303 44726 314
rect 44556 269 44557 303
rect 44557 269 44725 303
rect 44725 269 44726 303
rect 44556 258 44726 269
rect 44928 303 45098 314
rect 44928 269 44929 303
rect 44929 269 45097 303
rect 45097 269 45098 303
rect 44928 258 45098 269
rect 45300 303 45470 314
rect 45300 269 45301 303
rect 45301 269 45469 303
rect 45469 269 45470 303
rect 45300 258 45470 269
rect 45672 303 45842 314
rect 45672 269 45673 303
rect 45673 269 45841 303
rect 45841 269 45842 303
rect 45672 258 45842 269
rect 46044 303 46214 314
rect 46044 269 46045 303
rect 46045 269 46213 303
rect 46213 269 46214 303
rect 46044 258 46214 269
rect 46416 303 46586 314
rect 46416 269 46417 303
rect 46417 269 46585 303
rect 46585 269 46586 303
rect 46416 258 46586 269
rect 46788 303 46958 314
rect 46788 269 46789 303
rect 46789 269 46957 303
rect 46957 269 46958 303
rect 46788 258 46958 269
rect 47160 303 47330 314
rect 47160 269 47161 303
rect 47161 269 47329 303
rect 47329 269 47330 303
rect 47160 258 47330 269
rect 47532 303 47702 314
rect 47532 269 47533 303
rect 47533 269 47701 303
rect 47701 269 47702 303
rect 47532 258 47702 269
rect 47904 303 48074 314
rect 47904 269 47905 303
rect 47905 269 48073 303
rect 48073 269 48074 303
rect 47904 258 48074 269
rect 48276 303 48446 314
rect 48276 269 48277 303
rect 48277 269 48445 303
rect 48445 269 48446 303
rect 48276 258 48446 269
rect 48648 303 48818 314
rect 48648 269 48649 303
rect 48649 269 48817 303
rect 48817 269 48818 303
rect 48648 258 48818 269
rect 49020 303 49190 314
rect 49020 269 49021 303
rect 49021 269 49189 303
rect 49189 269 49190 303
rect 49020 258 49190 269
rect 49392 303 49562 314
rect 49392 269 49393 303
rect 49393 269 49561 303
rect 49561 269 49562 303
rect 49392 258 49562 269
rect 40656 -96 40856 104
rect 41380 -96 41580 104
rect 42124 -96 42324 104
rect 42868 -96 43068 104
rect 43612 -96 43812 104
rect 44356 -96 44556 104
rect 45100 -96 45300 104
rect 45844 -96 46044 104
rect 46588 -96 46788 104
rect 47332 -96 47532 104
rect 48076 -96 48276 104
rect 48820 -96 49020 104
rect 49564 -96 49764 104
<< metal2 >>
rect 40656 19961 40856 19971
rect 40656 19751 40856 19761
rect 41380 19961 41580 19971
rect 41380 19751 41580 19761
rect 42124 19961 42324 19971
rect 42124 19751 42324 19761
rect 42868 19961 43068 19971
rect 42868 19751 43068 19761
rect 43612 19961 43812 19971
rect 43612 19751 43812 19761
rect 44356 19961 44556 19971
rect 44356 19751 44556 19761
rect 45100 19961 45300 19971
rect 45100 19751 45300 19761
rect 45844 19961 46044 19971
rect 45844 19751 46044 19761
rect 46588 19961 46788 19971
rect 46588 19751 46788 19761
rect 47332 19961 47532 19971
rect 47332 19751 47532 19761
rect 48076 19961 48276 19971
rect 48076 19751 48276 19761
rect 48820 19961 49020 19971
rect 48820 19751 49020 19761
rect 49564 19961 49764 19971
rect 49564 19751 49764 19761
rect 40836 19607 43622 19617
rect 41006 19551 41208 19607
rect 41378 19551 41580 19607
rect 41750 19551 41952 19607
rect 42122 19551 42324 19607
rect 42494 19551 42696 19607
rect 42866 19551 43068 19607
rect 43238 19551 43440 19607
rect 43610 19551 43622 19607
rect 40836 19541 43622 19551
rect 43670 19607 49562 19617
rect 43670 19551 43812 19607
rect 43982 19551 44184 19607
rect 44354 19551 44556 19607
rect 44726 19551 44928 19607
rect 45098 19551 45300 19607
rect 45470 19551 45672 19607
rect 45842 19551 46044 19607
rect 46214 19551 46416 19607
rect 46586 19551 46788 19607
rect 46958 19551 47160 19607
rect 47330 19551 47532 19607
rect 47702 19551 47904 19607
rect 48074 19551 48276 19607
rect 48446 19551 48648 19607
rect 48818 19551 49020 19607
rect 49190 19551 49392 19607
rect 43670 19541 49562 19551
rect 43670 19297 43796 19541
rect 40836 19287 43622 19297
rect 41006 19143 41208 19287
rect 41378 19143 41580 19287
rect 41750 19143 41952 19287
rect 42122 19143 42324 19287
rect 42494 19143 42696 19287
rect 42866 19143 43068 19287
rect 43238 19143 43440 19287
rect 43610 19143 43622 19287
rect 40836 19133 43622 19143
rect 43670 19287 49562 19297
rect 43670 19143 43812 19287
rect 43982 19143 44184 19287
rect 44354 19143 44556 19287
rect 44726 19143 44928 19287
rect 45098 19143 45300 19287
rect 45470 19143 45672 19287
rect 45842 19143 46044 19287
rect 46214 19143 46416 19287
rect 46586 19143 46788 19287
rect 46958 19143 47160 19287
rect 47330 19143 47532 19287
rect 47702 19143 47904 19287
rect 48074 19143 48276 19287
rect 48446 19143 48648 19287
rect 48818 19143 49020 19287
rect 49190 19143 49392 19287
rect 43670 19133 49562 19143
rect 43670 18879 43796 19133
rect 40836 18869 43622 18879
rect 41006 18725 41208 18869
rect 41378 18725 41580 18869
rect 41750 18725 41952 18869
rect 42122 18725 42324 18869
rect 42494 18725 42696 18869
rect 42866 18725 43068 18869
rect 43238 18725 43440 18869
rect 43610 18725 43622 18869
rect 40836 18715 43622 18725
rect 43670 18869 49562 18879
rect 43670 18725 43812 18869
rect 43982 18725 44184 18869
rect 44354 18725 44556 18869
rect 44726 18725 44928 18869
rect 45098 18725 45300 18869
rect 45470 18725 45672 18869
rect 45842 18725 46044 18869
rect 46214 18725 46416 18869
rect 46586 18725 46788 18869
rect 46958 18725 47160 18869
rect 47330 18725 47532 18869
rect 47702 18725 47904 18869
rect 48074 18725 48276 18869
rect 48446 18725 48648 18869
rect 48818 18725 49020 18869
rect 49190 18725 49392 18869
rect 43670 18715 49562 18725
rect 43670 18461 43796 18715
rect 40836 18451 43622 18461
rect 41006 18307 41208 18451
rect 41378 18307 41580 18451
rect 41750 18307 41952 18451
rect 42122 18307 42324 18451
rect 42494 18307 42696 18451
rect 42866 18307 43068 18451
rect 43238 18307 43440 18451
rect 43610 18307 43622 18451
rect 40836 18297 43622 18307
rect 43670 18451 49562 18461
rect 43670 18307 43812 18451
rect 43982 18307 44184 18451
rect 44354 18307 44556 18451
rect 44726 18307 44928 18451
rect 45098 18307 45300 18451
rect 45470 18307 45672 18451
rect 45842 18307 46044 18451
rect 46214 18307 46416 18451
rect 46586 18307 46788 18451
rect 46958 18307 47160 18451
rect 47330 18307 47532 18451
rect 47702 18307 47904 18451
rect 48074 18307 48276 18451
rect 48446 18307 48648 18451
rect 48818 18307 49020 18451
rect 49190 18307 49392 18451
rect 43670 18297 49562 18307
rect 43670 18053 43796 18297
rect 40836 18043 43622 18053
rect 41006 17987 41208 18043
rect 41378 17987 41580 18043
rect 41750 17987 41952 18043
rect 42122 17987 42324 18043
rect 42494 17987 42696 18043
rect 42866 17987 43068 18043
rect 43238 17987 43440 18043
rect 43610 17987 43622 18043
rect 40836 17977 43622 17987
rect 43670 18043 49562 18053
rect 43670 17987 43812 18043
rect 43982 17987 44184 18043
rect 44354 17987 44556 18043
rect 44726 17987 44928 18043
rect 45098 17987 45300 18043
rect 45470 17987 45672 18043
rect 45842 17987 46044 18043
rect 46214 17987 46416 18043
rect 46586 17987 46788 18043
rect 46958 17987 47160 18043
rect 47330 17987 47532 18043
rect 47702 17987 47904 18043
rect 48074 17987 48276 18043
rect 48446 17987 48648 18043
rect 48818 17987 49020 18043
rect 49190 17987 49392 18043
rect 43670 17977 49562 17987
rect 43670 17859 43796 17977
rect 41816 17849 43796 17859
rect 42630 17803 43796 17849
rect 45826 17815 46104 17825
rect 42630 17669 45826 17803
rect 41816 17659 45826 17669
rect 38314 17616 38800 17626
rect 38800 17591 40714 17592
rect 38800 17493 42680 17591
rect 46104 17659 46118 17803
rect 38800 17492 40714 17493
rect 41766 17393 41936 17493
rect 42510 17393 42680 17493
rect 43942 17525 44224 17535
rect 40836 17383 41378 17393
rect 41006 17329 41208 17383
rect 40836 17319 41378 17329
rect 41580 17383 42866 17393
rect 41750 17329 41952 17383
rect 42122 17329 42324 17383
rect 42494 17329 42696 17383
rect 41580 17319 42866 17329
rect 43068 17383 43610 17393
rect 43238 17329 43440 17383
rect 43068 17319 43610 17329
rect 38314 17098 38800 17108
rect 41080 16457 41134 17319
rect 41824 16457 41878 17319
rect 42568 16457 42622 17319
rect 43312 16457 43366 17319
rect 44686 17525 44968 17535
rect 44224 17253 44686 17417
rect 45430 17525 45712 17535
rect 45826 17531 46104 17541
rect 44968 17253 45430 17417
rect 46174 17525 46456 17535
rect 45712 17253 46174 17417
rect 46918 17525 47200 17535
rect 46456 17253 46918 17417
rect 47662 17525 47944 17535
rect 47200 17253 47662 17417
rect 48406 17525 48688 17535
rect 47944 17253 48406 17417
rect 49150 17525 49432 17535
rect 48688 17253 49150 17417
rect 49432 17253 49442 17417
rect 43942 17243 49442 17253
rect 45566 16470 45734 16480
rect 40836 16447 41378 16457
rect 41006 16303 41208 16447
rect 40836 16293 41378 16303
rect 41580 16447 42866 16457
rect 41750 16303 41952 16447
rect 42122 16303 42324 16447
rect 42494 16303 42696 16447
rect 41580 16293 42866 16303
rect 43068 16447 43610 16457
rect 43238 16303 43440 16447
rect 43068 16293 43610 16303
rect 45566 16294 45734 16304
rect 41080 15421 41134 16293
rect 41824 15421 41878 16293
rect 42568 15421 42622 16293
rect 43312 15421 43366 16293
rect 45566 16070 45734 16080
rect 45566 15894 45734 15904
rect 45566 15670 45734 15680
rect 45566 15494 45734 15504
rect 40836 15411 41378 15421
rect 41006 15267 41208 15411
rect 40836 15257 41378 15267
rect 41580 15411 42866 15421
rect 41750 15267 41952 15411
rect 42122 15267 42324 15411
rect 42494 15267 42696 15411
rect 41580 15257 42866 15267
rect 43068 15411 43610 15421
rect 43238 15267 43440 15411
rect 43068 15257 43610 15267
rect 41080 14385 41134 15257
rect 41824 14385 41878 15257
rect 42568 14385 42622 15257
rect 43312 14385 43366 15257
rect 45852 15117 46134 15127
rect 45852 14835 46134 14845
rect 45964 14453 46448 14463
rect 40836 14375 41378 14385
rect 41006 14231 41208 14375
rect 40836 14221 41378 14231
rect 41580 14375 42866 14385
rect 41750 14231 41952 14375
rect 42122 14231 42324 14375
rect 42494 14231 42696 14375
rect 41580 14221 42866 14231
rect 43068 14375 43610 14385
rect 43238 14231 43440 14375
rect 43068 14221 43610 14231
rect 41080 13363 41134 14221
rect 41824 13363 41878 14221
rect 42568 13363 42622 14221
rect 43312 13363 43366 14221
rect 44422 14095 45964 14307
rect 40836 13353 41378 13363
rect 41006 13289 41208 13353
rect 40836 13279 41378 13289
rect 41580 13353 42866 13363
rect 41750 13289 41952 13353
rect 42122 13289 42324 13353
rect 42494 13289 42696 13353
rect 41580 13279 42866 13289
rect 43068 13353 43610 13363
rect 43238 13289 43440 13353
rect 43068 13279 43610 13289
rect 41022 13189 41192 13279
rect 43254 13219 43424 13279
rect 44422 13219 44602 14095
rect 45964 13943 46448 13953
rect 43254 13189 44602 13219
rect 40356 13091 44602 13189
rect 45432 13343 50922 13353
rect 45714 13071 46176 13343
rect 46458 13071 46920 13343
rect 47202 13071 47664 13343
rect 47946 13071 48408 13343
rect 48690 13071 49152 13343
rect 49434 13071 49896 13343
rect 50178 13071 50640 13343
rect 45432 13061 50922 13071
rect 39348 12763 51050 12773
rect 39518 12703 39720 12763
rect 39890 12703 40092 12763
rect 40262 12703 40464 12763
rect 40634 12703 40836 12763
rect 41006 12703 41208 12763
rect 41378 12703 41580 12763
rect 41750 12703 41952 12763
rect 42122 12703 42324 12763
rect 42494 12703 42696 12763
rect 42866 12703 43068 12763
rect 43238 12703 43440 12763
rect 43610 12703 43812 12763
rect 43982 12703 44184 12763
rect 44354 12703 44556 12763
rect 44726 12703 44928 12763
rect 45098 12703 45300 12763
rect 45470 12703 45672 12763
rect 45842 12703 46044 12763
rect 46214 12703 46416 12763
rect 46586 12703 46788 12763
rect 46958 12703 47160 12763
rect 47330 12703 47532 12763
rect 47702 12703 47904 12763
rect 48074 12703 48276 12763
rect 48446 12703 48648 12763
rect 48818 12703 49020 12763
rect 49190 12703 49392 12763
rect 49562 12703 49764 12763
rect 49934 12703 50136 12763
rect 50306 12703 50508 12763
rect 50678 12703 50880 12763
rect 39348 12693 51050 12703
rect 39348 12223 51050 12233
rect 39518 12079 39720 12223
rect 39890 12079 40092 12223
rect 40262 12079 40464 12223
rect 40634 12079 40836 12223
rect 41006 12079 41208 12223
rect 41378 12079 41580 12223
rect 41750 12079 41952 12223
rect 42122 12079 42324 12223
rect 42494 12079 42696 12223
rect 42866 12079 43068 12223
rect 43238 12079 43440 12223
rect 43610 12079 43812 12223
rect 43982 12079 44184 12223
rect 44354 12079 44556 12223
rect 44726 12079 44928 12223
rect 45098 12079 45300 12223
rect 45470 12079 45672 12223
rect 45842 12079 46044 12223
rect 46214 12079 46416 12223
rect 46586 12079 46788 12223
rect 46958 12079 47160 12223
rect 47330 12079 47532 12223
rect 47702 12079 47904 12223
rect 48074 12079 48276 12223
rect 48446 12079 48648 12223
rect 48818 12079 49020 12223
rect 49190 12079 49392 12223
rect 49562 12079 49764 12223
rect 49934 12079 50136 12223
rect 50306 12079 50508 12223
rect 50678 12079 50880 12223
rect 39348 12069 51050 12079
rect 39348 11587 51050 11597
rect 39518 11443 39720 11587
rect 39890 11443 40092 11587
rect 40262 11443 40464 11587
rect 40634 11443 40836 11587
rect 41006 11443 41208 11587
rect 41378 11443 41580 11587
rect 41750 11443 41952 11587
rect 42122 11443 42324 11587
rect 42494 11443 42696 11587
rect 42866 11443 43068 11587
rect 43238 11443 43440 11587
rect 43610 11443 43812 11587
rect 43982 11443 44184 11587
rect 44354 11443 44556 11587
rect 44726 11443 44928 11587
rect 45098 11443 45300 11587
rect 45470 11443 45672 11587
rect 45842 11443 46044 11587
rect 46214 11443 46416 11587
rect 46586 11443 46788 11587
rect 46958 11443 47160 11587
rect 47330 11443 47532 11587
rect 47702 11443 47904 11587
rect 48074 11443 48276 11587
rect 48446 11443 48648 11587
rect 48818 11443 49020 11587
rect 49190 11443 49392 11587
rect 49562 11443 49764 11587
rect 49934 11443 50136 11587
rect 50306 11443 50508 11587
rect 50678 11443 50880 11587
rect 39348 11433 51050 11443
rect 39348 10963 51060 10973
rect 39518 10903 39720 10963
rect 39890 10903 40092 10963
rect 40262 10903 40464 10963
rect 40634 10903 40836 10963
rect 41006 10903 41208 10963
rect 41378 10903 41580 10963
rect 41750 10903 41952 10963
rect 42122 10903 42324 10963
rect 42494 10903 42696 10963
rect 42866 10903 43068 10963
rect 43238 10903 43440 10963
rect 43610 10903 43812 10963
rect 43982 10903 44184 10963
rect 44354 10903 44556 10963
rect 44726 10903 44928 10963
rect 45098 10903 45300 10963
rect 45470 10903 45672 10963
rect 45842 10903 46044 10963
rect 46214 10903 46416 10963
rect 46586 10903 46788 10963
rect 46958 10903 47160 10963
rect 47330 10903 47532 10963
rect 47702 10903 47904 10963
rect 48074 10903 48276 10963
rect 48446 10903 48648 10963
rect 48818 10903 49020 10963
rect 49190 10903 49392 10963
rect 49562 10903 49764 10963
rect 49934 10903 50136 10963
rect 50306 10903 50508 10963
rect 50678 10903 50880 10963
rect 51050 10903 51060 10963
rect 39348 10893 51060 10903
rect 39518 10715 39718 10725
rect 39518 10505 39718 10515
rect 40262 10715 40462 10725
rect 40262 10505 40462 10515
rect 41006 10715 41206 10725
rect 41006 10505 41206 10515
rect 41750 10715 41950 10725
rect 41750 10505 41950 10515
rect 42494 10715 42694 10725
rect 42494 10505 42694 10515
rect 43238 10715 43438 10725
rect 43238 10505 43438 10515
rect 43982 10715 44182 10725
rect 43982 10505 44182 10515
rect 44726 10715 44926 10725
rect 44726 10505 44926 10515
rect 45098 10715 45298 10725
rect 45098 10505 45298 10515
rect 45842 10715 46042 10725
rect 45842 10505 46042 10515
rect 46586 10715 46786 10725
rect 46586 10505 46786 10515
rect 47330 10715 47530 10725
rect 47330 10505 47530 10515
rect 48074 10715 48274 10725
rect 48074 10505 48274 10515
rect 48818 10715 49018 10725
rect 48818 10505 49018 10515
rect 49562 10715 49762 10725
rect 49562 10505 49762 10515
rect 50306 10715 50506 10725
rect 50306 10505 50506 10515
rect 51050 10715 51250 10725
rect 51050 10505 51250 10515
rect 39518 9350 39718 9360
rect 39518 9140 39718 9150
rect 40262 9350 40462 9360
rect 40262 9140 40462 9150
rect 41006 9350 41206 9360
rect 41006 9140 41206 9150
rect 41750 9350 41950 9360
rect 41750 9140 41950 9150
rect 42494 9350 42694 9360
rect 42494 9140 42694 9150
rect 43238 9350 43438 9360
rect 43238 9140 43438 9150
rect 43982 9350 44182 9360
rect 43982 9140 44182 9150
rect 44726 9350 44926 9360
rect 44726 9140 44926 9150
rect 45098 9350 45298 9360
rect 45098 9140 45298 9150
rect 45842 9350 46042 9360
rect 45842 9140 46042 9150
rect 46586 9350 46786 9360
rect 46586 9140 46786 9150
rect 47330 9350 47530 9360
rect 47330 9140 47530 9150
rect 48074 9350 48274 9360
rect 48074 9140 48274 9150
rect 48818 9350 49018 9360
rect 48818 9140 49018 9150
rect 49562 9350 49762 9360
rect 49562 9140 49762 9150
rect 50306 9350 50506 9360
rect 50306 9140 50506 9150
rect 51050 9350 51250 9360
rect 51050 9140 51250 9150
rect 39348 8962 51060 8972
rect 39518 8902 39720 8962
rect 39890 8902 40092 8962
rect 40262 8902 40464 8962
rect 40634 8902 40836 8962
rect 41006 8902 41208 8962
rect 41378 8902 41580 8962
rect 41750 8902 41952 8962
rect 42122 8902 42324 8962
rect 42494 8902 42696 8962
rect 42866 8902 43068 8962
rect 43238 8902 43440 8962
rect 43610 8902 43812 8962
rect 43982 8902 44184 8962
rect 44354 8902 44556 8962
rect 44726 8902 44928 8962
rect 45098 8902 45300 8962
rect 45470 8902 45672 8962
rect 45842 8902 46044 8962
rect 46214 8902 46416 8962
rect 46586 8902 46788 8962
rect 46958 8902 47160 8962
rect 47330 8902 47532 8962
rect 47702 8902 47904 8962
rect 48074 8902 48276 8962
rect 48446 8902 48648 8962
rect 48818 8902 49020 8962
rect 49190 8902 49392 8962
rect 49562 8902 49764 8962
rect 49934 8902 50136 8962
rect 50306 8902 50508 8962
rect 50678 8902 50880 8962
rect 51050 8902 51060 8962
rect 39348 8892 51060 8902
rect 39348 8422 51050 8432
rect 39518 8278 39720 8422
rect 39890 8278 40092 8422
rect 40262 8278 40464 8422
rect 40634 8278 40836 8422
rect 41006 8278 41208 8422
rect 41378 8278 41580 8422
rect 41750 8278 41952 8422
rect 42122 8278 42324 8422
rect 42494 8278 42696 8422
rect 42866 8278 43068 8422
rect 43238 8278 43440 8422
rect 43610 8278 43812 8422
rect 43982 8278 44184 8422
rect 44354 8278 44556 8422
rect 44726 8278 44928 8422
rect 45098 8278 45300 8422
rect 45470 8278 45672 8422
rect 45842 8278 46044 8422
rect 46214 8278 46416 8422
rect 46586 8278 46788 8422
rect 46958 8278 47160 8422
rect 47330 8278 47532 8422
rect 47702 8278 47904 8422
rect 48074 8278 48276 8422
rect 48446 8278 48648 8422
rect 48818 8278 49020 8422
rect 49190 8278 49392 8422
rect 49562 8278 49764 8422
rect 49934 8278 50136 8422
rect 50306 8278 50508 8422
rect 50678 8278 50880 8422
rect 39348 8268 51050 8278
rect 39348 7786 51050 7796
rect 39518 7642 39720 7786
rect 39890 7642 40092 7786
rect 40262 7642 40464 7786
rect 40634 7642 40836 7786
rect 41006 7642 41208 7786
rect 41378 7642 41580 7786
rect 41750 7642 41952 7786
rect 42122 7642 42324 7786
rect 42494 7642 42696 7786
rect 42866 7642 43068 7786
rect 43238 7642 43440 7786
rect 43610 7642 43812 7786
rect 43982 7642 44184 7786
rect 44354 7642 44556 7786
rect 44726 7642 44928 7786
rect 45098 7642 45300 7786
rect 45470 7642 45672 7786
rect 45842 7642 46044 7786
rect 46214 7642 46416 7786
rect 46586 7642 46788 7786
rect 46958 7642 47160 7786
rect 47330 7642 47532 7786
rect 47702 7642 47904 7786
rect 48074 7642 48276 7786
rect 48446 7642 48648 7786
rect 48818 7642 49020 7786
rect 49190 7642 49392 7786
rect 49562 7642 49764 7786
rect 49934 7642 50136 7786
rect 50306 7642 50508 7786
rect 50678 7642 50880 7786
rect 39348 7632 51050 7642
rect 39348 7162 51050 7172
rect 39518 7102 39720 7162
rect 39890 7102 40092 7162
rect 40262 7102 40464 7162
rect 40634 7102 40836 7162
rect 41006 7102 41208 7162
rect 41378 7102 41580 7162
rect 41750 7102 41952 7162
rect 42122 7102 42324 7162
rect 42494 7102 42696 7162
rect 42866 7102 43068 7162
rect 43238 7102 43440 7162
rect 43610 7102 43812 7162
rect 43982 7102 44184 7162
rect 44354 7102 44556 7162
rect 44726 7102 44928 7162
rect 45098 7102 45300 7162
rect 45470 7102 45672 7162
rect 45842 7102 46044 7162
rect 46214 7102 46416 7162
rect 46586 7102 46788 7162
rect 46958 7102 47160 7162
rect 47330 7102 47532 7162
rect 47702 7102 47904 7162
rect 48074 7102 48276 7162
rect 48446 7102 48648 7162
rect 48818 7102 49020 7162
rect 49190 7102 49392 7162
rect 49562 7102 49764 7162
rect 49934 7102 50136 7162
rect 50306 7102 50508 7162
rect 50678 7102 50880 7162
rect 39348 7092 51050 7102
rect 44616 6831 44898 6841
rect 40122 6774 40404 6775
rect 40122 6773 43424 6774
rect 40122 6676 44616 6773
rect 40122 6675 40404 6676
rect 41022 6586 41192 6676
rect 43254 6639 44616 6676
rect 43254 6586 43424 6639
rect 40836 6576 41378 6586
rect 41006 6512 41208 6576
rect 40836 6502 41378 6512
rect 41580 6576 42866 6586
rect 41750 6512 41952 6576
rect 42122 6512 42324 6576
rect 42494 6512 42696 6576
rect 41580 6502 42866 6512
rect 43068 6576 43610 6586
rect 43238 6512 43440 6576
rect 44616 6547 44898 6557
rect 45432 6794 50922 6804
rect 45714 6522 46176 6794
rect 46458 6522 46920 6794
rect 47202 6522 47664 6794
rect 47946 6522 48408 6794
rect 48690 6522 49152 6794
rect 49434 6522 49896 6794
rect 50178 6522 50640 6794
rect 45432 6512 50922 6522
rect 43068 6502 43610 6512
rect 40122 6391 40404 6401
rect 40246 6259 40392 6269
rect 40246 6099 40392 6109
rect 40246 5859 40392 5869
rect 40246 5699 40392 5709
rect 41080 5644 41134 6502
rect 41824 5644 41878 6502
rect 42568 5644 42622 6502
rect 43312 5644 43366 6502
rect 45638 6135 46122 6145
rect 44162 5719 44308 5729
rect 40836 5634 41378 5644
rect 41006 5490 41208 5634
rect 40836 5480 41378 5490
rect 41580 5634 42866 5644
rect 41750 5490 41952 5634
rect 42122 5490 42324 5634
rect 42494 5490 42696 5634
rect 41580 5480 42866 5490
rect 43068 5634 43610 5644
rect 43238 5490 43440 5634
rect 45638 5625 46122 5635
rect 44162 5559 44308 5569
rect 43068 5480 43610 5490
rect 40246 5459 40392 5469
rect 40246 5299 40392 5309
rect 40246 5059 40392 5069
rect 40246 4899 40392 4909
rect 41080 4608 41134 5480
rect 41824 4608 41878 5480
rect 42568 4608 42622 5480
rect 43312 4608 43366 5480
rect 44162 5319 44308 5329
rect 44162 5159 44308 5169
rect 45852 5020 46134 5030
rect 44162 4919 44308 4929
rect 44162 4759 44308 4769
rect 45852 4738 46134 4748
rect 40836 4598 41378 4608
rect 41006 4454 41208 4598
rect 40836 4444 41378 4454
rect 41580 4598 42866 4608
rect 41750 4454 41952 4598
rect 42122 4454 42324 4598
rect 42494 4454 42696 4598
rect 41580 4444 42866 4454
rect 43068 4598 43610 4608
rect 43238 4454 43440 4598
rect 43068 4444 43610 4454
rect 44162 4519 44308 4529
rect 41080 3572 41134 4444
rect 41824 3572 41878 4444
rect 42568 3572 42622 4444
rect 43312 3572 43366 4444
rect 44162 4359 44308 4369
rect 45556 4306 45730 4316
rect 45556 4122 45730 4132
rect 45556 3906 45730 3916
rect 45556 3722 45730 3732
rect 40836 3562 41378 3572
rect 41006 3418 41208 3562
rect 40836 3408 41378 3418
rect 41580 3562 42866 3572
rect 41750 3418 41952 3562
rect 42122 3418 42324 3562
rect 42494 3418 42696 3562
rect 41580 3408 42866 3418
rect 43068 3562 43610 3572
rect 43238 3418 43440 3562
rect 43068 3408 43610 3418
rect 45556 3506 45730 3516
rect 41080 2546 41134 3408
rect 41824 2546 41878 3408
rect 42568 2546 42622 3408
rect 43312 2546 43366 3408
rect 45556 3322 45730 3332
rect 43942 2612 49442 2622
rect 40836 2536 41378 2546
rect 41006 2482 41208 2536
rect 40836 2472 41378 2482
rect 41580 2536 42866 2546
rect 41750 2482 41952 2536
rect 42122 2482 42324 2536
rect 42494 2482 42696 2536
rect 41580 2472 42866 2482
rect 43068 2536 43610 2546
rect 43238 2482 43440 2536
rect 43068 2472 43610 2482
rect 41766 2372 41936 2472
rect 42510 2372 42680 2472
rect 40356 2274 42680 2372
rect 44224 2448 44686 2612
rect 43942 2330 44224 2340
rect 44968 2448 45430 2612
rect 44686 2330 44968 2340
rect 45712 2448 46174 2612
rect 45430 2330 45712 2340
rect 46456 2448 46918 2612
rect 45826 2324 46104 2334
rect 46174 2330 46456 2340
rect 47200 2448 47662 2612
rect 46918 2330 47200 2340
rect 47944 2448 48406 2612
rect 47662 2330 47944 2340
rect 48688 2448 49150 2612
rect 48406 2330 48688 2340
rect 49432 2448 49442 2612
rect 49150 2330 49432 2340
rect 41816 2196 45826 2206
rect 42630 2062 45826 2196
rect 42630 2016 43796 2062
rect 46104 2062 46118 2206
rect 45826 2040 46104 2050
rect 41816 2006 43796 2016
rect 43670 1888 43796 2006
rect 40836 1878 43622 1888
rect 41006 1822 41208 1878
rect 41378 1822 41580 1878
rect 41750 1822 41952 1878
rect 42122 1822 42324 1878
rect 42494 1822 42696 1878
rect 42866 1822 43068 1878
rect 43238 1822 43440 1878
rect 43610 1822 43622 1878
rect 40836 1812 43622 1822
rect 43670 1878 49562 1888
rect 43670 1822 43812 1878
rect 43982 1822 44184 1878
rect 44354 1822 44556 1878
rect 44726 1822 44928 1878
rect 45098 1822 45300 1878
rect 45470 1822 45672 1878
rect 45842 1822 46044 1878
rect 46214 1822 46416 1878
rect 46586 1822 46788 1878
rect 46958 1822 47160 1878
rect 47330 1822 47532 1878
rect 47702 1822 47904 1878
rect 48074 1822 48276 1878
rect 48446 1822 48648 1878
rect 48818 1822 49020 1878
rect 49190 1822 49392 1878
rect 43670 1812 49562 1822
rect 43670 1568 43796 1812
rect 40836 1558 43622 1568
rect 41006 1414 41208 1558
rect 41378 1414 41580 1558
rect 41750 1414 41952 1558
rect 42122 1414 42324 1558
rect 42494 1414 42696 1558
rect 42866 1414 43068 1558
rect 43238 1414 43440 1558
rect 43610 1414 43622 1558
rect 40836 1404 43622 1414
rect 43670 1558 49562 1568
rect 43670 1414 43812 1558
rect 43982 1414 44184 1558
rect 44354 1414 44556 1558
rect 44726 1414 44928 1558
rect 45098 1414 45300 1558
rect 45470 1414 45672 1558
rect 45842 1414 46044 1558
rect 46214 1414 46416 1558
rect 46586 1414 46788 1558
rect 46958 1414 47160 1558
rect 47330 1414 47532 1558
rect 47702 1414 47904 1558
rect 48074 1414 48276 1558
rect 48446 1414 48648 1558
rect 48818 1414 49020 1558
rect 49190 1414 49392 1558
rect 43670 1404 49562 1414
rect 43670 1150 43796 1404
rect 40836 1140 43622 1150
rect 41006 996 41208 1140
rect 41378 996 41580 1140
rect 41750 996 41952 1140
rect 42122 996 42324 1140
rect 42494 996 42696 1140
rect 42866 996 43068 1140
rect 43238 996 43440 1140
rect 43610 996 43622 1140
rect 40836 986 43622 996
rect 43670 1140 49562 1150
rect 43670 996 43812 1140
rect 43982 996 44184 1140
rect 44354 996 44556 1140
rect 44726 996 44928 1140
rect 45098 996 45300 1140
rect 45470 996 45672 1140
rect 45842 996 46044 1140
rect 46214 996 46416 1140
rect 46586 996 46788 1140
rect 46958 996 47160 1140
rect 47330 996 47532 1140
rect 47702 996 47904 1140
rect 48074 996 48276 1140
rect 48446 996 48648 1140
rect 48818 996 49020 1140
rect 49190 996 49392 1140
rect 43670 986 49562 996
rect 43670 732 43796 986
rect 40836 722 43622 732
rect 41006 578 41208 722
rect 41378 578 41580 722
rect 41750 578 41952 722
rect 42122 578 42324 722
rect 42494 578 42696 722
rect 42866 578 43068 722
rect 43238 578 43440 722
rect 43610 578 43622 722
rect 40836 568 43622 578
rect 43670 722 49562 732
rect 43670 578 43812 722
rect 43982 578 44184 722
rect 44354 578 44556 722
rect 44726 578 44928 722
rect 45098 578 45300 722
rect 45470 578 45672 722
rect 45842 578 46044 722
rect 46214 578 46416 722
rect 46586 578 46788 722
rect 46958 578 47160 722
rect 47330 578 47532 722
rect 47702 578 47904 722
rect 48074 578 48276 722
rect 48446 578 48648 722
rect 48818 578 49020 722
rect 49190 578 49392 722
rect 43670 568 49562 578
rect 43670 324 43796 568
rect 40836 314 43622 324
rect 41006 258 41208 314
rect 41378 258 41580 314
rect 41750 258 41952 314
rect 42122 258 42324 314
rect 42494 258 42696 314
rect 42866 258 43068 314
rect 43238 258 43440 314
rect 43610 258 43622 314
rect 40836 248 43622 258
rect 43670 314 49562 324
rect 43670 258 43812 314
rect 43982 258 44184 314
rect 44354 258 44556 314
rect 44726 258 44928 314
rect 45098 258 45300 314
rect 45470 258 45672 314
rect 45842 258 46044 314
rect 46214 258 46416 314
rect 46586 258 46788 314
rect 46958 258 47160 314
rect 47330 258 47532 314
rect 47702 258 47904 314
rect 48074 258 48276 314
rect 48446 258 48648 314
rect 48818 258 49020 314
rect 49190 258 49392 314
rect 43670 248 49562 258
rect 40656 104 40856 114
rect 40656 -106 40856 -96
rect 41380 104 41580 114
rect 41380 -106 41580 -96
rect 42124 104 42324 114
rect 42124 -106 42324 -96
rect 42868 104 43068 114
rect 42868 -106 43068 -96
rect 43612 104 43812 114
rect 43612 -106 43812 -96
rect 44356 104 44556 114
rect 44356 -106 44556 -96
rect 45100 104 45300 114
rect 45100 -106 45300 -96
rect 45844 104 46044 114
rect 45844 -106 46044 -96
rect 46588 104 46788 114
rect 46588 -106 46788 -96
rect 47332 104 47532 114
rect 47332 -106 47532 -96
rect 48076 104 48276 114
rect 48076 -106 48276 -96
rect 48820 104 49020 114
rect 48820 -106 49020 -96
rect 49564 104 49764 114
rect 49564 -106 49764 -96
<< via2 >>
rect 40656 19761 40856 19961
rect 41380 19761 41580 19961
rect 42124 19761 42324 19961
rect 42868 19761 43068 19961
rect 43612 19761 43812 19961
rect 44356 19761 44556 19961
rect 45100 19761 45300 19961
rect 45844 19761 46044 19961
rect 46588 19761 46788 19961
rect 47332 19761 47532 19961
rect 48076 19761 48276 19961
rect 48820 19761 49020 19961
rect 49564 19761 49764 19961
rect 46918 17253 47200 17525
rect 47662 17253 47944 17525
rect 48406 17253 48688 17525
rect 49150 17253 49432 17525
rect 45566 16304 45734 16470
rect 45566 15904 45734 16070
rect 45566 15504 45734 15670
rect 45852 14845 46134 15117
rect 45964 13953 46448 14453
rect 46920 13071 47202 13343
rect 47664 13071 47946 13343
rect 48408 13071 48690 13343
rect 49152 13071 49434 13343
rect 39518 10515 39718 10715
rect 40262 10515 40462 10715
rect 41006 10515 41206 10715
rect 41750 10515 41950 10715
rect 42494 10515 42694 10715
rect 43238 10515 43438 10715
rect 43982 10515 44182 10715
rect 44726 10515 44926 10715
rect 45098 10515 45298 10715
rect 45842 10515 46042 10715
rect 46586 10515 46786 10715
rect 47330 10515 47530 10715
rect 48074 10515 48274 10715
rect 48818 10515 49018 10715
rect 49562 10515 49762 10715
rect 50306 10515 50506 10715
rect 51050 10515 51250 10715
rect 39518 9150 39718 9350
rect 40262 9150 40462 9350
rect 41006 9150 41206 9350
rect 41750 9150 41950 9350
rect 42494 9150 42694 9350
rect 43238 9150 43438 9350
rect 43982 9150 44182 9350
rect 44726 9150 44926 9350
rect 45098 9150 45298 9350
rect 45842 9150 46042 9350
rect 46586 9150 46786 9350
rect 47330 9150 47530 9350
rect 48074 9150 48274 9350
rect 48818 9150 49018 9350
rect 49562 9150 49762 9350
rect 50306 9150 50506 9350
rect 51050 9150 51250 9350
rect 46920 6522 47202 6794
rect 47664 6522 47946 6794
rect 48408 6522 48690 6794
rect 49152 6522 49434 6794
rect 40246 6109 40392 6259
rect 40246 5709 40392 5859
rect 44162 5569 44308 5719
rect 45638 5635 46122 6135
rect 40246 5309 40392 5459
rect 40246 4909 40392 5059
rect 44162 5169 44308 5319
rect 44162 4769 44308 4919
rect 45852 4748 46134 5020
rect 44162 4369 44308 4519
rect 45556 4132 45730 4306
rect 45556 3732 45730 3906
rect 45556 3332 45730 3506
rect 46918 2340 47200 2612
rect 47662 2340 47944 2612
rect 48406 2340 48688 2612
rect 49150 2340 49432 2612
rect 40656 -96 40856 104
rect 41380 -96 41580 104
rect 42124 -96 42324 104
rect 42868 -96 43068 104
rect 43612 -96 43812 104
rect 44356 -96 44556 104
rect 45100 -96 45300 104
rect 45844 -96 46044 104
rect 46588 -96 46788 104
rect 47332 -96 47532 104
rect 48076 -96 48276 104
rect 48820 -96 49020 104
rect 49564 -96 49764 104
<< metal3 >>
rect 40646 19961 40866 19966
rect 40646 19761 40656 19961
rect 40856 19761 40866 19961
rect 40646 19756 40866 19761
rect 41370 19961 41590 19966
rect 41370 19761 41380 19961
rect 41580 19761 41590 19961
rect 41370 19756 41590 19761
rect 42114 19961 42334 19966
rect 42114 19761 42124 19961
rect 42324 19761 42334 19961
rect 42114 19756 42334 19761
rect 42858 19961 43078 19966
rect 42858 19761 42868 19961
rect 43068 19761 43078 19961
rect 42858 19756 43078 19761
rect 43602 19961 43822 19966
rect 43602 19761 43612 19961
rect 43812 19761 43822 19961
rect 43602 19756 43822 19761
rect 44346 19961 44566 19966
rect 44346 19761 44356 19961
rect 44556 19761 44566 19961
rect 44346 19756 44566 19761
rect 45090 19961 45310 19966
rect 45090 19761 45100 19961
rect 45300 19761 45310 19961
rect 45090 19756 45310 19761
rect 45834 19961 46054 19966
rect 45834 19761 45844 19961
rect 46044 19761 46054 19961
rect 45834 19756 46054 19761
rect 46578 19961 46798 19966
rect 46578 19761 46588 19961
rect 46788 19761 46798 19961
rect 46578 19756 46798 19761
rect 47322 19961 47542 19966
rect 47322 19761 47332 19961
rect 47532 19761 47542 19961
rect 47322 19756 47542 19761
rect 48066 19961 48286 19966
rect 48066 19761 48076 19961
rect 48276 19761 48286 19961
rect 48066 19756 48286 19761
rect 48810 19961 49030 19966
rect 48810 19761 48820 19961
rect 49020 19761 49030 19961
rect 48810 19756 49030 19761
rect 49554 19961 49774 19966
rect 49554 19761 49564 19961
rect 49764 19761 49774 19961
rect 49554 19756 49774 19761
rect 46908 17525 47210 17530
rect 46908 17253 46918 17525
rect 47200 17253 47210 17525
rect 46908 16585 47210 17253
rect 47652 17525 47954 17530
rect 47652 17253 47662 17525
rect 47944 17253 47954 17525
rect 47652 16585 47954 17253
rect 48396 17525 48698 17530
rect 48396 17253 48406 17525
rect 48688 17253 48698 17525
rect 48396 16585 48698 17253
rect 49140 17525 49442 17530
rect 49140 17253 49150 17525
rect 49432 17253 49442 17525
rect 49140 16585 49442 17253
rect 45556 16470 45744 16475
rect 45556 16304 45566 16470
rect 45734 16304 45744 16470
rect 45556 16299 45744 16304
rect 45556 16070 45744 16075
rect 45556 15904 45566 16070
rect 45734 15904 45744 16070
rect 45556 15899 45744 15904
rect 45556 15670 45744 15675
rect 45556 15504 45566 15670
rect 45734 15504 45744 15670
rect 45556 15499 45744 15504
rect 46648 15483 49632 16585
rect 45842 15117 46144 15122
rect 45842 14845 45852 15117
rect 46134 14845 46144 15117
rect 45842 14840 46144 14845
rect 46648 14743 50144 15483
rect 45954 14453 46458 14458
rect 45954 13953 45964 14453
rect 46448 14345 46458 14453
rect 46648 14345 49632 14743
rect 46448 14089 49632 14345
rect 46448 13953 46458 14089
rect 45954 13948 46458 13953
rect 46648 13585 49632 14089
rect 46910 13343 47212 13585
rect 46910 13071 46920 13343
rect 47202 13071 47212 13343
rect 46910 13066 47212 13071
rect 47654 13343 47956 13585
rect 47654 13071 47664 13343
rect 47946 13071 47956 13343
rect 47654 13066 47956 13071
rect 48398 13343 48700 13585
rect 48398 13071 48408 13343
rect 48690 13071 48700 13343
rect 48398 13066 48700 13071
rect 49142 13343 49444 13585
rect 49142 13071 49152 13343
rect 49434 13071 49444 13343
rect 49142 13066 49444 13071
rect 39508 10715 39728 10720
rect 39508 10515 39518 10715
rect 39718 10515 39728 10715
rect 39508 10510 39728 10515
rect 40252 10715 40472 10720
rect 40252 10515 40262 10715
rect 40462 10515 40472 10715
rect 40252 10510 40472 10515
rect 40996 10715 41216 10720
rect 40996 10515 41006 10715
rect 41206 10515 41216 10715
rect 40996 10510 41216 10515
rect 41740 10715 41960 10720
rect 41740 10515 41750 10715
rect 41950 10515 41960 10715
rect 41740 10510 41960 10515
rect 42484 10715 42704 10720
rect 42484 10515 42494 10715
rect 42694 10515 42704 10715
rect 42484 10510 42704 10515
rect 43228 10715 43448 10720
rect 43228 10515 43238 10715
rect 43438 10515 43448 10715
rect 43228 10510 43448 10515
rect 43972 10715 44192 10720
rect 43972 10515 43982 10715
rect 44182 10515 44192 10715
rect 43972 10510 44192 10515
rect 44716 10715 44936 10720
rect 44716 10515 44726 10715
rect 44926 10515 44936 10715
rect 44716 10510 44936 10515
rect 45088 10715 45308 10720
rect 45088 10515 45098 10715
rect 45298 10515 45308 10715
rect 45088 10510 45308 10515
rect 45832 10715 46052 10720
rect 45832 10515 45842 10715
rect 46042 10515 46052 10715
rect 45832 10510 46052 10515
rect 46576 10715 46796 10720
rect 46576 10515 46586 10715
rect 46786 10515 46796 10715
rect 46576 10510 46796 10515
rect 47320 10715 47540 10720
rect 47320 10515 47330 10715
rect 47530 10515 47540 10715
rect 47320 10510 47540 10515
rect 48064 10715 48284 10720
rect 48064 10515 48074 10715
rect 48274 10515 48284 10715
rect 48064 10510 48284 10515
rect 48808 10715 49028 10720
rect 48808 10515 48818 10715
rect 49018 10515 49028 10715
rect 48808 10510 49028 10515
rect 49552 10715 49772 10720
rect 49552 10515 49562 10715
rect 49762 10515 49772 10715
rect 49552 10510 49772 10515
rect 50296 10715 50516 10720
rect 50296 10515 50306 10715
rect 50506 10515 50516 10715
rect 50296 10510 50516 10515
rect 51040 10715 51260 10720
rect 51040 10515 51050 10715
rect 51250 10515 51260 10715
rect 51040 10510 51260 10515
rect 39508 9350 39728 9355
rect 39508 9150 39518 9350
rect 39718 9150 39728 9350
rect 39508 9145 39728 9150
rect 40252 9350 40472 9355
rect 40252 9150 40262 9350
rect 40462 9150 40472 9350
rect 40252 9145 40472 9150
rect 40996 9350 41216 9355
rect 40996 9150 41006 9350
rect 41206 9150 41216 9350
rect 40996 9145 41216 9150
rect 41740 9350 41960 9355
rect 41740 9150 41750 9350
rect 41950 9150 41960 9350
rect 41740 9145 41960 9150
rect 42484 9350 42704 9355
rect 42484 9150 42494 9350
rect 42694 9150 42704 9350
rect 42484 9145 42704 9150
rect 43228 9350 43448 9355
rect 43228 9150 43238 9350
rect 43438 9150 43448 9350
rect 43228 9145 43448 9150
rect 43972 9350 44192 9355
rect 43972 9150 43982 9350
rect 44182 9150 44192 9350
rect 43972 9145 44192 9150
rect 44716 9350 44936 9355
rect 44716 9150 44726 9350
rect 44926 9150 44936 9350
rect 44716 9145 44936 9150
rect 45088 9350 45308 9355
rect 45088 9150 45098 9350
rect 45298 9150 45308 9350
rect 45088 9145 45308 9150
rect 45832 9350 46052 9355
rect 45832 9150 45842 9350
rect 46042 9150 46052 9350
rect 45832 9145 46052 9150
rect 46576 9350 46796 9355
rect 46576 9150 46586 9350
rect 46786 9150 46796 9350
rect 46576 9145 46796 9150
rect 47320 9350 47540 9355
rect 47320 9150 47330 9350
rect 47530 9150 47540 9350
rect 47320 9145 47540 9150
rect 48064 9350 48284 9355
rect 48064 9150 48074 9350
rect 48274 9150 48284 9350
rect 48064 9145 48284 9150
rect 48808 9350 49028 9355
rect 48808 9150 48818 9350
rect 49018 9150 49028 9350
rect 48808 9145 49028 9150
rect 49552 9350 49772 9355
rect 49552 9150 49562 9350
rect 49762 9150 49772 9350
rect 49552 9145 49772 9150
rect 50296 9350 50516 9355
rect 50296 9150 50306 9350
rect 50506 9150 50516 9350
rect 50296 9145 50516 9150
rect 51040 9350 51260 9355
rect 51040 9150 51050 9350
rect 51250 9150 51260 9350
rect 51040 9145 51260 9150
rect 46910 6794 47212 6799
rect 46910 6522 46920 6794
rect 47202 6522 47212 6794
rect 46910 6280 47212 6522
rect 47654 6794 47956 6799
rect 47654 6522 47664 6794
rect 47946 6522 47956 6794
rect 47654 6280 47956 6522
rect 48398 6794 48700 6799
rect 48398 6522 48408 6794
rect 48690 6522 48700 6794
rect 48398 6280 48700 6522
rect 49142 6794 49444 6799
rect 49142 6522 49152 6794
rect 49434 6522 49444 6794
rect 49142 6280 49444 6522
rect 40236 6259 40402 6264
rect 40236 6109 40246 6259
rect 40392 6109 40402 6259
rect 40236 6104 40402 6109
rect 45628 6135 46132 6140
rect 40236 5859 40402 5864
rect 40236 5709 40246 5859
rect 40392 5709 40402 5859
rect 40236 5704 40402 5709
rect 44152 5719 44318 5724
rect 44152 5569 44162 5719
rect 44308 5569 44318 5719
rect 45628 5635 45638 6135
rect 46122 6057 46132 6135
rect 46648 6057 49632 6280
rect 46122 5693 49632 6057
rect 46122 5635 46132 5693
rect 45628 5630 46132 5635
rect 44152 5564 44318 5569
rect 40236 5459 40402 5464
rect 40236 5309 40246 5459
rect 40392 5309 40402 5459
rect 40236 5304 40402 5309
rect 44152 5319 44318 5324
rect 44152 5169 44162 5319
rect 44308 5169 44318 5319
rect 44152 5164 44318 5169
rect 46648 5122 49632 5693
rect 40236 5059 40402 5064
rect 40236 4909 40246 5059
rect 40392 4909 40402 5059
rect 45842 5020 46144 5025
rect 40236 4904 40402 4909
rect 44152 4919 44318 4924
rect 44152 4769 44162 4919
rect 44308 4769 44318 4919
rect 44152 4764 44318 4769
rect 45842 4748 45852 5020
rect 46134 4748 46144 5020
rect 45842 4743 46144 4748
rect 44152 4519 44318 4524
rect 44152 4369 44162 4519
rect 44308 4369 44318 4519
rect 44152 4364 44318 4369
rect 46648 4382 50144 5122
rect 45546 4306 45740 4311
rect 45546 4132 45556 4306
rect 45730 4132 45740 4306
rect 45546 4127 45740 4132
rect 45546 3906 45740 3911
rect 45546 3732 45556 3906
rect 45730 3732 45740 3906
rect 45546 3727 45740 3732
rect 45546 3506 45740 3511
rect 45546 3332 45556 3506
rect 45730 3332 45740 3506
rect 45546 3327 45740 3332
rect 46648 3280 49632 4382
rect 46908 2612 47210 3280
rect 46908 2340 46918 2612
rect 47200 2340 47210 2612
rect 46908 2335 47210 2340
rect 47652 2612 47954 3280
rect 47652 2340 47662 2612
rect 47944 2340 47954 2612
rect 47652 2335 47954 2340
rect 48396 2612 48698 3280
rect 48396 2340 48406 2612
rect 48688 2340 48698 2612
rect 48396 2335 48698 2340
rect 49140 2612 49442 3280
rect 49140 2340 49150 2612
rect 49432 2340 49442 2612
rect 49140 2335 49442 2340
rect 40646 104 40866 109
rect 40646 -96 40656 104
rect 40856 -96 40866 104
rect 40646 -101 40866 -96
rect 41370 104 41590 109
rect 41370 -96 41380 104
rect 41580 -96 41590 104
rect 41370 -101 41590 -96
rect 42114 104 42334 109
rect 42114 -96 42124 104
rect 42324 -96 42334 104
rect 42114 -101 42334 -96
rect 42858 104 43078 109
rect 42858 -96 42868 104
rect 43068 -96 43078 104
rect 42858 -101 43078 -96
rect 43602 104 43822 109
rect 43602 -96 43612 104
rect 43812 -96 43822 104
rect 43602 -101 43822 -96
rect 44346 104 44566 109
rect 44346 -96 44356 104
rect 44556 -96 44566 104
rect 44346 -101 44566 -96
rect 45090 104 45310 109
rect 45090 -96 45100 104
rect 45300 -96 45310 104
rect 45090 -101 45310 -96
rect 45834 104 46054 109
rect 45834 -96 45844 104
rect 46044 -96 46054 104
rect 45834 -101 46054 -96
rect 46578 104 46798 109
rect 46578 -96 46588 104
rect 46788 -96 46798 104
rect 46578 -101 46798 -96
rect 47322 104 47542 109
rect 47322 -96 47332 104
rect 47532 -96 47542 104
rect 47322 -101 47542 -96
rect 48066 104 48286 109
rect 48066 -96 48076 104
rect 48276 -96 48286 104
rect 48066 -101 48286 -96
rect 48810 104 49030 109
rect 48810 -96 48820 104
rect 49020 -96 49030 104
rect 48810 -101 49030 -96
rect 49554 104 49774 109
rect 49554 -96 49564 104
rect 49764 -96 49774 104
rect 49554 -101 49774 -96
<< via3 >>
rect 40656 19761 40856 19961
rect 41380 19761 41580 19961
rect 42124 19761 42324 19961
rect 42868 19761 43068 19961
rect 43612 19761 43812 19961
rect 44356 19761 44556 19961
rect 45100 19761 45300 19961
rect 45844 19761 46044 19961
rect 46588 19761 46788 19961
rect 47332 19761 47532 19961
rect 48076 19761 48276 19961
rect 48820 19761 49020 19961
rect 49564 19761 49764 19961
rect 45566 16304 45734 16470
rect 45566 15904 45734 16070
rect 45566 15504 45734 15670
rect 45852 14845 46134 15117
rect 39518 10515 39718 10715
rect 40262 10515 40462 10715
rect 41006 10515 41206 10715
rect 41750 10515 41950 10715
rect 42494 10515 42694 10715
rect 43238 10515 43438 10715
rect 43982 10515 44182 10715
rect 44726 10515 44926 10715
rect 45098 10515 45298 10715
rect 45842 10515 46042 10715
rect 46586 10515 46786 10715
rect 47330 10515 47530 10715
rect 48074 10515 48274 10715
rect 48818 10515 49018 10715
rect 49562 10515 49762 10715
rect 50306 10515 50506 10715
rect 51050 10515 51250 10715
rect 39518 9150 39718 9350
rect 40262 9150 40462 9350
rect 41006 9150 41206 9350
rect 41750 9150 41950 9350
rect 42494 9150 42694 9350
rect 43238 9150 43438 9350
rect 43982 9150 44182 9350
rect 44726 9150 44926 9350
rect 45098 9150 45298 9350
rect 45842 9150 46042 9350
rect 46586 9150 46786 9350
rect 47330 9150 47530 9350
rect 48074 9150 48274 9350
rect 48818 9150 49018 9350
rect 49562 9150 49762 9350
rect 50306 9150 50506 9350
rect 51050 9150 51250 9350
rect 40246 6109 40392 6259
rect 40246 5709 40392 5859
rect 44162 5569 44308 5719
rect 40246 5309 40392 5459
rect 44162 5169 44308 5319
rect 40246 4909 40392 5059
rect 44162 4769 44308 4919
rect 45852 4748 46134 5020
rect 44162 4369 44308 4519
rect 45556 4132 45730 4306
rect 45556 3732 45730 3906
rect 45556 3332 45730 3506
rect 40656 -96 40856 104
rect 41380 -96 41580 104
rect 42124 -96 42324 104
rect 42868 -96 43068 104
rect 43612 -96 43812 104
rect 44356 -96 44556 104
rect 45100 -96 45300 104
rect 45844 -96 46044 104
rect 46588 -96 46788 104
rect 47332 -96 47532 104
rect 48076 -96 48276 104
rect 48820 -96 49020 104
rect 49564 -96 49764 104
<< mimcap >>
rect 46748 16445 49548 16485
rect 46748 13725 46788 16445
rect 49508 13725 49548 16445
rect 46748 13685 49548 13725
rect 46748 6140 49548 6180
rect 46748 3420 46788 6140
rect 49508 3420 49548 6140
rect 46748 3380 49548 3420
<< mimcapcontact >>
rect 46788 13725 49508 16445
rect 46788 3420 49508 6140
<< metal4 >>
rect 38912 19961 51436 20741
rect 38912 19761 40656 19961
rect 40856 19761 41380 19961
rect 41580 19761 42124 19961
rect 42324 19761 42868 19961
rect 43068 19761 43612 19961
rect 43812 19761 44356 19961
rect 44556 19761 45100 19961
rect 45300 19761 45844 19961
rect 46044 19761 46588 19961
rect 46788 19761 47332 19961
rect 47532 19761 48076 19961
rect 48276 19761 48820 19961
rect 49020 19761 49564 19961
rect 49764 19761 51436 19961
rect 38912 19737 51436 19761
rect 45530 16470 45768 19737
rect 45530 16304 45566 16470
rect 45734 16304 45768 16470
rect 45530 16070 45768 16304
rect 45530 15904 45566 16070
rect 45734 15904 45768 16070
rect 45530 15670 45768 15904
rect 45530 15504 45566 15670
rect 45734 15504 45768 15670
rect 45530 15395 45768 15504
rect 46787 16445 49509 16446
rect 45851 15117 46135 15118
rect 45851 14845 45852 15117
rect 46134 15091 46135 15117
rect 46787 15091 46788 16445
rect 46134 14873 46788 15091
rect 46134 14845 46135 14873
rect 45851 14844 46135 14845
rect 46787 13725 46788 14873
rect 49508 13725 49509 16445
rect 46787 13724 49509 13725
rect 38912 10715 51436 10741
rect 38912 10515 39518 10715
rect 39718 10515 40262 10715
rect 40462 10515 41006 10715
rect 41206 10515 41750 10715
rect 41950 10515 42494 10715
rect 42694 10515 43238 10715
rect 43438 10515 43982 10715
rect 44182 10515 44726 10715
rect 44926 10515 45098 10715
rect 45298 10515 45842 10715
rect 46042 10515 46586 10715
rect 46786 10515 47330 10715
rect 47530 10515 48074 10715
rect 48274 10515 48818 10715
rect 49018 10515 49562 10715
rect 49762 10515 50306 10715
rect 50506 10515 51050 10715
rect 51250 10515 51436 10715
rect 38912 9350 51436 10515
rect 38912 9150 39518 9350
rect 39718 9150 40262 9350
rect 40462 9150 41006 9350
rect 41206 9150 41750 9350
rect 41950 9150 42494 9350
rect 42694 9150 43238 9350
rect 43438 9150 43982 9350
rect 44182 9150 44726 9350
rect 44926 9150 45098 9350
rect 45298 9150 45842 9350
rect 46042 9150 46586 9350
rect 46786 9150 47330 9350
rect 47530 9150 48074 9350
rect 48274 9150 48818 9350
rect 49018 9150 49562 9350
rect 49762 9150 50306 9350
rect 50506 9150 51050 9350
rect 51250 9150 51436 9350
rect 38912 9124 51436 9150
rect 40148 6259 40478 6303
rect 40148 6109 40246 6259
rect 40392 6109 40478 6259
rect 40148 5859 40478 6109
rect 40148 5709 40246 5859
rect 40392 5709 40478 5859
rect 46787 6140 49509 6141
rect 40148 5459 40478 5709
rect 40148 5309 40246 5459
rect 40392 5309 40478 5459
rect 40148 5059 40478 5309
rect 40148 4909 40246 5059
rect 40392 4909 40478 5059
rect 40148 128 40478 4909
rect 44122 5719 44344 5801
rect 44122 5569 44162 5719
rect 44308 5569 44344 5719
rect 44122 5319 44344 5569
rect 44122 5169 44162 5319
rect 44308 5169 44344 5319
rect 44122 4919 44344 5169
rect 44122 4769 44162 4919
rect 44308 4769 44344 4919
rect 44122 4519 44344 4769
rect 45851 5020 46135 5021
rect 45851 4748 45852 5020
rect 46134 4992 46135 5020
rect 46787 4992 46788 6140
rect 46134 4774 46788 4992
rect 46134 4748 46135 4774
rect 45851 4747 46135 4748
rect 44122 4369 44162 4519
rect 44308 4369 44344 4519
rect 44122 128 44344 4369
rect 45522 4306 45760 4470
rect 45522 4132 45556 4306
rect 45730 4132 45760 4306
rect 45522 3906 45760 4132
rect 45522 3732 45556 3906
rect 45730 3732 45760 3906
rect 45522 3506 45760 3732
rect 45522 3332 45556 3506
rect 45730 3332 45760 3506
rect 46787 3420 46788 4774
rect 49508 3420 49509 6140
rect 46787 3419 49509 3420
rect 45522 128 45760 3332
rect 38912 104 51436 128
rect 38912 -96 40656 104
rect 40856 -96 41380 104
rect 41580 -96 42124 104
rect 42324 -96 42868 104
rect 43068 -96 43612 104
rect 43812 -96 44356 104
rect 44556 -96 45100 104
rect 45300 -96 45844 104
rect 46044 -96 46588 104
rect 46788 -96 47332 104
rect 47532 -96 48076 104
rect 48276 -96 48820 104
rect 49020 -96 49564 104
rect 49764 -96 51436 104
rect 38912 -876 51436 -96
<< end >>
