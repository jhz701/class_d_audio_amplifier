magic
tech sky130A
magscale 1 2
timestamp 1629189290
<< nwell >>
rect 368 1522 402 1660
rect 368 -1618 402 -1500
<< pwell >>
rect 417 -5206 1137 -3010
rect 5573 -5846 6293 -3650
<< psubdiff >>
rect 453 -3080 549 -3046
rect 1005 -3080 1101 -3046
rect 453 -3142 487 -3080
rect 1067 -3142 1101 -3080
rect 453 -5136 487 -5074
rect 1067 -5136 1101 -5074
rect 453 -5170 549 -5136
rect 1005 -5170 1101 -5136
rect 5609 -3720 5705 -3686
rect 6161 -3720 6257 -3686
rect 5609 -3782 5643 -3720
rect 6223 -3782 6257 -3720
rect 5609 -5776 5643 -5714
rect 6223 -5776 6257 -5714
rect 5609 -5810 5705 -5776
rect 6161 -5810 6257 -5776
<< psubdiffcont >>
rect 549 -3080 1005 -3046
rect 453 -5074 487 -3142
rect 1067 -5074 1101 -3142
rect 549 -5170 1005 -5136
rect 5705 -3720 6161 -3686
rect 5609 -5714 5643 -3782
rect 6223 -5714 6257 -3782
rect 5705 -5810 6161 -5776
<< xpolycontact >>
rect 583 -3608 653 -3176
rect 583 -5040 653 -4608
rect 901 -3608 971 -3176
rect 901 -5040 971 -4608
rect 5739 -4248 5809 -3816
rect 5739 -5680 5809 -5248
rect 6057 -4248 6127 -3816
rect 6057 -5680 6127 -5248
<< xpolyres >>
rect 583 -4608 653 -3608
rect 901 -4608 971 -3608
rect 5739 -5248 5809 -4248
rect 6057 -5248 6127 -4248
<< locali >>
rect 453 -3080 549 -3046
rect 1005 -3080 1101 -3046
rect 453 -3142 487 -3080
rect 1067 -3142 1101 -3080
rect 5609 -3720 5705 -3686
rect 6161 -3720 6257 -3686
rect 5609 -3782 5643 -3720
rect 6223 -3782 6257 -3720
rect 453 -5136 487 -5074
rect 1067 -5136 1101 -5074
rect 453 -5170 549 -5136
rect 1005 -5170 1101 -5136
rect 5609 -5776 5643 -5714
rect 6223 -5776 6257 -5714
rect 5609 -5810 5705 -5776
rect 6161 -5810 6257 -5776
<< viali >>
rect 599 -3591 637 -3194
rect 917 -3591 955 -3194
rect 1048 -3763 1067 -3697
rect 1067 -3763 1101 -3697
rect 1101 -3763 1120 -3697
rect 1048 -4161 1067 -4097
rect 1067 -4161 1101 -4097
rect 1101 -4161 1120 -4097
rect 5755 -4231 5793 -3834
rect 5590 -4303 5609 -4237
rect 5609 -4303 5643 -4237
rect 5643 -4303 5662 -4237
rect 6073 -4231 6111 -3834
rect 1048 -4561 1067 -4497
rect 1067 -4561 1101 -4497
rect 1101 -4561 1120 -4497
rect 599 -5022 637 -4625
rect 917 -5022 955 -4625
rect 5590 -4701 5609 -4637
rect 5609 -4701 5643 -4637
rect 5643 -4701 5662 -4637
rect 1048 -4961 1067 -4897
rect 1067 -4961 1101 -4897
rect 1101 -4961 1120 -4897
rect 5590 -5101 5609 -5037
rect 5609 -5101 5643 -5037
rect 5643 -5101 5662 -5037
rect 5590 -5501 5609 -5437
rect 5609 -5501 5643 -5437
rect 5643 -5501 5662 -5437
rect 5755 -5662 5793 -5265
rect 6073 -5662 6111 -5265
<< metal1 >>
rect -618 7192 -608 7700
rect -122 7192 -112 7700
rect -532 -3218 -194 7192
rect 368 1522 402 1660
rect 368 -1618 402 -1500
rect 582 -3194 654 -3177
rect -532 -3219 342 -3218
rect 582 -3219 599 -3194
rect -532 -3535 599 -3219
rect -532 -3536 342 -3535
rect 593 -3591 599 -3535
rect 637 -3421 654 -3194
rect 902 -3194 970 -3177
rect 637 -3591 643 -3421
rect 593 -3603 643 -3591
rect 902 -3591 917 -3194
rect 955 -3269 970 -3194
rect 1190 -3269 1200 -3241
rect 955 -3475 1200 -3269
rect 955 -3591 970 -3475
rect 1190 -3515 1200 -3475
rect 1482 -3515 1492 -3241
rect 5684 -3359 5694 -3085
rect 5976 -3359 5986 -3085
rect 902 -3607 970 -3591
rect 1314 -3691 1324 -3657
rect 1036 -3697 1324 -3691
rect 1036 -3763 1048 -3697
rect 1120 -3763 1324 -3697
rect 1036 -3767 1324 -3763
rect 1036 -3769 1132 -3767
rect 1314 -3807 1324 -3767
rect 1470 -3807 1480 -3657
rect 5738 -3834 5810 -3359
rect 6706 -3815 6716 -3781
rect 1314 -4091 1324 -4057
rect 1036 -4097 1324 -4091
rect 1036 -4161 1048 -4097
rect 1120 -4161 1324 -4097
rect 1036 -4167 1324 -4161
rect 1314 -4207 1324 -4167
rect 1470 -4207 1480 -4057
rect 5738 -4061 5755 -3834
rect 5230 -4347 5240 -4197
rect 5386 -4231 5396 -4197
rect 5749 -4231 5755 -4061
rect 5793 -4061 5810 -3834
rect 6056 -3834 6716 -3815
rect 5793 -4231 5799 -4061
rect 5386 -4237 5674 -4231
rect 5386 -4303 5590 -4237
rect 5662 -4303 5674 -4237
rect 5749 -4243 5799 -4231
rect 6056 -4231 6073 -3834
rect 6111 -4231 6716 -3834
rect 6056 -4249 6716 -4231
rect 6706 -4281 6716 -4249
rect 7200 -4281 7210 -3781
rect 5386 -4307 5674 -4303
rect 5386 -4347 5396 -4307
rect 5578 -4309 5674 -4307
rect 1314 -4491 1324 -4457
rect 1036 -4497 1324 -4491
rect 1036 -4561 1048 -4497
rect 1120 -4561 1324 -4497
rect 1036 -4567 1324 -4561
rect 1314 -4607 1324 -4567
rect 1470 -4607 1480 -4457
rect 582 -4625 972 -4607
rect 582 -5022 599 -4625
rect 637 -5022 917 -4625
rect 955 -5022 972 -4625
rect 5230 -4747 5240 -4597
rect 5386 -4631 5396 -4597
rect 5386 -4637 5674 -4631
rect 5386 -4701 5590 -4637
rect 5662 -4701 5674 -4637
rect 5386 -4707 5674 -4701
rect 5386 -4747 5396 -4707
rect 1314 -4891 1324 -4857
rect 1036 -4897 1324 -4891
rect 1036 -4961 1048 -4897
rect 1120 -4961 1324 -4897
rect 1036 -4967 1324 -4961
rect 1314 -5007 1324 -4967
rect 1470 -5007 1480 -4857
rect 582 -5041 972 -5022
rect 5230 -5147 5240 -4997
rect 5386 -5031 5396 -4997
rect 5386 -5037 5674 -5031
rect 5386 -5101 5590 -5037
rect 5662 -5101 5674 -5037
rect 5386 -5107 5674 -5101
rect 5386 -5147 5396 -5107
rect 5738 -5265 6128 -5247
rect 5230 -5547 5240 -5397
rect 5386 -5431 5396 -5397
rect 5386 -5437 5674 -5431
rect 5386 -5501 5590 -5437
rect 5662 -5501 5674 -5437
rect 5386 -5507 5674 -5501
rect 5386 -5547 5396 -5507
rect 5738 -5662 5755 -5265
rect 5793 -5662 6073 -5265
rect 6111 -5662 6128 -5265
rect 5738 -5681 6128 -5662
<< via1 >>
rect -608 7192 -122 7700
rect 1200 -3515 1482 -3241
rect 5694 -3359 5976 -3085
rect 1324 -3807 1470 -3657
rect 1324 -4207 1470 -4057
rect 5240 -4347 5386 -4197
rect 6716 -4281 7200 -3781
rect 1324 -4607 1470 -4457
rect 5240 -4747 5386 -4597
rect 1324 -5007 1470 -4857
rect 5240 -5147 5386 -4997
rect 5240 -5547 5386 -5397
<< metal2 >>
rect -608 7700 -122 7710
rect -122 7576 1792 7676
rect -608 7182 -122 7192
rect 7042 4537 7526 4547
rect 5500 4179 7042 4391
rect 5500 3303 5680 4179
rect 7042 4027 7526 4037
rect 4468 3175 5680 3303
rect 5694 -3085 5976 -3075
rect 1200 -3241 1482 -3141
rect 4492 -3277 5694 -3143
rect 5694 -3369 5976 -3359
rect 1200 -3525 1482 -3515
rect 1324 -3657 1470 -3647
rect 1324 -3817 1470 -3807
rect 6716 -3781 7200 -3771
rect 1324 -4057 1470 -4047
rect 1324 -4217 1470 -4207
rect 5240 -4197 5386 -4187
rect 6716 -4291 7200 -4281
rect 5240 -4357 5386 -4347
rect 1324 -4457 1470 -4447
rect 1324 -4617 1470 -4607
rect 5240 -4597 5386 -4587
rect 5240 -4757 5386 -4747
rect 1324 -4857 1470 -4847
rect 1324 -5017 1470 -5007
rect 5240 -4997 5386 -4987
rect 5240 -5157 5386 -5147
rect 5240 -5397 5386 -5387
rect 5240 -5557 5386 -5547
rect 1754 -7628 2044 -7556
<< via2 >>
rect 7042 4037 7526 4537
rect 1324 -3807 1470 -3657
rect 1324 -4207 1470 -4057
rect 5240 -4347 5386 -4197
rect 6716 -4281 7200 -3781
rect 1324 -4607 1470 -4457
rect 5240 -4747 5386 -4597
rect 1324 -5007 1470 -4857
rect 5240 -5147 5386 -4997
rect 5240 -5547 5386 -5397
<< metal3 >>
rect 10842 4852 11180 5292
rect 7032 4537 7536 4542
rect 7032 4037 7042 4537
rect 7526 4429 7536 4537
rect 7526 4173 8112 4429
rect 7526 4037 7536 4173
rect 7032 4032 7536 4037
rect 1314 -3657 1480 -3652
rect 1314 -3807 1324 -3657
rect 1470 -3807 1480 -3657
rect 1314 -3812 1480 -3807
rect 6706 -3781 7210 -3776
rect 1314 -4057 1480 -4052
rect 1314 -4207 1324 -4057
rect 1470 -4207 1480 -4057
rect 1314 -4212 1480 -4207
rect 5230 -4197 5396 -4192
rect 5230 -4347 5240 -4197
rect 5386 -4347 5396 -4197
rect 6706 -4281 6716 -3781
rect 7200 -3859 7210 -3781
rect 7200 -4223 7910 -3859
rect 7200 -4281 7210 -4223
rect 6706 -4286 7210 -4281
rect 5230 -4352 5396 -4347
rect 1314 -4457 1480 -4452
rect 1314 -4607 1324 -4457
rect 1470 -4607 1480 -4457
rect 1314 -4612 1480 -4607
rect 5230 -4597 5396 -4592
rect 5230 -4747 5240 -4597
rect 5386 -4747 5396 -4597
rect 5230 -4752 5396 -4747
rect 1314 -4857 1480 -4852
rect 1314 -5007 1324 -4857
rect 1470 -5007 1480 -4857
rect 1314 -5012 1480 -5007
rect 5230 -4997 5396 -4992
rect 5230 -5147 5240 -4997
rect 5386 -5147 5396 -4997
rect 5230 -5152 5396 -5147
rect 5230 -5397 5396 -5392
rect 5230 -5547 5240 -5397
rect 5386 -5547 5396 -5397
rect 10770 -5522 11014 -4974
rect 5230 -5552 5396 -5547
<< via3 >>
rect 1324 -3807 1470 -3657
rect 1324 -4207 1470 -4057
rect 5240 -4347 5386 -4197
rect 1324 -4607 1470 -4457
rect 5240 -4747 5386 -4597
rect 1324 -5007 1470 -4857
rect 5240 -5147 5386 -4997
rect 5240 -5547 5386 -5397
<< metal4 >>
rect 11650 9904 17120 10772
rect 258 -378 12038 336
rect 1226 -3657 1556 -3613
rect 1226 -3807 1324 -3657
rect 1470 -3807 1556 -3657
rect 1226 -4057 1556 -3807
rect 1226 -4207 1324 -4057
rect 1470 -4207 1556 -4057
rect 1226 -4457 1556 -4207
rect 1226 -4607 1324 -4457
rect 1470 -4607 1556 -4457
rect 1226 -4857 1556 -4607
rect 1226 -5007 1324 -4857
rect 1470 -5007 1556 -4857
rect 1226 -10227 1556 -5007
rect 5200 -4197 5422 -4115
rect 5200 -4347 5240 -4197
rect 5386 -4347 5422 -4197
rect 5200 -4597 5422 -4347
rect 5200 -4747 5240 -4597
rect 5386 -4747 5422 -4597
rect 5200 -4997 5422 -4747
rect 5200 -5147 5240 -4997
rect 5386 -5147 5422 -4997
rect 5200 -5397 5422 -5147
rect 5200 -5547 5240 -5397
rect 5386 -5547 5422 -5397
rect 5200 -10417 5422 -5547
rect 15930 -9812 17024 9904
rect 11898 -10766 17424 -9812
use OTA_revised  OTA_revised_1 ~/magic/class_d_audio_amplifier/OTA
timestamp 1629189150
transform 1 0 918 0 1 -2080
box -928 -8712 11596 2292
use OTA_revised  OTA_revised_0
timestamp 1629189150
transform 1 0 918 0 -1 2113
box -928 -8712 11596 2292
<< labels >>
flabel metal4 4606 -30 4606 -30 0 FreeSans 8000 0 0 0 vdd
port 0 nsew
flabel metal4 16216 2364 16216 2364 0 FreeSans 8000 0 0 0 vss
port 5 nsew
flabel metal3 10944 5046 10944 5046 0 FreeSans 8000 0 0 0 vp
port 7 nsew
flabel metal3 10912 -5226 10912 -5226 0 FreeSans 8000 0 0 0 vn
port 6 nsew
flabel metal1 -312 4004 -312 4004 0 FreeSans 8000 0 0 0 vi
port 3 nsew
flabel metal2 1874 -7600 1874 -7600 0 FreeSans 8000 0 0 0 vref
port 4 nsew
flabel metal1 382 1596 382 1596 0 FreeSans 8000 0 0 0 vbias1
port 1 nsew
flabel metal1 388 -1546 388 -1546 0 FreeSans 8000 0 0 0 vbias2
port 2 nsew
<< end >>
