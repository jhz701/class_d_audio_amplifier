* NGSPICE file created from /home/eda/magic/class_d_audio_amplifier/comparator/comparator_revised.ext - technology: sky130A

.subckt comparator_revised_post vdd vp vn vbias vss vout
X0 w_20679_4119.t42 vbias.t48 vdd.t95 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1 w_20679_4119.t41 vbias.t49 vdd.t94 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2 w_20679_4119.t18 vp.t0 a_21819_2107.t15 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3 vout.t63 a_21819_2107.t32 vss.t78 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4 vout.t111 vbias.t50 vdd.t93 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5 vout.t62 a_21819_2107.t33 vss.t77 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6 vdd.t92 vbias.t46 vbias.t47 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7 vdd.t91 vbias.t51 vout.t110 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8 vout.t109 vbias.t52 vdd.t90 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9 a_21819_2107.t16 a_20875_2019.t48 vss.t80 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10 w_20679_4119.t55 vn.t0 a_20875_2019.t47 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X11 a_21819_2107.t17 a_20875_2019.t49 vss.t81 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X12 vss.t76 a_21819_2107.t34 vout.t61 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X13 w_20679_4119.t16 vp.t1 a_21819_2107.t14 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X14 a_21819_2107.t13 vp.t2 w_20679_4119.t17 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X15 vdd.t89 vbias.t53 vout.t108 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X16 vbias.t45 vbias.t44 vdd.t88 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X17 vout.t60 a_21819_2107.t35 vss.t75 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X18 vdd.t87 vbias.t42 vbias.t43 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X19 vbias.t41 vbias.t40 vdd.t86 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X20 vout.t107 vbias.t54 vdd.t85 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X21 vbias.t39 vbias.t38 vdd.t84 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X22 vdd.t83 vbias.t55 vout.t106 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X23 vss.t74 a_21819_2107.t36 vout.t59 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X24 vout.t105 vbias.t56 vdd.t82 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X25 vdd.t81 vbias.t57 vout.t104 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X26 vout.t58 a_21819_2107.t37 vss.t73 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X27 vss.t72 a_21819_2107.t38 vout.t57 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X28 vout.t103 vbias.t58 vdd.t80 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X29 w_20679_4119.t53 vn.t1 a_20875_2019.t45 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X30 vout.t56 a_21819_2107.t39 vss.t71 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X31 vout.t55 a_21819_2107.t40 vss.t70 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X32 a_21819_2107.t12 vp.t3 w_20679_4119.t4 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X33 vss.t69 a_21819_2107.t41 vout.t54 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X34 w_20679_4119.t3 vp.t4 a_21819_2107.t11 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X35 vss.t68 a_21819_2107.t42 vout.t53 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X36 vdd.t79 vbias.t59 vout.t102 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X37 vout.t52 a_21819_2107.t43 vss.t67 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X38 vss.t66 a_21819_2107.t44 vout.t51 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X39 vout.t101 vbias.t60 vdd.t78 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X40 vdd.t77 vbias.t61 vout.t100 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X41 w_20679_4119.t40 vbias.t62 vdd.t76 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X42 vdd.t75 vbias.t63 w_20679_4119.t39 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X43 a_20875_2019.t34 a_20875_2019.t33 vss.t79 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X44 vdd.t74 vbias.t36 vbias.t37 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X45 a_20875_2019.t32 a_20875_2019.t31 vss.t14 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X46 vss.t65 a_21819_2107.t45 vout.t50 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X47 vout.t99 vbias.t64 vdd.t73 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X48 a_20875_2019.t30 a_20875_2019.t29 vss.t13 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X49 a_20875_2019.t28 a_20875_2019.t27 vss.t12 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X50 a_21819_2107.t10 vp.t5 w_20679_4119.t15 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X51 vss.t64 a_21819_2107.t46 vout.t49 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X52 vss.t63 a_21819_2107.t47 vout.t48 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X53 w_20679_4119.t43 vp.t6 a_21819_2107.t9 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X54 vdd.t72 vbias.t34 vbias.t35 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X55 vdd.t71 vbias.t65 vout.t98 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X56 vss.t62 a_21819_2107.t48 vout.t47 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X57 w_20679_4119.t38 vbias.t66 vdd.t70 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X58 vdd.t69 vbias.t67 vout.t97 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X59 vdd.t68 vbias.t32 vbias.t33 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X60 vout.t46 a_21819_2107.t49 vss.t61 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X61 vss.t60 a_21819_2107.t50 vout.t45 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X62 vss.t82 a_20875_2019.t50 a_21819_2107.t18 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X63 vss.t83 a_20875_2019.t51 a_21819_2107.t19 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X64 vss.t59 a_21819_2107.t51 vout.t44 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X65 vout.t96 vbias.t68 vdd.t67 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X66 vss.t58 a_21819_2107.t52 vout.t43 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X67 vout.t42 a_21819_2107.t53 vss.t57 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X68 vout.t41 a_21819_2107.t54 vss.t56 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X69 vdd.t66 vbias.t69 vout.t95 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X70 vout.t40 a_21819_2107.t55 vss.t55 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X71 vss.t54 a_21819_2107.t56 vout.t39 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X72 vdd.t65 vbias.t30 vbias.t31 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X73 vdd.t64 vbias.t70 vout.t94 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X74 vdd.t63 vbias.t71 w_20679_4119.t37 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X75 vout.t93 vbias.t72 vdd.t62 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X76 vss.t11 a_20875_2019.t25 a_20875_2019.t26 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X77 vout.t92 vbias.t73 vdd.t61 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X78 a_21819_2107.t20 a_20875_2019.t52 vss.t84 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X79 vdd.t60 vbias.t74 vout.t91 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X80 vdd.t59 vbias.t75 vout.t90 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X81 a_21819_2107.t21 a_20875_2019.t53 vss.t85 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X82 a_20875_2019.t46 vn.t2 w_20679_4119.t54 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X83 vout.t38 a_21819_2107.t57 vss.t53 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X84 vss.t52 a_21819_2107.t58 vout.t37 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X85 a_20875_2019.t1 vn.t3 w_20679_4119.t1 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X86 vss.t51 a_21819_2107.t59 vout.t36 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X87 vss.t10 a_20875_2019.t23 a_20875_2019.t24 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X88 vdd.t58 vbias.t76 w_20679_4119.t36 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X89 vbias.t29 vbias.t28 vdd.t57 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X90 vdd.t56 vbias.t77 vout.t89 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X91 vdd.t55 vbias.t26 vbias.t27 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X92 w_20679_4119.t2 vn.t4 a_20875_2019.t2 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X93 vout.t35 a_21819_2107.t60 vss.t50 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X94 vss.t9 a_20875_2019.t21 a_20875_2019.t22 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X95 vout.t88 vbias.t78 vdd.t54 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X96 vdd.t53 vbias.t79 w_20679_4119.t35 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X97 vout.t34 a_21819_2107.t61 vss.t49 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X98 w_20679_4119.t34 vbias.t80 vdd.t52 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X99 vdd.t51 vbias.t81 vout.t87 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X100 vss.t86 a_20875_2019.t54 a_21819_2107.t22 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X101 vbias.t25 vbias.t24 vdd.t50 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X102 vss.t87 a_20875_2019.t55 a_21819_2107.t23 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X103 w_20679_4119.t44 vp.t7 a_21819_2107.t8 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X104 vout.t86 vbias.t82 vdd.t49 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X105 vss.t8 a_20875_2019.t19 a_20875_2019.t20 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X106 vout.t33 a_21819_2107.t62 vss.t48 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X107 vout.t32 a_21819_2107.t63 vss.t47 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X108 w_20679_4119.t33 vbias.t83 vdd.t48 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X109 vout.t31 a_21819_2107.t64 vss.t46 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X110 vdd.t47 vbias.t84 w_20679_4119.t32 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X111 w_20679_4119.t0 vn.t5 a_20875_2019.t0 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X112 vbias.t23 vbias.t22 vdd.t46 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X113 vout.t85 vbias.t85 vdd.t45 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X114 a_21819_2107.t24 a_20875_2019.t56 vss.t88 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X115 vout.t84 vbias.t86 vdd.t44 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X116 w_20679_4119.t31 vbias.t87 vdd.t43 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X117 vout.t83 vbias.t88 vdd.t42 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X118 a_21819_2107.t7 vp.t8 w_20679_4119.t45 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X119 vout.t30 a_21819_2107.t65 vss.t45 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X120 vout.t29 a_21819_2107.t66 vss.t44 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X121 vbias.t21 vbias.t20 vdd.t41 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X122 w_20679_4119.t5 vn.t6 a_20875_2019.t35 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X123 a_21819_2107.t25 a_20875_2019.t57 vss.t89 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X124 vss.t43 a_21819_2107.t67 vout.t28 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X125 vss.t42 a_21819_2107.t68 vout.t27 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X126 vdd.t40 vbias.t18 vbias.t19 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X127 vbias.t17 vbias.t16 vdd.t39 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X128 vdd.t38 vbias.t89 w_20679_4119.t30 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X129 vout.t82 vbias.t90 vdd.t37 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X130 vbias.t15 vbias.t14 vdd.t36 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X131 a_21819_2107.t6 vp.t9 w_20679_4119.t46 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X132 vdd.t35 vbias.t12 vbias.t13 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X133 vout.t26 a_21819_2107.t69 vss.t41 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X134 vss.t40 a_21819_2107.t70 vout.t25 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X135 vdd.t34 vbias.t91 vout.t81 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X136 w_20679_4119.t47 vp.t10 a_21819_2107.t5 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X137 vout.t24 a_21819_2107.t71 vss.t39 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X138 vss.t38 a_21819_2107.t72 vout.t23 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X139 vout.t22 a_21819_2107.t73 vss.t37 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X140 vss.t36 a_21819_2107.t74 vout.t21 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X141 w_20679_4119.t29 vbias.t92 vdd.t33 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X142 w_20679_4119.t6 vn.t7 a_20875_2019.t36 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X143 w_20679_4119.t7 vn.t8 a_20875_2019.t37 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X144 vdd.t32 vbias.t93 w_20679_4119.t28 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X145 vdd.t31 vbias.t94 w_20679_4119.t27 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X146 vout.t20 a_21819_2107.t75 vss.t35 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X147 vout.t80 vbias.t95 vdd.t30 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X148 vss.t34 a_21819_2107.t76 vout.t19 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X149 a_20875_2019.t18 a_20875_2019.t17 vss.t7 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X150 w_20679_4119.t26 vbias.t96 vdd.t29 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X151 vdd.t28 vbias.t97 w_20679_4119.t25 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X152 vdd.t27 vbias.t98 vout.t79 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X153 a_20875_2019.t16 a_20875_2019.t15 vss.t6 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X154 vss.t33 a_21819_2107.t77 vout.t18 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X155 vout.t78 vbias.t99 vdd.t26 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X156 vdd.t25 vbias.t100 vout.t77 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X157 vout.t76 vbias.t101 vdd.t24 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X158 w_20679_4119.t8 vn.t9 a_20875_2019.t38 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X159 a_20875_2019.t14 a_20875_2019.t13 vss.t5 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X160 vss.t32 a_21819_2107.t78 vout.t17 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X161 vss.t31 a_21819_2107.t79 vout.t16 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X162 a_21819_2107.t4 vp.t11 w_20679_4119.t48 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X163 a_20875_2019.t12 a_20875_2019.t11 vss.t4 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X164 vdd.t23 vbias.t10 vbias.t11 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X165 vdd.t22 vbias.t102 w_20679_4119.t24 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X166 a_20875_2019.t39 vn.t10 w_20679_4119.t9 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X167 vss.t30 a_21819_2107.t80 vout.t15 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X168 w_20679_4119.t23 vbias.t103 vdd.t21 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X169 vbias.t9 vbias.t8 vdd.t20 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X170 vdd.t19 vbias.t104 vout.t75 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X171 a_20875_2019.t40 vn.t11 w_20679_4119.t10 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X172 vss.t90 a_20875_2019.t58 a_21819_2107.t26 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X173 vdd.t18 vbias.t6 vbias.t7 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X174 vss.t29 a_21819_2107.t81 vout.t14 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X175 vdd.t17 vbias.t105 vout.t74 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X176 vout.t13 a_21819_2107.t82 vss.t28 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X177 vdd.t16 vbias.t106 w_20679_4119.t22 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X178 vdd.t15 vbias.t107 vout.t73 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X179 vout.t72 vbias.t108 vdd.t14 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X180 vss.t27 a_21819_2107.t83 vout.t12 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X181 vout.t11 a_21819_2107.t84 vss.t26 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X182 vss.t25 a_21819_2107.t85 vout.t10 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X183 vout.t9 a_21819_2107.t86 vss.t24 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X184 a_21819_2107.t3 vp.t12 w_20679_4119.t49 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X185 vss.t91 a_20875_2019.t59 a_21819_2107.t27 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X186 vbias.t5 vbias.t4 vdd.t13 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X187 vout.t71 vbias.t109 vdd.t12 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X188 vss.t23 a_21819_2107.t87 vout.t8 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X189 vdd.t11 vbias.t110 vout.t70 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X190 w_20679_4119.t21 vbias.t111 vdd.t10 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X191 w_20679_4119.t50 vp.t13 a_21819_2107.t2 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X192 vout.t7 a_21819_2107.t88 vss.t22 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X193 a_21819_2107.t28 a_20875_2019.t60 vss.t92 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X194 vout.t69 vbias.t112 vdd.t9 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X195 vss.t21 a_21819_2107.t89 vout.t6 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X196 vout.t68 vbias.t113 vdd.t8 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X197 vdd.t7 vbias.t114 vout.t67 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X198 vss.t3 a_20875_2019.t9 a_20875_2019.t10 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X199 vss.t2 a_20875_2019.t7 a_20875_2019.t8 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X200 a_20875_2019.t41 vn.t12 w_20679_4119.t11 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X201 a_21819_2107.t29 a_20875_2019.t61 vss.t93 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X202 vout.t5 a_21819_2107.t90 vss.t20 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X203 vout.t4 a_21819_2107.t91 vss.t19 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X204 vdd.t6 vbias.t115 w_20679_4119.t20 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X205 a_20875_2019.t42 vn.t13 w_20679_4119.t12 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X206 vss.t18 a_21819_2107.t92 vout.t3 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X207 vbias.t3 vbias.t2 vdd.t5 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X208 a_21819_2107.t1 vp.t14 w_20679_4119.t51 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X209 vdd.t4 vbias.t116 vout.t66 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X210 vss.t94 a_20875_2019.t62 a_21819_2107.t30 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X211 vout.t65 vbias.t117 vdd.t3 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X212 vdd.t2 vbias.t118 vout.t64 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X213 vss.t1 a_20875_2019.t5 a_20875_2019.t6 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X214 vout.t2 a_21819_2107.t93 vss.t17 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X215 vss.t0 a_20875_2019.t3 a_20875_2019.t4 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X216 vout.t1 a_21819_2107.t94 vss.t16 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X217 w_20679_4119.t19 vbias.t119 vdd.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X218 vout.t0 a_21819_2107.t95 vss.t15 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X219 a_20875_2019.t43 vn.t14 w_20679_4119.t13 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X220 a_20875_2019.t44 vn.t15 w_20679_4119.t14 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X221 w_20679_4119.t52 vp.t15 a_21819_2107.t0 w_20679_4119# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X222 vss.t95 a_20875_2019.t63 a_21819_2107.t31 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X223 vdd.t0 vbias.t0 vbias.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
C0 vn vp 1.91fF
C1 vdd vbias 34.89fF
C2 vdd vout 13.38fF
C3 vbias vout 9.42fF
R0 vbias.n128 vbias.t6 63.632
R1 vbias.n195 vbias.t30 63.63
R2 vbias.n87 vbias.t36 63.63
R3 vbias.n194 vbias.t103 63.63
R4 vbias.n19 vbias.t90 63.63
R5 vbias.n105 vbias.t109 63.63
R6 vbias.n105 vbias.t85 63.63
R7 vbias.n20 vbias.t110 63.63
R8 vbias.n106 vbias.t77 63.63
R9 vbias.n106 vbias.t55 63.63
R10 vbias.n18 vbias.t74 63.63
R11 vbias.n104 vbias.t65 63.63
R12 vbias.n104 vbias.t116 63.63
R13 vbias.n21 vbias.t54 63.63
R14 vbias.n107 vbias.t86 63.63
R15 vbias.n107 vbias.t64 63.63
R16 vbias.n23 vbias.t108 63.63
R17 vbias.n109 vbias.t78 63.63
R18 vbias.n109 vbias.t58 63.63
R19 vbias.n24 vbias.t59 63.63
R20 vbias.n110 vbias.t98 63.63
R21 vbias.n110 vbias.t75 63.63
R22 vbias.n22 vbias.t69 63.63
R23 vbias.n108 vbias.t57 63.63
R24 vbias.n108 vbias.t107 63.63
R25 vbias.n25 vbias.t101 63.63
R26 vbias.n111 vbias.t50 63.63
R27 vbias.n111 vbias.t99 63.63
R28 vbias.n27 vbias.t68 63.63
R29 vbias.n113 vbias.t112 63.63
R30 vbias.n113 vbias.t88 63.63
R31 vbias.n28 vbias.t105 63.63
R32 vbias.n114 vbias.t61 63.63
R33 vbias.n114 vbias.t114 63.63
R34 vbias.n26 vbias.t53 63.63
R35 vbias.n112 vbias.t67 63.63
R36 vbias.n112 vbias.t118 63.63
R37 vbias.n29 vbias.t82 63.63
R38 vbias.n115 vbias.t60 63.63
R39 vbias.n115 vbias.t113 63.63
R40 vbias.n31 vbias.t117 63.63
R41 vbias.n117 vbias.t72 63.63
R42 vbias.n117 vbias.t52 63.63
R43 vbias.n32 vbias.t91 63.63
R44 vbias.n118 vbias.t70 63.63
R45 vbias.n118 vbias.t51 63.63
R46 vbias.n30 vbias.t100 63.63
R47 vbias.n116 vbias.t104 63.63
R48 vbias.n116 vbias.t81 63.63
R49 vbias.n63 vbias.t66 63.63
R50 vbias.n126 vbias.t111 63.63
R51 vbias.n126 vbias.t87 63.63
R52 vbias.n159 vbias.t38 63.63
R53 vbias.n159 vbias.t28 63.63
R54 vbias.n77 vbias.t40 63.63
R55 vbias.n64 vbias.t12 63.63
R56 vbias.n103 vbias.t42 63.63
R57 vbias.n62 vbias.t97 63.63
R58 vbias.n125 vbias.t84 63.63
R59 vbias.n125 vbias.t63 63.63
R60 vbias.n33 vbias.t56 63.63
R61 vbias.n119 vbias.t95 63.63
R62 vbias.n119 vbias.t73 63.63
R63 vbias.n123 vbias.t14 63.63
R64 vbias.n35 vbias.t24 63.63
R65 vbias.n123 vbias.t2 63.63
R66 vbias.n78 vbias.t94 63.63
R67 vbias.n161 vbias.t102 63.63
R68 vbias.n161 vbias.t79 63.63
R69 vbias.n83 vbias.t76 63.63
R70 vbias.n188 vbias.t115 63.63
R71 vbias.n188 vbias.t89 63.63
R72 vbias.n189 vbias.t62 63.63
R73 vbias.n190 vbias.t26 63.63
R74 vbias.n192 vbias.t8 63.63
R75 vbias.n192 vbias.t44 63.63
R76 vbias.n85 vbias.t0 63.63
R77 vbias.n190 vbias.t10 63.63
R78 vbias.n163 vbias.t18 63.63
R79 vbias.n80 vbias.t34 63.63
R80 vbias.n82 vbias.t16 63.63
R81 vbias.n186 vbias.t4 63.63
R82 vbias.n163 vbias.t32 63.63
R83 vbias.n186 vbias.t22 63.63
R84 vbias.n79 vbias.t49 63.63
R85 vbias.n162 vbias.t48 63.63
R86 vbias.n162 vbias.t96 63.63
R87 vbias.n90 vbias.t106 63.63
R88 vbias.n193 vbias.t93 63.63
R89 vbias.n193 vbias.t71 63.63
R90 vbias.n194 vbias.t80 63.63
R91 vbias.n189 vbias.t83 63.63
R92 vbias.n84 vbias.t92 63.63
R93 vbias.n91 vbias.t20 63.63
R94 vbias.n89 vbias.t119 63.63
R95 vbias.n195 vbias.t46 63.63
R96 vbias.n0 vbias.t31 14.295
R97 vbias.n9 vbias.t37 14.295
R98 vbias.n156 vbias.t39 14.295
R99 vbias.n156 vbias.t7 14.295
R100 vbias.n132 vbias.t43 14.295
R101 vbias.n132 vbias.t29 14.295
R102 vbias.n74 vbias.t13 14.295
R103 vbias.n74 vbias.t41 14.295
R104 vbias.n134 vbias.t15 14.295
R105 vbias.n53 vbias.t25 14.295
R106 vbias.n56 vbias.t3 14.295
R107 vbias.n101 vbias.t9 14.295
R108 vbias.n101 vbias.t27 14.295
R109 vbias.n94 vbias.t11 14.295
R110 vbias.n94 vbias.t45 14.295
R111 vbias.n17 vbias.t1 14.295
R112 vbias.n17 vbias.t21 14.295
R113 vbias.n183 vbias.t33 14.295
R114 vbias.n183 vbias.t23 14.295
R115 vbias.n173 vbias.t19 14.295
R116 vbias.n173 vbias.t5 14.295
R117 vbias.n171 vbias.t17 14.295
R118 vbias.n171 vbias.t35 14.295
R119 vbias.n3 vbias.t47 14.295
R120 vbias.n196 vbias.n0 3.25
R121 vbias.n196 vbias.n3 1.139
R122 vbias.n3 vbias.n2 0.874
R123 vbias.n10 vbias.n9 0.87
R124 vbias.n53 vbias.n52 0.823
R125 vbias.n150 vbias.n134 0.823
R126 vbias.n54 vbias.n53 0.594
R127 vbias.n57 vbias.n56 0.58
R128 vbias.n13 vbias.n12 0.577
R129 vbias.n37 vbias.n36 0.575
R130 vbias.n38 vbias.n37 0.575
R131 vbias.n39 vbias.n38 0.575
R132 vbias.n41 vbias.n40 0.575
R133 vbias.n42 vbias.n41 0.575
R134 vbias.n40 vbias.n39 0.575
R135 vbias.n43 vbias.n42 0.575
R136 vbias.n45 vbias.n44 0.575
R137 vbias.n46 vbias.n45 0.575
R138 vbias.n44 vbias.n43 0.575
R139 vbias.n47 vbias.n46 0.575
R140 vbias.n49 vbias.n48 0.575
R141 vbias.n50 vbias.n49 0.575
R142 vbias.n48 vbias.n47 0.575
R143 vbias.n66 vbias.n65 0.575
R144 vbias.n152 vbias.n151 0.575
R145 vbias.n167 vbias.n166 0.575
R146 vbias.n5 vbias.n4 0.575
R147 vbias.n2 vbias.n1 0.575
R148 vbias.n138 vbias.n137 0.574
R149 vbias.n139 vbias.n138 0.574
R150 vbias.n142 vbias.n141 0.574
R151 vbias.n143 vbias.n142 0.574
R152 vbias.n146 vbias.n145 0.574
R153 vbias.n147 vbias.n146 0.574
R154 vbias.n67 vbias.n66 0.574
R155 vbias.n153 vbias.n152 0.574
R156 vbias.n96 vbias.n95 0.574
R157 vbias.n168 vbias.n167 0.574
R158 vbias.n175 vbias.n174 0.574
R159 vbias.n176 vbias.n175 0.574
R160 vbias.n12 vbias.n11 0.574
R161 vbias.n6 vbias.n5 0.574
R162 vbias.n11 vbias.n10 0.574
R163 vbias.n137 vbias.n136 0.574
R164 vbias.n141 vbias.n140 0.574
R165 vbias.n145 vbias.n144 0.574
R166 vbias.n149 vbias.n148 0.574
R167 vbias.n136 vbias.n135 0.573
R168 vbias.n140 vbias.n139 0.573
R169 vbias.n144 vbias.n143 0.573
R170 vbias.n148 vbias.n147 0.573
R171 vbias.n154 vbias.n153 0.573
R172 vbias.n98 vbias.n97 0.573
R173 vbias.n99 vbias.n98 0.573
R174 vbias.n52 vbias.n50 0.57
R175 vbias.n150 vbias.n149 0.569
R176 vbias.n73 vbias.n68 0.376
R177 vbias.n16 vbias.n7 0.376
R178 vbias.n182 vbias.n177 0.376
R179 vbias.n156 vbias.n155 0.337
R180 vbias.n171 vbias.n170 0.337
R181 vbias.n101 vbias.n100 0.332
R182 vbias.n188 vbias.n187 0.284
R183 vbias.n161 vbias.n160 0.284
R184 vbias.n125 vbias.n124 0.284
R185 vbias.n78 vbias.n77 0.281
R186 vbias.n193 vbias.n192 0.281
R187 vbias.n83 vbias.n82 0.281
R188 vbias.n20 vbias.n19 0.281
R189 vbias.n106 vbias.n105 0.281
R190 vbias.n21 vbias.n20 0.281
R191 vbias.n107 vbias.n106 0.281
R192 vbias.n19 vbias.n18 0.281
R193 vbias.n105 vbias.n104 0.281
R194 vbias.n22 vbias.n21 0.281
R195 vbias.n108 vbias.n107 0.281
R196 vbias.n24 vbias.n23 0.281
R197 vbias.n110 vbias.n109 0.281
R198 vbias.n25 vbias.n24 0.281
R199 vbias.n111 vbias.n110 0.281
R200 vbias.n23 vbias.n22 0.281
R201 vbias.n109 vbias.n108 0.281
R202 vbias.n26 vbias.n25 0.281
R203 vbias.n112 vbias.n111 0.281
R204 vbias.n28 vbias.n27 0.281
R205 vbias.n114 vbias.n113 0.281
R206 vbias.n29 vbias.n28 0.281
R207 vbias.n115 vbias.n114 0.281
R208 vbias.n27 vbias.n26 0.281
R209 vbias.n113 vbias.n112 0.281
R210 vbias.n30 vbias.n29 0.281
R211 vbias.n116 vbias.n115 0.281
R212 vbias.n32 vbias.n31 0.281
R213 vbias.n118 vbias.n117 0.281
R214 vbias.n33 vbias.n32 0.281
R215 vbias.n119 vbias.n118 0.281
R216 vbias.n31 vbias.n30 0.281
R217 vbias.n117 vbias.n116 0.281
R218 vbias.n63 vbias.n62 0.281
R219 vbias.n126 vbias.n125 0.281
R220 vbias.n79 vbias.n78 0.281
R221 vbias.n162 vbias.n161 0.281
R222 vbias.n84 vbias.n83 0.281
R223 vbias.n189 vbias.n188 0.281
R224 vbias.n91 vbias.n90 0.281
R225 vbias.n194 vbias.n193 0.281
R226 vbias.n85 vbias.n84 0.281
R227 vbias.n90 vbias.n89 0.281
R228 vbias.n64 vbias.n63 0.281
R229 vbias.n89 vbias.n88 0.281
R230 vbias.n62 vbias.n61 0.281
R231 vbias.n190 vbias.n189 0.28
R232 vbias.n163 vbias.n162 0.28
R233 vbias.n80 vbias.n79 0.28
R234 vbias.n195 vbias.n194 0.28
R235 vbias.n102 vbias.n94 0.234
R236 vbias.n94 vbias.n93 0.231
R237 vbias.n93 vbias.n17 0.231
R238 vbias.n74 vbias.n73 0.229
R239 vbias.n17 vbias.n16 0.229
R240 vbias.n183 vbias.n182 0.229
R241 vbias.n157 vbias.n132 0.227
R242 vbias.n75 vbias.n74 0.227
R243 vbias.n157 vbias.n156 0.227
R244 vbias.n102 vbias.n101 0.227
R245 vbias.n184 vbias.n173 0.227
R246 vbias.n173 vbias.n172 0.227
R247 vbias.n172 vbias.n171 0.227
R248 vbias.n184 vbias.n183 0.227
R249 vbias.n127 vbias.n126 0.217
R250 vbias.n34 vbias.n33 0.217
R251 vbias.n120 vbias.n119 0.217
R252 vbias.n131 vbias.n130 0.215
R253 vbias.n165 vbias.n164 0.215
R254 vbias.n73 vbias.n72 0.212
R255 vbias.n16 vbias.n15 0.212
R256 vbias.n182 vbias.n181 0.212
R257 vbias.n72 vbias.n71 0.175
R258 vbias.n15 vbias.n14 0.175
R259 vbias.n181 vbias.n180 0.175
R260 vbias.n155 vbias.n133 0.167
R261 vbias.n170 vbias.n169 0.167
R262 vbias.n155 vbias.n154 0.167
R263 vbias.n170 vbias.n168 0.167
R264 vbias.n100 vbias.n96 0.165
R265 vbias.n100 vbias.n99 0.164
R266 vbias.n179 vbias.n178 0.132
R267 vbias.n70 vbias.n69 0.132
R268 vbias.n13 vbias.n8 0.132
R269 vbias.n88 vbias.n86 0.09
R270 vbias.n196 vbias.n195 0.085
R271 vbias.n158 vbias.n157 0.081
R272 vbias.n185 vbias.n184 0.081
R273 vbias.n92 vbias.n91 0.074
R274 vbias.n192 vbias.n191 0.074
R275 vbias.n191 vbias.n190 0.074
R276 vbias.n92 vbias.n85 0.074
R277 vbias.n77 vbias.n76 0.073
R278 vbias.n82 vbias.n81 0.073
R279 vbias.n76 vbias.n64 0.073
R280 vbias.n81 vbias.n80 0.073
R281 vbias.n123 vbias.n122 0.068
R282 vbias.n159 vbias.n158 0.067
R283 vbias.n186 vbias.n185 0.067
R284 vbias.n124 vbias.n120 0.065
R285 vbias.n160 vbias.n131 0.065
R286 vbias.n187 vbias.n165 0.065
R287 vbias.n128 vbias.n127 0.064
R288 vbias.n55 vbias.n34 0.064
R289 vbias.n93 vbias.n92 0.039
R290 vbias.n191 vbias.n102 0.038
R291 vbias.n76 vbias.n75 0.038
R292 vbias vbias.n196 0.021
R293 vbias.n58 vbias.n57 0.014
R294 vbias.n177 vbias.n176 0.005
R295 vbias.n68 vbias.n67 0.005
R296 vbias.n7 vbias.n6 0.005
R297 vbias.n151 vbias.n150 0.005
R298 vbias.n52 vbias.n51 0.005
R299 vbias.n164 vbias.n163 0.002
R300 vbias.n130 vbias.n129 0.002
R301 vbias.n55 vbias.n54 0.001
R302 vbias.n59 vbias.n58 0.001
R303 vbias.n180 vbias.n179 0.001
R304 vbias.n129 vbias.n128 0.001
R305 vbias.n122 vbias.n121 0.001
R306 vbias.n61 vbias.n60 0.001
R307 vbias.n88 vbias.n87 0.001
R308 vbias.n129 vbias.n103 0.001
R309 vbias.n54 vbias.n35 0.001
R310 vbias.n160 vbias.n159 0.001
R311 vbias.n71 vbias.n70 0.001
R312 vbias.n124 vbias.n123 0.001
R313 vbias.n14 vbias.n13 0.001
R314 vbias.n187 vbias.n186 0.001
R315 vbias.n60 vbias.n59 0.001
R316 vbias.n59 vbias.n55 0.001
R317 vdd.n118 vdd.n117 386.601
R318 vdd.n103 vdd.n101 127.023
R319 vdd.n98 vdd.n96 127.023
R320 vdd.n87 vdd.n85 127.023
R321 vdd.n82 vdd.n80 127.023
R322 vdd.n71 vdd.n69 127.023
R323 vdd.n66 vdd.n64 127.023
R324 vdd.n45 vdd.n43 127.023
R325 vdd.n40 vdd.n38 127.023
R326 vdd.n29 vdd.n27 127.023
R327 vdd.n24 vdd.n22 127.023
R328 vdd.n13 vdd.n11 127.023
R329 vdd.n8 vdd.n4 127.023
R330 vdd.n8 vdd.n6 127.023
R331 vdd.n122 vdd.n120 116.986
R332 vdd.n57 vdd.t61 15.566
R333 vdd.n114 vdd.t4 15.351
R334 vdd.n144 vdd.t1 14.295
R335 vdd.n144 vdd.t74 14.295
R336 vdd.n143 vdd.t21 14.295
R337 vdd.n143 vdd.t65 14.295
R338 vdd.n142 vdd.t52 14.295
R339 vdd.n142 vdd.t92 14.295
R340 vdd.n2 vdd.t41 14.295
R341 vdd.n2 vdd.t16 14.295
R342 vdd.n1 vdd.t88 14.295
R343 vdd.n1 vdd.t32 14.295
R344 vdd.n0 vdd.t20 14.295
R345 vdd.n0 vdd.t63 14.295
R346 vdd.n16 vdd.t33 14.295
R347 vdd.n16 vdd.t0 14.295
R348 vdd.n15 vdd.t48 14.295
R349 vdd.n15 vdd.t23 14.295
R350 vdd.n14 vdd.t76 14.295
R351 vdd.n14 vdd.t55 14.295
R352 vdd.n20 vdd.t39 14.295
R353 vdd.n20 vdd.t58 14.295
R354 vdd.n19 vdd.t13 14.295
R355 vdd.n19 vdd.t6 14.295
R356 vdd.n18 vdd.t46 14.295
R357 vdd.n18 vdd.t38 14.295
R358 vdd.n32 vdd.t94 14.295
R359 vdd.n32 vdd.t72 14.295
R360 vdd.n31 vdd.t95 14.295
R361 vdd.n31 vdd.t40 14.295
R362 vdd.n30 vdd.t29 14.295
R363 vdd.n30 vdd.t68 14.295
R364 vdd.n36 vdd.t86 14.295
R365 vdd.n36 vdd.t31 14.295
R366 vdd.n35 vdd.t57 14.295
R367 vdd.n35 vdd.t22 14.295
R368 vdd.n34 vdd.t84 14.295
R369 vdd.n34 vdd.t53 14.295
R370 vdd.n48 vdd.t70 14.295
R371 vdd.n48 vdd.t35 14.295
R372 vdd.n47 vdd.t10 14.295
R373 vdd.n47 vdd.t87 14.295
R374 vdd.n46 vdd.t43 14.295
R375 vdd.n46 vdd.t18 14.295
R376 vdd.n52 vdd.t50 14.295
R377 vdd.n52 vdd.t28 14.295
R378 vdd.n51 vdd.t5 14.295
R379 vdd.n51 vdd.t47 14.295
R380 vdd.n50 vdd.t36 14.295
R381 vdd.n50 vdd.t75 14.295
R382 vdd.n58 vdd.t82 14.295
R383 vdd.n57 vdd.t30 14.295
R384 vdd.n62 vdd.t3 14.295
R385 vdd.n62 vdd.t34 14.295
R386 vdd.n61 vdd.t62 14.295
R387 vdd.n61 vdd.t64 14.295
R388 vdd.n60 vdd.t90 14.295
R389 vdd.n60 vdd.t91 14.295
R390 vdd.n74 vdd.t49 14.295
R391 vdd.n74 vdd.t25 14.295
R392 vdd.n73 vdd.t78 14.295
R393 vdd.n73 vdd.t19 14.295
R394 vdd.n72 vdd.t8 14.295
R395 vdd.n72 vdd.t51 14.295
R396 vdd.n78 vdd.t67 14.295
R397 vdd.n78 vdd.t17 14.295
R398 vdd.n77 vdd.t9 14.295
R399 vdd.n77 vdd.t77 14.295
R400 vdd.n76 vdd.t42 14.295
R401 vdd.n76 vdd.t7 14.295
R402 vdd.n90 vdd.t24 14.295
R403 vdd.n90 vdd.t89 14.295
R404 vdd.n89 vdd.t93 14.295
R405 vdd.n89 vdd.t69 14.295
R406 vdd.n88 vdd.t26 14.295
R407 vdd.n88 vdd.t2 14.295
R408 vdd.n94 vdd.t14 14.295
R409 vdd.n94 vdd.t79 14.295
R410 vdd.n93 vdd.t54 14.295
R411 vdd.n93 vdd.t27 14.295
R412 vdd.n92 vdd.t80 14.295
R413 vdd.n92 vdd.t59 14.295
R414 vdd.n106 vdd.t85 14.295
R415 vdd.n106 vdd.t66 14.295
R416 vdd.n105 vdd.t44 14.295
R417 vdd.n105 vdd.t81 14.295
R418 vdd.n104 vdd.t73 14.295
R419 vdd.n104 vdd.t15 14.295
R420 vdd.n110 vdd.t37 14.295
R421 vdd.n110 vdd.t11 14.295
R422 vdd.n109 vdd.t12 14.295
R423 vdd.n109 vdd.t56 14.295
R424 vdd.n108 vdd.t45 14.295
R425 vdd.n108 vdd.t83 14.295
R426 vdd.n115 vdd.t60 14.295
R427 vdd.n114 vdd.t71 14.295
R428 vdd.n58 vdd.n57 1.271
R429 vdd.n115 vdd.n114 1.056
R430 vdd.n143 vdd.n142 0.733
R431 vdd.n144 vdd.n143 0.733
R432 vdd.n1 vdd.n0 0.733
R433 vdd.n2 vdd.n1 0.733
R434 vdd.n15 vdd.n14 0.733
R435 vdd.n16 vdd.n15 0.733
R436 vdd.n19 vdd.n18 0.733
R437 vdd.n20 vdd.n19 0.733
R438 vdd.n31 vdd.n30 0.733
R439 vdd.n32 vdd.n31 0.733
R440 vdd.n35 vdd.n34 0.733
R441 vdd.n36 vdd.n35 0.733
R442 vdd.n47 vdd.n46 0.733
R443 vdd.n48 vdd.n47 0.733
R444 vdd.n51 vdd.n50 0.733
R445 vdd.n52 vdd.n51 0.733
R446 vdd.n61 vdd.n60 0.733
R447 vdd.n62 vdd.n61 0.733
R448 vdd.n73 vdd.n72 0.733
R449 vdd.n74 vdd.n73 0.733
R450 vdd.n77 vdd.n76 0.733
R451 vdd.n78 vdd.n77 0.733
R452 vdd.n89 vdd.n88 0.733
R453 vdd.n90 vdd.n89 0.733
R454 vdd.n93 vdd.n92 0.733
R455 vdd.n94 vdd.n93 0.733
R456 vdd.n105 vdd.n104 0.733
R457 vdd.n106 vdd.n105 0.733
R458 vdd.n109 vdd.n108 0.733
R459 vdd.n110 vdd.n109 0.733
R460 vdd.n59 vdd.n58 0.698
R461 vdd.n116 vdd.n115 0.586
R462 vdd.n145 vdd.n144 0.477
R463 vdd.n17 vdd.n16 0.477
R464 vdd.n33 vdd.n32 0.477
R465 vdd.n49 vdd.n48 0.477
R466 vdd.n75 vdd.n74 0.477
R467 vdd.n91 vdd.n90 0.477
R468 vdd.n107 vdd.n106 0.477
R469 vdd.n113 vdd.n110 0.477
R470 vdd.n99 vdd.n94 0.477
R471 vdd.n83 vdd.n78 0.477
R472 vdd.n67 vdd.n62 0.477
R473 vdd.n55 vdd.n52 0.477
R474 vdd.n41 vdd.n36 0.477
R475 vdd.n25 vdd.n20 0.477
R476 vdd.n9 vdd.n2 0.477
R477 vdd.n133 vdd.n55 0.378
R478 vdd vdd.n145 0.296
R479 vdd.n132 vdd.n59 0.286
R480 vdd.n139 vdd.n9 0.274
R481 vdd.n137 vdd.n25 0.274
R482 vdd.n135 vdd.n41 0.274
R483 vdd.n131 vdd.n67 0.274
R484 vdd.n129 vdd.n83 0.274
R485 vdd.n127 vdd.n99 0.274
R486 vdd.n125 vdd.n113 0.274
R487 vdd.n126 vdd.n107 0.274
R488 vdd.n128 vdd.n91 0.274
R489 vdd.n130 vdd.n75 0.274
R490 vdd.n134 vdd.n49 0.274
R491 vdd.n136 vdd.n33 0.274
R492 vdd.n138 vdd.n17 0.274
R493 vdd.n125 vdd.n124 0.261
R494 vdd.n123 vdd.n122 0.212
R495 vdd.n122 vdd.n121 0.212
R496 vdd.n112 vdd.n111 0.195
R497 vdd.n103 vdd.n102 0.195
R498 vdd.n98 vdd.n97 0.195
R499 vdd.n87 vdd.n86 0.195
R500 vdd.n82 vdd.n81 0.195
R501 vdd.n71 vdd.n70 0.195
R502 vdd.n45 vdd.n44 0.195
R503 vdd.n40 vdd.n39 0.195
R504 vdd.n29 vdd.n28 0.195
R505 vdd.n24 vdd.n23 0.195
R506 vdd.n13 vdd.n12 0.195
R507 vdd.n8 vdd.n7 0.195
R508 vdd.n126 vdd.n125 0.034
R509 vdd.n127 vdd.n126 0.034
R510 vdd.n128 vdd.n127 0.034
R511 vdd.n129 vdd.n128 0.034
R512 vdd.n130 vdd.n129 0.034
R513 vdd.n131 vdd.n130 0.034
R514 vdd.n132 vdd.n131 0.034
R515 vdd.n134 vdd.n133 0.034
R516 vdd.n135 vdd.n134 0.034
R517 vdd.n136 vdd.n135 0.034
R518 vdd.n137 vdd.n136 0.034
R519 vdd.n138 vdd.n137 0.034
R520 vdd.n139 vdd.n138 0.034
R521 vdd.n124 vdd.n123 0.027
R522 vdd.n66 vdd.n65 0.018
R523 vdd.n133 vdd.n132 0.017
R524 vdd.n141 vdd.n140 0.017
R525 vdd.n54 vdd.n53 0.017
R526 vdd vdd.n139 0.011
R527 vdd.n123 vdd.n118 0.001
R528 vdd.n120 vdd.n119 0.001
R529 vdd.n101 vdd.n100 0.001
R530 vdd.n96 vdd.n95 0.001
R531 vdd.n85 vdd.n84 0.001
R532 vdd.n80 vdd.n79 0.001
R533 vdd.n69 vdd.n68 0.001
R534 vdd.n64 vdd.n63 0.001
R535 vdd.n43 vdd.n42 0.001
R536 vdd.n38 vdd.n37 0.001
R537 vdd.n27 vdd.n26 0.001
R538 vdd.n22 vdd.n21 0.001
R539 vdd.n11 vdd.n10 0.001
R540 vdd.n4 vdd.n3 0.001
R541 vdd.n6 vdd.n5 0.001
R542 vdd.n59 vdd.n56 0.001
R543 vdd.n113 vdd.n112 0.001
R544 vdd.n107 vdd.n103 0.001
R545 vdd.n99 vdd.n98 0.001
R546 vdd.n91 vdd.n87 0.001
R547 vdd.n83 vdd.n82 0.001
R548 vdd.n75 vdd.n71 0.001
R549 vdd.n67 vdd.n66 0.001
R550 vdd.n55 vdd.n54 0.001
R551 vdd.n49 vdd.n45 0.001
R552 vdd.n41 vdd.n40 0.001
R553 vdd.n33 vdd.n29 0.001
R554 vdd.n25 vdd.n24 0.001
R555 vdd.n17 vdd.n13 0.001
R556 vdd.n9 vdd.n8 0.001
R557 vdd.n145 vdd.n141 0.001
R558 vdd.n118 vdd.n116 0.001
R559 w_20679_4119.n27 w_20679_4119.n26 779.876
R560 w_20679_4119.n49 w_20679_4119.t24 14.295
R561 w_20679_4119.n3 w_20679_4119.t41 14.295
R562 w_20679_4119.n3 w_20679_4119.t27 14.295
R563 w_20679_4119.n48 w_20679_4119.t26 14.295
R564 w_20679_4119.n48 w_20679_4119.t35 14.295
R565 w_20679_4119.n11 w_20679_4119.t31 14.295
R566 w_20679_4119.n11 w_20679_4119.t39 14.295
R567 w_20679_4119.n10 w_20679_4119.t21 14.295
R568 w_20679_4119.n10 w_20679_4119.t32 14.295
R569 w_20679_4119.n9 w_20679_4119.t38 14.295
R570 w_20679_4119.n9 w_20679_4119.t25 14.295
R571 w_20679_4119.n35 w_20679_4119.t37 14.295
R572 w_20679_4119.n35 w_20679_4119.t34 14.295
R573 w_20679_4119.n34 w_20679_4119.t28 14.295
R574 w_20679_4119.n34 w_20679_4119.t23 14.295
R575 w_20679_4119.n33 w_20679_4119.t19 14.295
R576 w_20679_4119.n33 w_20679_4119.t22 14.295
R577 w_20679_4119.n20 w_20679_4119.t40 14.295
R578 w_20679_4119.n20 w_20679_4119.t30 14.295
R579 w_20679_4119.n19 w_20679_4119.t33 14.295
R580 w_20679_4119.n19 w_20679_4119.t20 14.295
R581 w_20679_4119.n18 w_20679_4119.t29 14.295
R582 w_20679_4119.n18 w_20679_4119.t36 14.295
R583 w_20679_4119.t42 w_20679_4119.n49 14.295
R584 w_20679_4119.n28 w_20679_4119.t54 8.834
R585 w_20679_4119.n12 w_20679_4119.t55 8.766
R586 w_20679_4119.n14 w_20679_4119.t6 7.146
R587 w_20679_4119.n13 w_20679_4119.t5 7.146
R588 w_20679_4119.n12 w_20679_4119.t2 7.146
R589 w_20679_4119.n30 w_20679_4119.t13 7.146
R590 w_20679_4119.n29 w_20679_4119.t11 7.146
R591 w_20679_4119.n28 w_20679_4119.t9 7.146
R592 w_20679_4119.n25 w_20679_4119.t4 7.146
R593 w_20679_4119.n25 w_20679_4119.t8 7.146
R594 w_20679_4119.n24 w_20679_4119.t17 7.146
R595 w_20679_4119.n24 w_20679_4119.t7 7.146
R596 w_20679_4119.n23 w_20679_4119.t51 7.146
R597 w_20679_4119.n23 w_20679_4119.t0 7.146
R598 w_20679_4119.n22 w_20679_4119.t45 7.146
R599 w_20679_4119.n22 w_20679_4119.t53 7.146
R600 w_20679_4119.n43 w_20679_4119.t49 7.146
R601 w_20679_4119.n43 w_20679_4119.t16 7.146
R602 w_20679_4119.n42 w_20679_4119.t48 7.146
R603 w_20679_4119.n42 w_20679_4119.t52 7.146
R604 w_20679_4119.n41 w_20679_4119.t46 7.146
R605 w_20679_4119.n41 w_20679_4119.t50 7.146
R606 w_20679_4119.n40 w_20679_4119.t15 7.146
R607 w_20679_4119.n40 w_20679_4119.t44 7.146
R608 w_20679_4119.n8 w_20679_4119.t14 7.146
R609 w_20679_4119.n8 w_20679_4119.t43 7.146
R610 w_20679_4119.n7 w_20679_4119.t12 7.146
R611 w_20679_4119.n7 w_20679_4119.t3 7.146
R612 w_20679_4119.n6 w_20679_4119.t10 7.146
R613 w_20679_4119.n6 w_20679_4119.t18 7.146
R614 w_20679_4119.n5 w_20679_4119.t1 7.146
R615 w_20679_4119.n5 w_20679_4119.t47 7.146
R616 w_20679_4119.n0 w_20679_4119.n27 5.228
R617 w_20679_4119.n15 w_20679_4119.n11 2.373
R618 w_20679_4119.n36 w_20679_4119.n35 2.373
R619 w_20679_4119.n29 w_20679_4119.n28 1.688
R620 w_20679_4119.n30 w_20679_4119.n29 1.688
R621 w_20679_4119.n13 w_20679_4119.n12 1.62
R622 w_20679_4119.n14 w_20679_4119.n13 1.62
R623 w_20679_4119.n15 w_20679_4119.n14 1.149
R624 w_20679_4119.n23 w_20679_4119.n22 1.045
R625 w_20679_4119.n24 w_20679_4119.n23 1.045
R626 w_20679_4119.n25 w_20679_4119.n24 1.045
R627 w_20679_4119.n41 w_20679_4119.n40 1.045
R628 w_20679_4119.n42 w_20679_4119.n41 1.045
R629 w_20679_4119.n43 w_20679_4119.n42 1.045
R630 w_20679_4119.n6 w_20679_4119.n5 1.045
R631 w_20679_4119.n7 w_20679_4119.n6 1.045
R632 w_20679_4119.n8 w_20679_4119.n7 1.045
R633 w_20679_4119.n39 w_20679_4119.n20 0.893
R634 w_20679_4119.n48 w_20679_4119.n47 0.893
R635 w_20679_4119.n44 w_20679_4119.n43 0.888
R636 w_20679_4119.n0 w_20679_4119.n30 0.871
R637 w_20679_4119.n44 w_20679_4119.n39 1.316
R638 w_20679_4119.n46 w_20679_4119.n44 0.748
R639 w_20679_4119.n47 w_20679_4119.n17 0.748
R640 w_20679_4119.n49 w_20679_4119.n3 0.733
R641 w_20679_4119.n10 w_20679_4119.n9 0.733
R642 w_20679_4119.n11 w_20679_4119.n10 0.733
R643 w_20679_4119.n34 w_20679_4119.n33 0.733
R644 w_20679_4119.n35 w_20679_4119.n34 0.733
R645 w_20679_4119.n19 w_20679_4119.n18 0.733
R646 w_20679_4119.n20 w_20679_4119.n19 0.733
R647 w_20679_4119.n49 w_20679_4119.n48 0.733
R648 w_20679_4119.n38 w_20679_4119.n36 0.72
R649 w_20679_4119.n2 w_20679_4119.n25 0.621
R650 w_20679_4119.n1 w_20679_4119.n8 0.621
R651 w_20679_4119.n39 w_20679_4119.n38 0.568
R652 w_20679_4119.n47 w_20679_4119.n46 0.568
R653 w_20679_4119.n17 w_20679_4119.n15 0.541
R654 w_20679_4119.n17 w_20679_4119.n16 0.491
R655 w_20679_4119.n46 w_20679_4119.n45 0.491
R656 w_20679_4119.n38 w_20679_4119.n37 0.491
R657 w_20679_4119.n36 w_20679_4119.n0 0.288
R658 w_20679_4119.n0 w_20679_4119.n32 0.28
R659 w_20679_4119.n32 w_20679_4119.n31 0.28
R660 w_20679_4119.n47 w_20679_4119.n1 0.267
R661 w_20679_4119.n39 w_20679_4119.n2 0.267
R662 w_20679_4119.n2 w_20679_4119.n21 0.196
R663 w_20679_4119.n1 w_20679_4119.n4 0.196
R664 vp.n0 vp.t10 111.996
R665 vp.n25 vp.t8 111.994
R666 vp.n6 vp.t12 111.83
R667 vp.n10 vp.t11 111.83
R668 vp.n21 vp.t9 111.83
R669 vp.n1 vp.t5 111.83
R670 vp.n15 vp.t6 111.83
R671 vp.n17 vp.t4 111.83
R672 vp.n19 vp.t0 111.83
R673 vp.n8 vp.t3 111.83
R674 vp.n12 vp.t2 111.83
R675 vp.n23 vp.t14 111.83
R676 vp.n2 vp.t7 111.83
R677 vp.n22 vp.t13 111.83
R678 vp.n11 vp.t15 111.83
R679 vp.n7 vp.t1 111.83
R680 vp.n25 vp.n24 2.022
R681 vp.n18 vp.n16 2.018
R682 vp.n13 vp.n9 2.018
R683 vp.n24 vp.n13 2.018
R684 vp.n20 vp.n18 2.018
R685 vp.n9 vp.n5 1.986
R686 vp.n16 vp.n14 1.986
R687 vp vp.n26 1.714
R688 vp.n26 vp.n0 0.868
R689 vp.n2 vp.n1 0.619
R690 vp.n4 vp.n3 0.547
R691 vp.n7 vp.n6 0.281
R692 vp.n11 vp.n10 0.281
R693 vp.n22 vp.n21 0.281
R694 vp.n5 vp.n4 0.273
R695 vp.n25 vp.n2 0.167
R696 vp.n21 vp.n20 0.14
R697 vp.n24 vp.n23 0.14
R698 vp.n13 vp.n12 0.14
R699 vp.n9 vp.n8 0.14
R700 vp.n16 vp.n15 0.139
R701 vp.n18 vp.n17 0.139
R702 vp.n20 vp.n19 0.139
R703 vp.n24 vp.n22 0.139
R704 vp.n13 vp.n11 0.139
R705 vp.n9 vp.n7 0.139
R706 vp.n26 vp.n25 0.136
R707 a_21819_2107.n55 a_21819_2107.t60 37.361
R708 a_21819_2107.n40 a_21819_2107.t90 37.361
R709 a_21819_2107.n25 a_21819_2107.t57 37.361
R710 a_21819_2107.n56 a_21819_2107.t76 37.361
R711 a_21819_2107.n41 a_21819_2107.t42 37.361
R712 a_21819_2107.n26 a_21819_2107.t70 37.361
R713 a_21819_2107.n57 a_21819_2107.t32 37.361
R714 a_21819_2107.n42 a_21819_2107.t63 37.361
R715 a_21819_2107.n27 a_21819_2107.t93 37.361
R716 a_21819_2107.n58 a_21819_2107.t48 37.361
R717 a_21819_2107.n43 a_21819_2107.t78 37.361
R718 a_21819_2107.n28 a_21819_2107.t45 37.361
R719 a_21819_2107.n59 a_21819_2107.t88 37.361
R720 a_21819_2107.n44 a_21819_2107.t53 37.361
R721 a_21819_2107.n29 a_21819_2107.t82 37.361
R722 a_21819_2107.n60 a_21819_2107.t44 37.361
R723 a_21819_2107.n45 a_21819_2107.t72 37.361
R724 a_21819_2107.n30 a_21819_2107.t38 37.361
R725 a_21819_2107.n61 a_21819_2107.t43 37.361
R726 a_21819_2107.n46 a_21819_2107.t73 37.361
R727 a_21819_2107.n31 a_21819_2107.t37 37.361
R728 a_21819_2107.n62 a_21819_2107.t80 37.361
R729 a_21819_2107.n47 a_21819_2107.t47 37.361
R730 a_21819_2107.n32 a_21819_2107.t77 37.361
R731 a_21819_2107.n63 a_21819_2107.t55 37.361
R732 a_21819_2107.n48 a_21819_2107.t86 37.361
R733 a_21819_2107.n33 a_21819_2107.t49 37.361
R734 a_21819_2107.n64 a_21819_2107.t56 37.361
R735 a_21819_2107.n49 a_21819_2107.t83 37.361
R736 a_21819_2107.n34 a_21819_2107.t50 37.361
R737 a_21819_2107.n65 a_21819_2107.t75 37.361
R738 a_21819_2107.n50 a_21819_2107.t39 37.361
R739 a_21819_2107.n35 a_21819_2107.t69 37.361
R740 a_21819_2107.n66 a_21819_2107.t92 37.361
R741 a_21819_2107.n51 a_21819_2107.t59 37.361
R742 a_21819_2107.n36 a_21819_2107.t89 37.361
R743 a_21819_2107.n67 a_21819_2107.t64 37.361
R744 a_21819_2107.n52 a_21819_2107.t95 37.361
R745 a_21819_2107.n37 a_21819_2107.t61 37.361
R746 a_21819_2107.n68 a_21819_2107.t87 37.361
R747 a_21819_2107.n53 a_21819_2107.t52 37.361
R748 a_21819_2107.n38 a_21819_2107.t81 37.361
R749 a_21819_2107.n0 a_21819_2107.t35 37.361
R750 a_21819_2107.n1 a_21819_2107.t65 37.361
R751 a_21819_2107.n2 a_21819_2107.t33 37.361
R752 a_21819_2107.n23 a_21819_2107.t66 37.361
R753 a_21819_2107.n24 a_21819_2107.t68 37.361
R754 a_21819_2107.n37 a_21819_2107.t94 37.361
R755 a_21819_2107.n38 a_21819_2107.t51 37.361
R756 a_21819_2107.n34 a_21819_2107.t85 37.361
R757 a_21819_2107.n35 a_21819_2107.t40 37.361
R758 a_21819_2107.n31 a_21819_2107.t71 37.361
R759 a_21819_2107.n32 a_21819_2107.t46 37.361
R760 a_21819_2107.n28 a_21819_2107.t79 37.361
R761 a_21819_2107.n29 a_21819_2107.t54 37.361
R762 a_21819_2107.n25 a_21819_2107.t91 37.361
R763 a_21819_2107.n26 a_21819_2107.t41 37.361
R764 a_21819_2107.n27 a_21819_2107.t62 37.361
R765 a_21819_2107.n30 a_21819_2107.t74 37.361
R766 a_21819_2107.n33 a_21819_2107.t84 37.361
R767 a_21819_2107.n36 a_21819_2107.t58 37.361
R768 a_21819_2107.n24 a_21819_2107.t34 37.361
R769 a_21819_2107.n39 a_21819_2107.t67 37.361
R770 a_21819_2107.n54 a_21819_2107.t36 37.361
R771 a_21819_2107.n8 a_21819_2107.t22 17.43
R772 a_21819_2107.n8 a_21819_2107.t16 17.43
R773 a_21819_2107.n7 a_21819_2107.t30 17.43
R774 a_21819_2107.n7 a_21819_2107.t24 17.43
R775 a_21819_2107.n6 a_21819_2107.t23 17.43
R776 a_21819_2107.n6 a_21819_2107.t17 17.43
R777 a_21819_2107.n5 a_21819_2107.t31 17.43
R778 a_21819_2107.n5 a_21819_2107.t25 17.43
R779 a_21819_2107.n92 a_21819_2107.t19 17.43
R780 a_21819_2107.n92 a_21819_2107.t20 17.43
R781 a_21819_2107.n91 a_21819_2107.t26 17.43
R782 a_21819_2107.n91 a_21819_2107.t28 17.43
R783 a_21819_2107.n90 a_21819_2107.t18 17.43
R784 a_21819_2107.n90 a_21819_2107.t21 17.43
R785 a_21819_2107.n89 a_21819_2107.t27 17.43
R786 a_21819_2107.n89 a_21819_2107.t29 17.43
R787 a_21819_2107.n97 a_21819_2107.t6 7.146
R788 a_21819_2107.n4 a_21819_2107.t4 7.146
R789 a_21819_2107.n4 a_21819_2107.t11 7.146
R790 a_21819_2107.n3 a_21819_2107.t3 7.146
R791 a_21819_2107.n3 a_21819_2107.t9 7.146
R792 a_21819_2107.n96 a_21819_2107.t10 7.146
R793 a_21819_2107.n96 a_21819_2107.t5 7.146
R794 a_21819_2107.n88 a_21819_2107.t8 7.146
R795 a_21819_2107.n88 a_21819_2107.t7 7.146
R796 a_21819_2107.n87 a_21819_2107.t2 7.146
R797 a_21819_2107.n87 a_21819_2107.t1 7.146
R798 a_21819_2107.n86 a_21819_2107.t0 7.146
R799 a_21819_2107.n86 a_21819_2107.t13 7.146
R800 a_21819_2107.n85 a_21819_2107.t12 7.146
R801 a_21819_2107.n85 a_21819_2107.t14 7.146
R802 a_21819_2107.t15 a_21819_2107.n97 7.146
R803 a_21819_2107.n94 a_21819_2107.n84 1.097
R804 a_21819_2107.n4 a_21819_2107.n3 1.045
R805 a_21819_2107.n97 a_21819_2107.n4 1.045
R806 a_21819_2107.n86 a_21819_2107.n85 1.045
R807 a_21819_2107.n87 a_21819_2107.n86 1.045
R808 a_21819_2107.n88 a_21819_2107.n87 1.045
R809 a_21819_2107.n97 a_21819_2107.n96 1.045
R810 a_21819_2107.n93 a_21819_2107.n88 0.983
R811 a_21819_2107.n96 a_21819_2107.n95 0.983
R812 a_21819_2107.n70 a_21819_2107.n69 0.604
R813 a_21819_2107.n10 a_21819_2107.n9 0.604
R814 a_21819_2107.n71 a_21819_2107.n70 0.604
R815 a_21819_2107.n72 a_21819_2107.n71 0.604
R816 a_21819_2107.n11 a_21819_2107.n10 0.604
R817 a_21819_2107.n12 a_21819_2107.n11 0.604
R818 a_21819_2107.n73 a_21819_2107.n72 0.604
R819 a_21819_2107.n13 a_21819_2107.n12 0.604
R820 a_21819_2107.n74 a_21819_2107.n73 0.604
R821 a_21819_2107.n75 a_21819_2107.n74 0.604
R822 a_21819_2107.n14 a_21819_2107.n13 0.604
R823 a_21819_2107.n15 a_21819_2107.n14 0.604
R824 a_21819_2107.n76 a_21819_2107.n75 0.604
R825 a_21819_2107.n16 a_21819_2107.n15 0.604
R826 a_21819_2107.n77 a_21819_2107.n76 0.604
R827 a_21819_2107.n78 a_21819_2107.n77 0.604
R828 a_21819_2107.n17 a_21819_2107.n16 0.604
R829 a_21819_2107.n18 a_21819_2107.n17 0.604
R830 a_21819_2107.n79 a_21819_2107.n78 0.604
R831 a_21819_2107.n19 a_21819_2107.n18 0.604
R832 a_21819_2107.n80 a_21819_2107.n79 0.604
R833 a_21819_2107.n81 a_21819_2107.n80 0.604
R834 a_21819_2107.n20 a_21819_2107.n19 0.604
R835 a_21819_2107.n21 a_21819_2107.n20 0.604
R836 a_21819_2107.n82 a_21819_2107.n81 0.604
R837 a_21819_2107.n83 a_21819_2107.n82 0.604
R838 a_21819_2107.n22 a_21819_2107.n21 0.604
R839 a_21819_2107.n23 a_21819_2107.n22 0.604
R840 a_21819_2107.n6 a_21819_2107.n5 0.545
R841 a_21819_2107.n7 a_21819_2107.n6 0.545
R842 a_21819_2107.n8 a_21819_2107.n7 0.545
R843 a_21819_2107.n90 a_21819_2107.n89 0.545
R844 a_21819_2107.n91 a_21819_2107.n90 0.545
R845 a_21819_2107.n92 a_21819_2107.n91 0.545
R846 a_21819_2107.n0 a_21819_2107.n83 0.523
R847 a_21819_2107.n95 a_21819_2107.n8 0.472
R848 a_21819_2107.n93 a_21819_2107.n92 0.472
R849 a_21819_2107.n2 a_21819_2107.n1 0.414
R850 a_21819_2107.n1 a_21819_2107.n0 0.414
R851 a_21819_2107.n84 a_21819_2107.n2 0.361
R852 a_21819_2107.n2 a_21819_2107.n38 0.356
R853 a_21819_2107.n1 a_21819_2107.n53 0.356
R854 a_21819_2107.n0 a_21819_2107.n68 0.356
R855 a_21819_2107.n56 a_21819_2107.n55 0.281
R856 a_21819_2107.n41 a_21819_2107.n40 0.281
R857 a_21819_2107.n42 a_21819_2107.n41 0.281
R858 a_21819_2107.n26 a_21819_2107.n25 0.281
R859 a_21819_2107.n57 a_21819_2107.n56 0.281
R860 a_21819_2107.n58 a_21819_2107.n57 0.281
R861 a_21819_2107.n43 a_21819_2107.n42 0.281
R862 a_21819_2107.n27 a_21819_2107.n26 0.281
R863 a_21819_2107.n28 a_21819_2107.n27 0.281
R864 a_21819_2107.n59 a_21819_2107.n58 0.281
R865 a_21819_2107.n44 a_21819_2107.n43 0.281
R866 a_21819_2107.n45 a_21819_2107.n44 0.281
R867 a_21819_2107.n29 a_21819_2107.n28 0.281
R868 a_21819_2107.n60 a_21819_2107.n59 0.281
R869 a_21819_2107.n61 a_21819_2107.n60 0.281
R870 a_21819_2107.n46 a_21819_2107.n45 0.281
R871 a_21819_2107.n30 a_21819_2107.n29 0.281
R872 a_21819_2107.n31 a_21819_2107.n30 0.281
R873 a_21819_2107.n62 a_21819_2107.n61 0.281
R874 a_21819_2107.n47 a_21819_2107.n46 0.281
R875 a_21819_2107.n48 a_21819_2107.n47 0.281
R876 a_21819_2107.n32 a_21819_2107.n31 0.281
R877 a_21819_2107.n63 a_21819_2107.n62 0.281
R878 a_21819_2107.n64 a_21819_2107.n63 0.281
R879 a_21819_2107.n49 a_21819_2107.n48 0.281
R880 a_21819_2107.n33 a_21819_2107.n32 0.281
R881 a_21819_2107.n34 a_21819_2107.n33 0.281
R882 a_21819_2107.n65 a_21819_2107.n64 0.281
R883 a_21819_2107.n50 a_21819_2107.n49 0.281
R884 a_21819_2107.n51 a_21819_2107.n50 0.281
R885 a_21819_2107.n35 a_21819_2107.n34 0.281
R886 a_21819_2107.n66 a_21819_2107.n65 0.281
R887 a_21819_2107.n67 a_21819_2107.n66 0.281
R888 a_21819_2107.n52 a_21819_2107.n51 0.281
R889 a_21819_2107.n36 a_21819_2107.n35 0.281
R890 a_21819_2107.n37 a_21819_2107.n36 0.281
R891 a_21819_2107.n68 a_21819_2107.n67 0.281
R892 a_21819_2107.n53 a_21819_2107.n52 0.281
R893 a_21819_2107.n38 a_21819_2107.n37 0.281
R894 a_21819_2107.n25 a_21819_2107.n24 0.281
R895 a_21819_2107.n40 a_21819_2107.n39 0.281
R896 a_21819_2107.n55 a_21819_2107.n54 0.281
R897 a_21819_2107.n95 a_21819_2107.n94 0.258
R898 a_21819_2107.n94 a_21819_2107.n93 0.258
R899 a_21819_2107.n84 a_21819_2107.n23 0.162
R900 vss.n87 vss.n85 127.023
R901 vss.n78 vss.n76 127.023
R902 vss.n69 vss.n67 127.023
R903 vss.n60 vss.n58 127.023
R904 vss.n38 vss.n36 127.023
R905 vss.n29 vss.n27 127.023
R906 vss.n20 vss.n18 127.023
R907 vss.n11 vss.n9 127.023
R908 vss.n6 vss.n4 113.388
R909 vss.n106 vss.n104 112.311
R910 vss.n0 vss.t79 18.06
R911 vss.n100 vss.t42 18.06
R912 vss.n2 vss.t5 17.43
R913 vss.n1 vss.t14 17.43
R914 vss.n0 vss.t7 17.43
R915 vss.n15 vss.t8 17.43
R916 vss.n15 vss.t93 17.43
R917 vss.n14 vss.t1 17.43
R918 vss.n14 vss.t85 17.43
R919 vss.n13 vss.t9 17.43
R920 vss.n13 vss.t92 17.43
R921 vss.n12 vss.t0 17.43
R922 vss.n12 vss.t84 17.43
R923 vss.n24 vss.t91 17.43
R924 vss.n24 vss.t89 17.43
R925 vss.n23 vss.t82 17.43
R926 vss.n23 vss.t81 17.43
R927 vss.n22 vss.t90 17.43
R928 vss.n22 vss.t88 17.43
R929 vss.n21 vss.t83 17.43
R930 vss.n21 vss.t80 17.43
R931 vss.n33 vss.t95 17.43
R932 vss.n33 vss.t4 17.43
R933 vss.n32 vss.t87 17.43
R934 vss.n32 vss.t13 17.43
R935 vss.n31 vss.t94 17.43
R936 vss.n31 vss.t6 17.43
R937 vss.n30 vss.t86 17.43
R938 vss.n30 vss.t12 17.43
R939 vss.n42 vss.t10 17.43
R940 vss.n42 vss.t75 17.43
R941 vss.n41 vss.t3 17.43
R942 vss.n41 vss.t45 17.43
R943 vss.n40 vss.t11 17.43
R944 vss.n40 vss.t77 17.43
R945 vss.n39 vss.t2 17.43
R946 vss.n39 vss.t44 17.43
R947 vss.n49 vss.t23 17.43
R948 vss.n49 vss.t46 17.43
R949 vss.n48 vss.t58 17.43
R950 vss.n48 vss.t15 17.43
R951 vss.n47 vss.t29 17.43
R952 vss.n47 vss.t49 17.43
R953 vss.n46 vss.t59 17.43
R954 vss.n46 vss.t16 17.43
R955 vss.n55 vss.t18 17.43
R956 vss.n55 vss.t35 17.43
R957 vss.n54 vss.t51 17.43
R958 vss.n54 vss.t71 17.43
R959 vss.n53 vss.t21 17.43
R960 vss.n53 vss.t41 17.43
R961 vss.n52 vss.t52 17.43
R962 vss.n52 vss.t70 17.43
R963 vss.n64 vss.t54 17.43
R964 vss.n64 vss.t55 17.43
R965 vss.n63 vss.t27 17.43
R966 vss.n63 vss.t24 17.43
R967 vss.n62 vss.t60 17.43
R968 vss.n62 vss.t61 17.43
R969 vss.n61 vss.t25 17.43
R970 vss.n61 vss.t26 17.43
R971 vss.n73 vss.t30 17.43
R972 vss.n73 vss.t67 17.43
R973 vss.n72 vss.t63 17.43
R974 vss.n72 vss.t37 17.43
R975 vss.n71 vss.t33 17.43
R976 vss.n71 vss.t73 17.43
R977 vss.n70 vss.t64 17.43
R978 vss.n70 vss.t39 17.43
R979 vss.n82 vss.t66 17.43
R980 vss.n82 vss.t22 17.43
R981 vss.n81 vss.t38 17.43
R982 vss.n81 vss.t57 17.43
R983 vss.n80 vss.t72 17.43
R984 vss.n80 vss.t28 17.43
R985 vss.n79 vss.t36 17.43
R986 vss.n79 vss.t56 17.43
R987 vss.n91 vss.t62 17.43
R988 vss.n91 vss.t78 17.43
R989 vss.n90 vss.t32 17.43
R990 vss.n90 vss.t47 17.43
R991 vss.n89 vss.t65 17.43
R992 vss.n89 vss.t17 17.43
R993 vss.n88 vss.t31 17.43
R994 vss.n88 vss.t48 17.43
R995 vss.n98 vss.t34 17.43
R996 vss.n98 vss.t50 17.43
R997 vss.n97 vss.t68 17.43
R998 vss.n97 vss.t20 17.43
R999 vss.n96 vss.t40 17.43
R1000 vss.n96 vss.t53 17.43
R1001 vss.n95 vss.t69 17.43
R1002 vss.n95 vss.t19 17.43
R1003 vss.n102 vss.t74 17.43
R1004 vss.n101 vss.t43 17.43
R1005 vss.n100 vss.t76 17.43
R1006 vss.n1 vss.n0 0.63
R1007 vss.n2 vss.n1 0.63
R1008 vss.n101 vss.n100 0.63
R1009 vss.n102 vss.n101 0.63
R1010 vss.n13 vss.n12 0.545
R1011 vss.n14 vss.n13 0.545
R1012 vss.n15 vss.n14 0.545
R1013 vss.n22 vss.n21 0.545
R1014 vss.n23 vss.n22 0.545
R1015 vss.n24 vss.n23 0.545
R1016 vss.n31 vss.n30 0.545
R1017 vss.n32 vss.n31 0.545
R1018 vss.n33 vss.n32 0.545
R1019 vss.n40 vss.n39 0.545
R1020 vss.n41 vss.n40 0.545
R1021 vss.n42 vss.n41 0.545
R1022 vss.n47 vss.n46 0.545
R1023 vss.n48 vss.n47 0.545
R1024 vss.n49 vss.n48 0.545
R1025 vss.n53 vss.n52 0.545
R1026 vss.n54 vss.n53 0.545
R1027 vss.n55 vss.n54 0.545
R1028 vss.n62 vss.n61 0.545
R1029 vss.n63 vss.n62 0.545
R1030 vss.n64 vss.n63 0.545
R1031 vss.n71 vss.n70 0.545
R1032 vss.n72 vss.n71 0.545
R1033 vss.n73 vss.n72 0.545
R1034 vss.n80 vss.n79 0.545
R1035 vss.n81 vss.n80 0.545
R1036 vss.n82 vss.n81 0.545
R1037 vss.n89 vss.n88 0.545
R1038 vss.n90 vss.n89 0.545
R1039 vss.n91 vss.n90 0.545
R1040 vss.n96 vss.n95 0.545
R1041 vss.n97 vss.n96 0.545
R1042 vss.n98 vss.n97 0.545
R1043 vss.n16 vss.n15 0.379
R1044 vss.n25 vss.n24 0.379
R1045 vss.n34 vss.n33 0.379
R1046 vss.n43 vss.n42 0.379
R1047 vss.n50 vss.n49 0.379
R1048 vss.n56 vss.n55 0.379
R1049 vss.n65 vss.n64 0.379
R1050 vss.n74 vss.n73 0.379
R1051 vss.n83 vss.n82 0.379
R1052 vss.n92 vss.n91 0.379
R1053 vss.n99 vss.n98 0.379
R1054 vss.n7 vss.n2 0.375
R1055 vss.n106 vss.n102 0.367
R1056 vss.n117 vss.n16 0.197
R1057 vss.n115 vss.n34 0.197
R1058 vss.n113 vss.n50 0.197
R1059 vss.n111 vss.n65 0.197
R1060 vss.n109 vss.n83 0.197
R1061 vss.n107 vss.n99 0.197
R1062 vss.n108 vss.n92 0.197
R1063 vss.n110 vss.n74 0.197
R1064 vss.n112 vss.n56 0.197
R1065 vss.n114 vss.n43 0.197
R1066 vss.n116 vss.n25 0.197
R1067 vss.n94 vss.n93 0.195
R1068 vss.n87 vss.n86 0.195
R1069 vss.n78 vss.n77 0.195
R1070 vss.n69 vss.n68 0.195
R1071 vss.n38 vss.n37 0.195
R1072 vss.n29 vss.n28 0.195
R1073 vss.n20 vss.n19 0.195
R1074 vss.n11 vss.n10 0.195
R1075 vss.n107 vss.n106 0.181
R1076 vss.n118 vss.n7 0.147
R1077 vss vss.n118 0.05
R1078 vss.n108 vss.n107 0.034
R1079 vss.n109 vss.n108 0.034
R1080 vss.n110 vss.n109 0.034
R1081 vss.n111 vss.n110 0.034
R1082 vss.n112 vss.n111 0.034
R1083 vss.n113 vss.n112 0.034
R1084 vss.n114 vss.n113 0.034
R1085 vss.n115 vss.n114 0.034
R1086 vss.n116 vss.n115 0.034
R1087 vss.n117 vss.n116 0.034
R1088 vss.n118 vss.n117 0.033
R1089 vss.n60 vss.n59 0.011
R1090 vss.n45 vss.n44 0.011
R1091 vss.n106 vss.n105 0.008
R1092 vss.n6 vss.n5 0.008
R1093 vss.n104 vss.n103 0.001
R1094 vss.n85 vss.n84 0.001
R1095 vss.n76 vss.n75 0.001
R1096 vss.n67 vss.n66 0.001
R1097 vss.n58 vss.n57 0.001
R1098 vss.n36 vss.n35 0.001
R1099 vss.n27 vss.n26 0.001
R1100 vss.n18 vss.n17 0.001
R1101 vss.n9 vss.n8 0.001
R1102 vss.n4 vss.n3 0.001
R1103 vss.n99 vss.n94 0.001
R1104 vss.n92 vss.n87 0.001
R1105 vss.n83 vss.n78 0.001
R1106 vss.n74 vss.n69 0.001
R1107 vss.n65 vss.n60 0.001
R1108 vss.n56 vss.n51 0.001
R1109 vss.n50 vss.n45 0.001
R1110 vss.n43 vss.n38 0.001
R1111 vss.n34 vss.n29 0.001
R1112 vss.n25 vss.n20 0.001
R1113 vss.n16 vss.n11 0.001
R1114 vss.n7 vss.n6 0.001
R1115 vout.n34 vout.t54 17.43
R1116 vout.n34 vout.t33 17.43
R1117 vout.n33 vout.t25 17.43
R1118 vout.n33 vout.t2 17.43
R1119 vout.n32 vout.t53 17.43
R1120 vout.n32 vout.t32 17.43
R1121 vout.n31 vout.t19 17.43
R1122 vout.n31 vout.t63 17.43
R1123 vout.n38 vout.t27 17.43
R1124 vout.n38 vout.t4 17.43
R1125 vout.n37 vout.t61 17.43
R1126 vout.n37 vout.t38 17.43
R1127 vout.n36 vout.t28 17.43
R1128 vout.n36 vout.t5 17.43
R1129 vout.n35 vout.t59 17.43
R1130 vout.n35 vout.t35 17.43
R1131 vout.n63 vout.t44 17.43
R1132 vout.n63 vout.t29 17.43
R1133 vout.n62 vout.t14 17.43
R1134 vout.n62 vout.t62 17.43
R1135 vout.n61 vout.t43 17.43
R1136 vout.n61 vout.t30 17.43
R1137 vout.n60 vout.t8 17.43
R1138 vout.n60 vout.t60 17.43
R1139 vout.n59 vout.t37 17.43
R1140 vout.n59 vout.t1 17.43
R1141 vout.n58 vout.t6 17.43
R1142 vout.n58 vout.t34 17.43
R1143 vout.n57 vout.t36 17.43
R1144 vout.n57 vout.t0 17.43
R1145 vout.n56 vout.t3 17.43
R1146 vout.n56 vout.t31 17.43
R1147 vout.n55 vout.t10 17.43
R1148 vout.n55 vout.t55 17.43
R1149 vout.n54 vout.t45 17.43
R1150 vout.n54 vout.t26 17.43
R1151 vout.n53 vout.t12 17.43
R1152 vout.n53 vout.t56 17.43
R1153 vout.n52 vout.t39 17.43
R1154 vout.n52 vout.t20 17.43
R1155 vout.n51 vout.t49 17.43
R1156 vout.n51 vout.t11 17.43
R1157 vout.n50 vout.t18 17.43
R1158 vout.n50 vout.t46 17.43
R1159 vout.n49 vout.t48 17.43
R1160 vout.n49 vout.t9 17.43
R1161 vout.n48 vout.t15 17.43
R1162 vout.n48 vout.t40 17.43
R1163 vout.n47 vout.t21 17.43
R1164 vout.n47 vout.t24 17.43
R1165 vout.n46 vout.t57 17.43
R1166 vout.n46 vout.t58 17.43
R1167 vout.n45 vout.t23 17.43
R1168 vout.n45 vout.t22 17.43
R1169 vout.n44 vout.t51 17.43
R1170 vout.n44 vout.t52 17.43
R1171 vout.n43 vout.t16 17.43
R1172 vout.n43 vout.t41 17.43
R1173 vout.n42 vout.t50 17.43
R1174 vout.n42 vout.t13 17.43
R1175 vout.n41 vout.t17 17.43
R1176 vout.n41 vout.t42 17.43
R1177 vout.n40 vout.t47 17.43
R1178 vout.n40 vout.t7 17.43
R1179 vout.n11 vout.t85 14.295
R1180 vout.n11 vout.t66 14.295
R1181 vout.n10 vout.t71 14.295
R1182 vout.n10 vout.t98 14.295
R1183 vout.n9 vout.t82 14.295
R1184 vout.n9 vout.t91 14.295
R1185 vout.n8 vout.t99 14.295
R1186 vout.n8 vout.t106 14.295
R1187 vout.n7 vout.t84 14.295
R1188 vout.n7 vout.t89 14.295
R1189 vout.n6 vout.t107 14.295
R1190 vout.n6 vout.t70 14.295
R1191 vout.n5 vout.t103 14.295
R1192 vout.n5 vout.t73 14.295
R1193 vout.n4 vout.t88 14.295
R1194 vout.n4 vout.t104 14.295
R1195 vout.n3 vout.t72 14.295
R1196 vout.n3 vout.t95 14.295
R1197 vout.n2 vout.t78 14.295
R1198 vout.n2 vout.t90 14.295
R1199 vout.n1 vout.t111 14.295
R1200 vout.n1 vout.t79 14.295
R1201 vout.n0 vout.t76 14.295
R1202 vout.n0 vout.t102 14.295
R1203 vout.n17 vout.t83 14.295
R1204 vout.n17 vout.t64 14.295
R1205 vout.n16 vout.t69 14.295
R1206 vout.n16 vout.t97 14.295
R1207 vout.n15 vout.t96 14.295
R1208 vout.n15 vout.t108 14.295
R1209 vout.n20 vout.t68 14.295
R1210 vout.n20 vout.t67 14.295
R1211 vout.n19 vout.t101 14.295
R1212 vout.n19 vout.t100 14.295
R1213 vout.n18 vout.t86 14.295
R1214 vout.n18 vout.t74 14.295
R1215 vout.n23 vout.t109 14.295
R1216 vout.n23 vout.t87 14.295
R1217 vout.n22 vout.t93 14.295
R1218 vout.n22 vout.t75 14.295
R1219 vout.n21 vout.t65 14.295
R1220 vout.n21 vout.t77 14.295
R1221 vout.n26 vout.t110 14.295
R1222 vout.n26 vout.t92 14.295
R1223 vout.n25 vout.t94 14.295
R1224 vout.n25 vout.t80 14.295
R1225 vout.n24 vout.t105 14.295
R1226 vout.n24 vout.t81 14.295
R1227 vout.n39 vout.n38 1.368
R1228 vout.n64 vout.n63 1.368
R1229 vout vout.n69 1.271
R1230 vout.n12 vout.n11 1.216
R1231 vout.n27 vout.n26 1.216
R1232 vout vout.n30 1.169
R1233 vout.n39 vout.n34 0.74
R1234 vout.n64 vout.n59 0.74
R1235 vout.n65 vout.n55 0.74
R1236 vout.n66 vout.n51 0.74
R1237 vout.n67 vout.n47 0.74
R1238 vout.n68 vout.n43 0.74
R1239 vout.n10 vout.n9 0.733
R1240 vout.n11 vout.n10 0.733
R1241 vout.n7 vout.n6 0.733
R1242 vout.n8 vout.n7 0.733
R1243 vout.n4 vout.n3 0.733
R1244 vout.n5 vout.n4 0.733
R1245 vout.n1 vout.n0 0.733
R1246 vout.n2 vout.n1 0.733
R1247 vout.n16 vout.n15 0.733
R1248 vout.n17 vout.n16 0.733
R1249 vout.n19 vout.n18 0.733
R1250 vout.n20 vout.n19 0.733
R1251 vout.n22 vout.n21 0.733
R1252 vout.n23 vout.n22 0.733
R1253 vout.n25 vout.n24 0.733
R1254 vout.n26 vout.n25 0.733
R1255 vout.n13 vout.n12 0.628
R1256 vout.n14 vout.n13 0.628
R1257 vout.n29 vout.n28 0.628
R1258 vout.n28 vout.n27 0.628
R1259 vout.n68 vout.n67 0.628
R1260 vout.n67 vout.n66 0.628
R1261 vout.n66 vout.n65 0.628
R1262 vout.n65 vout.n64 0.628
R1263 vout.n12 vout.n8 0.588
R1264 vout.n13 vout.n5 0.588
R1265 vout.n14 vout.n2 0.588
R1266 vout.n29 vout.n17 0.588
R1267 vout.n28 vout.n20 0.588
R1268 vout.n27 vout.n23 0.588
R1269 vout.n32 vout.n31 0.545
R1270 vout.n33 vout.n32 0.545
R1271 vout.n34 vout.n33 0.545
R1272 vout.n36 vout.n35 0.545
R1273 vout.n37 vout.n36 0.545
R1274 vout.n38 vout.n37 0.545
R1275 vout.n61 vout.n60 0.545
R1276 vout.n62 vout.n61 0.545
R1277 vout.n63 vout.n62 0.545
R1278 vout.n57 vout.n56 0.545
R1279 vout.n58 vout.n57 0.545
R1280 vout.n59 vout.n58 0.545
R1281 vout.n53 vout.n52 0.545
R1282 vout.n54 vout.n53 0.545
R1283 vout.n55 vout.n54 0.545
R1284 vout.n49 vout.n48 0.545
R1285 vout.n50 vout.n49 0.545
R1286 vout.n51 vout.n50 0.545
R1287 vout.n45 vout.n44 0.545
R1288 vout.n46 vout.n45 0.545
R1289 vout.n47 vout.n46 0.545
R1290 vout.n41 vout.n40 0.545
R1291 vout.n42 vout.n41 0.545
R1292 vout.n43 vout.n42 0.545
R1293 vout.n30 vout.n14 0.53
R1294 vout.n69 vout.n39 0.53
R1295 vout.n30 vout.n29 0.097
R1296 vout.n69 vout.n68 0.097
R1297 a_20875_2019.n2 a_20875_2019.t11 37.645
R1298 a_20875_2019.n2 a_20875_2019.t63 37.361
R1299 a_20875_2019.n6 a_20875_2019.t55 37.361
R1300 a_20875_2019.n5 a_20875_2019.t62 37.361
R1301 a_20875_2019.n5 a_20875_2019.t54 37.361
R1302 a_20875_2019.n2 a_20875_2019.t57 37.361
R1303 a_20875_2019.n0 a_20875_2019.t49 37.361
R1304 a_20875_2019.n1 a_20875_2019.t56 37.361
R1305 a_20875_2019.n1 a_20875_2019.t48 37.361
R1306 a_20875_2019.n5 a_20875_2019.t7 37.361
R1307 a_20875_2019.n5 a_20875_2019.t27 37.361
R1308 a_20875_2019.n4 a_20875_2019.t23 37.361
R1309 a_20875_2019.n6 a_20875_2019.t9 37.361
R1310 a_20875_2019.n6 a_20875_2019.t29 37.361
R1311 a_20875_2019.n5 a_20875_2019.t15 37.361
R1312 a_20875_2019.n5 a_20875_2019.t25 37.361
R1313 a_20875_2019.n1 a_20875_2019.t52 37.361
R1314 a_20875_2019.n1 a_20875_2019.t33 37.361
R1315 a_20875_2019.n1 a_20875_2019.t3 37.361
R1316 a_20875_2019.n1 a_20875_2019.t51 37.361
R1317 a_20875_2019.n1 a_20875_2019.t58 37.361
R1318 a_20875_2019.n0 a_20875_2019.t50 37.361
R1319 a_20875_2019.n3 a_20875_2019.t59 37.361
R1320 a_20875_2019.n3 a_20875_2019.t61 37.361
R1321 a_20875_2019.n3 a_20875_2019.t13 37.361
R1322 a_20875_2019.n3 a_20875_2019.t19 37.361
R1323 a_20875_2019.n1 a_20875_2019.t31 37.361
R1324 a_20875_2019.n1 a_20875_2019.t5 37.361
R1325 a_20875_2019.n1 a_20875_2019.t53 37.361
R1326 a_20875_2019.n1 a_20875_2019.t60 37.361
R1327 a_20875_2019.n1 a_20875_2019.t17 37.361
R1328 a_20875_2019.n1 a_20875_2019.t21 37.361
R1329 a_20875_2019.n1 a_20875_2019.t4 17.43
R1330 a_20875_2019.n3 a_20875_2019.t6 17.43
R1331 a_20875_2019.n3 a_20875_2019.t32 17.43
R1332 a_20875_2019.n5 a_20875_2019.t8 17.43
R1333 a_20875_2019.n5 a_20875_2019.t28 17.43
R1334 a_20875_2019.n4 a_20875_2019.t30 17.43
R1335 a_20875_2019.n4 a_20875_2019.t10 17.43
R1336 a_20875_2019.n4 a_20875_2019.t12 17.43
R1337 a_20875_2019.n4 a_20875_2019.t24 17.43
R1338 a_20875_2019.n5 a_20875_2019.t16 17.43
R1339 a_20875_2019.n5 a_20875_2019.t26 17.43
R1340 a_20875_2019.n3 a_20875_2019.t20 17.43
R1341 a_20875_2019.n3 a_20875_2019.t14 17.43
R1342 a_20875_2019.n1 a_20875_2019.t22 17.43
R1343 a_20875_2019.n1 a_20875_2019.t18 17.43
R1344 a_20875_2019.t34 a_20875_2019.n1 17.43
R1345 a_20875_2019.n22 a_20875_2019.t1 7.146
R1346 a_20875_2019.n22 a_20875_2019.t47 7.146
R1347 a_20875_2019.n21 a_20875_2019.t40 7.146
R1348 a_20875_2019.n21 a_20875_2019.t2 7.146
R1349 a_20875_2019.n20 a_20875_2019.t42 7.146
R1350 a_20875_2019.n20 a_20875_2019.t35 7.146
R1351 a_20875_2019.n19 a_20875_2019.t44 7.146
R1352 a_20875_2019.n19 a_20875_2019.t36 7.146
R1353 a_20875_2019.n15 a_20875_2019.t45 7.146
R1354 a_20875_2019.n15 a_20875_2019.t46 7.146
R1355 a_20875_2019.n14 a_20875_2019.t0 7.146
R1356 a_20875_2019.n14 a_20875_2019.t39 7.146
R1357 a_20875_2019.n13 a_20875_2019.t37 7.146
R1358 a_20875_2019.n13 a_20875_2019.t41 7.146
R1359 a_20875_2019.n12 a_20875_2019.t43 7.146
R1360 a_20875_2019.n12 a_20875_2019.t38 7.146
R1361 a_20875_2019.n5 a_20875_2019.n22 1.777
R1362 a_20875_2019.n1 a_20875_2019.n15 1.583
R1363 a_20875_2019.n3 a_20875_2019.n2 1.388
R1364 a_20875_2019.n5 a_20875_2019.n4 1.13
R1365 a_20875_2019.n1 a_20875_2019.n0 1.122
R1366 a_20875_2019.n3 a_20875_2019.n18 1.076
R1367 a_20875_2019.n20 a_20875_2019.n19 1.045
R1368 a_20875_2019.n21 a_20875_2019.n20 1.045
R1369 a_20875_2019.n22 a_20875_2019.n21 1.045
R1370 a_20875_2019.n13 a_20875_2019.n12 1.045
R1371 a_20875_2019.n14 a_20875_2019.n13 1.045
R1372 a_20875_2019.n15 a_20875_2019.n14 1.045
R1373 a_20875_2019.n0 a_20875_2019.n6 0.989
R1374 a_20875_2019.n1 a_20875_2019.n3 0.901
R1375 a_20875_2019.n1 a_20875_2019.n5 0.841
R1376 a_20875_2019.n1 a_20875_2019.n7 0.82
R1377 a_20875_2019.n17 a_20875_2019.n16 0.603
R1378 a_20875_2019.n10 a_20875_2019.n9 0.603
R1379 a_20875_2019.n11 a_20875_2019.n10 0.603
R1380 a_20875_2019.n18 a_20875_2019.n17 0.603
R1381 a_20875_2019.n7 a_20875_2019.n11 0.603
R1382 a_20875_2019.n9 a_20875_2019.n8 0.602
R1383 vn.n10 vn.t15 111.977
R1384 vn.n21 vn.t14 111.977
R1385 vn.n10 vn.t7 111.975
R1386 vn.n21 vn.t9 111.975
R1387 vn.n1 vn.t0 111.83
R1388 vn.n7 vn.t6 111.83
R1389 vn.n12 vn.t1 111.83
R1390 vn.n18 vn.t8 111.83
R1391 vn.n8 vn.t13 111.83
R1392 vn.n5 vn.t11 111.83
R1393 vn.n2 vn.t3 111.83
R1394 vn.n4 vn.t4 111.83
R1395 vn.n19 vn.t12 111.83
R1396 vn.n16 vn.t10 111.83
R1397 vn.n13 vn.t2 111.83
R1398 vn.n15 vn.t5 111.83
R1399 vn.n22 vn.n10 2.763
R1400 vn.n9 vn.n6 2.018
R1401 vn.n6 vn.n3 2.018
R1402 vn.n20 vn.n17 2.018
R1403 vn.n17 vn.n14 2.018
R1404 vn.n10 vn.n9 2.016
R1405 vn.n21 vn.n20 2.016
R1406 vn.n3 vn.n0 1.995
R1407 vn.n14 vn.n11 1.995
R1408 vn vn.n22 0.811
R1409 vn.n9 vn.n8 0.14
R1410 vn.n6 vn.n5 0.14
R1411 vn.n3 vn.n2 0.14
R1412 vn.n20 vn.n19 0.14
R1413 vn.n17 vn.n16 0.14
R1414 vn.n14 vn.n13 0.14
R1415 vn.n3 vn.n1 0.139
R1416 vn.n6 vn.n4 0.139
R1417 vn.n9 vn.n7 0.139
R1418 vn.n14 vn.n12 0.139
R1419 vn.n17 vn.n15 0.139
R1420 vn.n20 vn.n18 0.139
R1421 vn.n22 vn.n21 0.133
C4 vp vss 7.41fF
C5 vn vss 6.69fF
C6 vout vss 30.11fF
C7 vbias vss 43.40fF
C8 vdd vss 123.75fF
C9 vn.n10 vss 1.27fF $ **FLOATING
C10 a_20875_2019.n0 vss 1.60fF $ **FLOATING
C11 a_20875_2019.n1 vss 7.74fF $ **FLOATING
C12 a_20875_2019.n2 vss 2.47fF $ **FLOATING
C13 a_20875_2019.n3 vss 4.50fF $ **FLOATING
C14 a_20875_2019.n4 vss 2.77fF $ **FLOATING
C15 a_20875_2019.n5 vss 4.15fF $ **FLOATING
C16 a_20875_2019.n6 vss 2.33fF $ **FLOATING
C17 a_20875_2019.n12 vss 1.41fF $ **FLOATING
C18 a_20875_2019.n13 vss 1.46fF $ **FLOATING
C19 a_20875_2019.n14 vss 1.46fF $ **FLOATING
C20 a_20875_2019.n15 vss 1.49fF $ **FLOATING
C21 a_20875_2019.n19 vss 1.41fF $ **FLOATING
C22 a_20875_2019.n20 vss 1.46fF $ **FLOATING
C23 a_20875_2019.n21 vss 1.46fF $ **FLOATING
C24 a_20875_2019.n22 vss 1.59fF $ **FLOATING
C25 vout.n11 vss 1.18fF $ **FLOATING
C26 vout.n12 vss 1.09fF $ **FLOATING
C27 vout.n26 vss 1.18fF $ **FLOATING
C28 vout.n27 vss 1.09fF $ **FLOATING
C29 vout.n30 vss 2.04fF $ **FLOATING
C30 vout.n39 vss 1.06fF $ **FLOATING
C31 vout.n64 vss 1.12fF $ **FLOATING
C32 vout.n69 vss 2.18fF $ **FLOATING
C33 a_21819_2107.n0 vss 1.10fF $ **FLOATING
C34 a_21819_2107.n1 vss 1.06fF $ **FLOATING
C35 a_21819_2107.n2 vss 1.04fF $ **FLOATING
C36 a_21819_2107.n3 vss 1.48fF $ **FLOATING
C37 a_21819_2107.n4 vss 1.53fF $ **FLOATING
C38 a_21819_2107.n84 vss 1.06fF $ **FLOATING
C39 a_21819_2107.n85 vss 1.48fF $ **FLOATING
C40 a_21819_2107.n86 vss 1.53fF $ **FLOATING
C41 a_21819_2107.n87 vss 1.53fF $ **FLOATING
C42 a_21819_2107.n88 vss 1.48fF $ **FLOATING
C43 a_21819_2107.n94 vss 1.84fF $ **FLOATING
C44 a_21819_2107.n96 vss 1.48fF $ **FLOATING
C45 a_21819_2107.n97 vss 1.53fF $ **FLOATING
C46 w_20679_4119.n3 vss 1.58fF $ **FLOATING
C47 w_20679_4119.n5 vss 3.06fF $ **FLOATING
C48 w_20679_4119.n6 vss 3.16fF $ **FLOATING
C49 w_20679_4119.n7 vss 3.16fF $ **FLOATING
C50 w_20679_4119.n8 vss 2.90fF $ **FLOATING
C51 w_20679_4119.n9 vss 1.58fF $ **FLOATING
C52 w_20679_4119.n10 vss 1.68fF $ **FLOATING
C53 w_20679_4119.n11 vss 1.94fF $ **FLOATING
C54 w_20679_4119.n12 vss 3.12fF $ **FLOATING
C55 w_20679_4119.n13 vss 1.76fF $ **FLOATING
C56 w_20679_4119.n14 vss 2.61fF $ **FLOATING
C57 w_20679_4119.n15 vss 3.82fF $ **FLOATING
C58 w_20679_4119.n18 vss 1.58fF $ **FLOATING
C59 w_20679_4119.n19 vss 1.68fF $ **FLOATING
C60 w_20679_4119.n20 vss 1.65fF $ **FLOATING
C61 w_20679_4119.n22 vss 3.06fF $ **FLOATING
C62 w_20679_4119.n23 vss 3.16fF $ **FLOATING
C63 w_20679_4119.n24 vss 3.16fF $ **FLOATING
C64 w_20679_4119.n25 vss 2.90fF $ **FLOATING
C65 w_20679_4119.n26 vss 4.69fF $ **FLOATING
C66 w_20679_4119.n28 vss 3.09fF $ **FLOATING
C67 w_20679_4119.n29 vss 1.74fF $ **FLOATING
C68 w_20679_4119.n30 vss 1.56fF $ **FLOATING
C69 w_20679_4119.n33 vss 1.58fF $ **FLOATING
C70 w_20679_4119.n34 vss 1.68fF $ **FLOATING
C71 w_20679_4119.n35 vss 1.94fF $ **FLOATING
C72 w_20679_4119.n40 vss 3.06fF $ **FLOATING
C73 w_20679_4119.n41 vss 3.16fF $ **FLOATING
C74 w_20679_4119.n42 vss 3.16fF $ **FLOATING
C75 w_20679_4119.n43 vss 3.09fF $ **FLOATING
C76 w_20679_4119.n44 vss 1.25fF $ **FLOATING
C77 w_20679_4119.n48 vss 1.65fF $ **FLOATING
C78 w_20679_4119.n49 vss 1.68fF $ **FLOATING
C79 vdd.n114 vss 1.05fF $ **FLOATING
C80 vdd.n117 vss 3.91fF $ **FLOATING
C81 vdd.n125 vss 10.96fF $ **FLOATING
C82 vdd.n126 vss 6.14fF $ **FLOATING
C83 vdd.n127 vss 6.14fF $ **FLOATING
C84 vdd.n128 vss 6.14fF $ **FLOATING
C85 vdd.n129 vss 6.14fF $ **FLOATING
C86 vdd.n130 vss 6.14fF $ **FLOATING
C87 vdd.n131 vss 6.14fF $ **FLOATING
C88 vdd.n132 vss 4.84fF $ **FLOATING
C89 vdd.n133 vss 4.84fF $ **FLOATING
C90 vdd.n134 vss 6.14fF $ **FLOATING
C91 vdd.n135 vss 6.14fF $ **FLOATING
C92 vdd.n136 vss 6.14fF $ **FLOATING
C93 vdd.n137 vss 6.14fF $ **FLOATING
C94 vdd.n138 vss 6.14fF $ **FLOATING
C95 vdd.n139 vss 4.43fF $ **FLOATING
C96 vdd.n140 vss 3.69fF $ **FLOATING
.ends
