magic
tech sky130A
magscale 1 2
timestamp 1629274976
<< pwell >>
rect -4801 -3309 5715 965
<< nmoslvt >>
rect -4605 -45 -4205 755
rect -4033 -45 -3633 755
rect -3461 -45 -3061 755
rect -2889 -45 -2489 755
rect -2317 -45 -1917 755
rect -1745 -45 -1345 755
rect -1173 -45 -773 755
rect -601 -45 -201 755
rect -29 -45 371 755
rect 543 -45 943 755
rect 1115 -45 1515 755
rect 1687 -45 2087 755
rect 2259 -45 2659 755
rect 2831 -45 3231 755
rect 3403 -45 3803 755
rect 3975 -45 4375 755
rect 4547 -45 4947 755
rect 5119 -45 5519 755
rect -4605 -1063 -4205 -263
rect -4033 -1063 -3633 -263
rect -3461 -1063 -3061 -263
rect -2889 -1063 -2489 -263
rect -2317 -1063 -1917 -263
rect -1745 -1063 -1345 -263
rect -1173 -1063 -773 -263
rect -601 -1063 -201 -263
rect -29 -1063 371 -263
rect 543 -1063 943 -263
rect 1115 -1063 1515 -263
rect 1687 -1063 2087 -263
rect 2259 -1063 2659 -263
rect 2831 -1063 3231 -263
rect 3403 -1063 3803 -263
rect 3975 -1063 4375 -263
rect 4547 -1063 4947 -263
rect 5119 -1063 5519 -263
rect -4605 -2081 -4205 -1281
rect -4033 -2081 -3633 -1281
rect -3461 -2081 -3061 -1281
rect -2889 -2081 -2489 -1281
rect -2317 -2081 -1917 -1281
rect -1745 -2081 -1345 -1281
rect -1173 -2081 -773 -1281
rect -601 -2081 -201 -1281
rect -29 -2081 371 -1281
rect 543 -2081 943 -1281
rect 1115 -2081 1515 -1281
rect 1687 -2081 2087 -1281
rect 2259 -2081 2659 -1281
rect 2831 -2081 3231 -1281
rect 3403 -2081 3803 -1281
rect 3975 -2081 4375 -1281
rect 4547 -2081 4947 -1281
rect 5119 -2081 5519 -1281
rect -4605 -3099 -4205 -2299
rect -4033 -3099 -3633 -2299
rect -3461 -3099 -3061 -2299
rect -2889 -3099 -2489 -2299
rect -2317 -3099 -1917 -2299
rect -1745 -3099 -1345 -2299
rect -1173 -3099 -773 -2299
rect -601 -3099 -201 -2299
rect -29 -3099 371 -2299
rect 543 -3099 943 -2299
rect 1115 -3099 1515 -2299
rect 1687 -3099 2087 -2299
rect 2259 -3099 2659 -2299
rect 2831 -3099 3231 -2299
rect 3403 -3099 3803 -2299
rect 3975 -3099 4375 -2299
rect 4547 -3099 4947 -2299
rect 5119 -3099 5519 -2299
<< ndiff >>
rect -4663 743 -4605 755
rect -4663 -33 -4651 743
rect -4617 -33 -4605 743
rect -4663 -45 -4605 -33
rect -4205 743 -4147 755
rect -4205 -33 -4193 743
rect -4159 -33 -4147 743
rect -4205 -45 -4147 -33
rect -4091 743 -4033 755
rect -4091 -33 -4079 743
rect -4045 -33 -4033 743
rect -4091 -45 -4033 -33
rect -3633 743 -3575 755
rect -3633 -33 -3621 743
rect -3587 -33 -3575 743
rect -3633 -45 -3575 -33
rect -3519 743 -3461 755
rect -3519 -33 -3507 743
rect -3473 -33 -3461 743
rect -3519 -45 -3461 -33
rect -3061 743 -3003 755
rect -3061 -33 -3049 743
rect -3015 -33 -3003 743
rect -3061 -45 -3003 -33
rect -2947 743 -2889 755
rect -2947 -33 -2935 743
rect -2901 -33 -2889 743
rect -2947 -45 -2889 -33
rect -2489 743 -2431 755
rect -2489 -33 -2477 743
rect -2443 -33 -2431 743
rect -2489 -45 -2431 -33
rect -2375 743 -2317 755
rect -2375 -33 -2363 743
rect -2329 -33 -2317 743
rect -2375 -45 -2317 -33
rect -1917 743 -1859 755
rect -1917 -33 -1905 743
rect -1871 -33 -1859 743
rect -1917 -45 -1859 -33
rect -1803 743 -1745 755
rect -1803 -33 -1791 743
rect -1757 -33 -1745 743
rect -1803 -45 -1745 -33
rect -1345 743 -1287 755
rect -1345 -33 -1333 743
rect -1299 -33 -1287 743
rect -1345 -45 -1287 -33
rect -1231 743 -1173 755
rect -1231 -33 -1219 743
rect -1185 -33 -1173 743
rect -1231 -45 -1173 -33
rect -773 743 -715 755
rect -773 -33 -761 743
rect -727 -33 -715 743
rect -773 -45 -715 -33
rect -659 743 -601 755
rect -659 -33 -647 743
rect -613 -33 -601 743
rect -659 -45 -601 -33
rect -201 743 -143 755
rect -201 -33 -189 743
rect -155 -33 -143 743
rect -201 -45 -143 -33
rect -87 743 -29 755
rect -87 -33 -75 743
rect -41 -33 -29 743
rect -87 -45 -29 -33
rect 371 743 429 755
rect 371 -33 383 743
rect 417 -33 429 743
rect 371 -45 429 -33
rect 485 743 543 755
rect 485 -33 497 743
rect 531 -33 543 743
rect 485 -45 543 -33
rect 943 743 1001 755
rect 943 -33 955 743
rect 989 -33 1001 743
rect 943 -45 1001 -33
rect 1057 743 1115 755
rect 1057 -33 1069 743
rect 1103 -33 1115 743
rect 1057 -45 1115 -33
rect 1515 743 1573 755
rect 1515 -33 1527 743
rect 1561 -33 1573 743
rect 1515 -45 1573 -33
rect 1629 743 1687 755
rect 1629 -33 1641 743
rect 1675 -33 1687 743
rect 1629 -45 1687 -33
rect 2087 743 2145 755
rect 2087 -33 2099 743
rect 2133 -33 2145 743
rect 2087 -45 2145 -33
rect 2201 743 2259 755
rect 2201 -33 2213 743
rect 2247 -33 2259 743
rect 2201 -45 2259 -33
rect 2659 743 2717 755
rect 2659 -33 2671 743
rect 2705 -33 2717 743
rect 2659 -45 2717 -33
rect 2773 743 2831 755
rect 2773 -33 2785 743
rect 2819 -33 2831 743
rect 2773 -45 2831 -33
rect 3231 743 3289 755
rect 3231 -33 3243 743
rect 3277 -33 3289 743
rect 3231 -45 3289 -33
rect 3345 743 3403 755
rect 3345 -33 3357 743
rect 3391 -33 3403 743
rect 3345 -45 3403 -33
rect 3803 743 3861 755
rect 3803 -33 3815 743
rect 3849 -33 3861 743
rect 3803 -45 3861 -33
rect 3917 743 3975 755
rect 3917 -33 3929 743
rect 3963 -33 3975 743
rect 3917 -45 3975 -33
rect 4375 743 4433 755
rect 4375 -33 4387 743
rect 4421 -33 4433 743
rect 4375 -45 4433 -33
rect 4489 743 4547 755
rect 4489 -33 4501 743
rect 4535 -33 4547 743
rect 4489 -45 4547 -33
rect 4947 743 5005 755
rect 4947 -33 4959 743
rect 4993 -33 5005 743
rect 4947 -45 5005 -33
rect 5061 743 5119 755
rect 5061 -33 5073 743
rect 5107 -33 5119 743
rect 5061 -45 5119 -33
rect 5519 743 5577 755
rect 5519 -33 5531 743
rect 5565 -33 5577 743
rect 5519 -45 5577 -33
rect -4663 -275 -4605 -263
rect -4663 -1051 -4651 -275
rect -4617 -1051 -4605 -275
rect -4663 -1063 -4605 -1051
rect -4205 -275 -4147 -263
rect -4205 -1051 -4193 -275
rect -4159 -1051 -4147 -275
rect -4205 -1063 -4147 -1051
rect -4091 -275 -4033 -263
rect -4091 -1051 -4079 -275
rect -4045 -1051 -4033 -275
rect -4091 -1063 -4033 -1051
rect -3633 -275 -3575 -263
rect -3633 -1051 -3621 -275
rect -3587 -1051 -3575 -275
rect -3633 -1063 -3575 -1051
rect -3519 -275 -3461 -263
rect -3519 -1051 -3507 -275
rect -3473 -1051 -3461 -275
rect -3519 -1063 -3461 -1051
rect -3061 -275 -3003 -263
rect -3061 -1051 -3049 -275
rect -3015 -1051 -3003 -275
rect -3061 -1063 -3003 -1051
rect -2947 -275 -2889 -263
rect -2947 -1051 -2935 -275
rect -2901 -1051 -2889 -275
rect -2947 -1063 -2889 -1051
rect -2489 -275 -2431 -263
rect -2489 -1051 -2477 -275
rect -2443 -1051 -2431 -275
rect -2489 -1063 -2431 -1051
rect -2375 -275 -2317 -263
rect -2375 -1051 -2363 -275
rect -2329 -1051 -2317 -275
rect -2375 -1063 -2317 -1051
rect -1917 -275 -1859 -263
rect -1917 -1051 -1905 -275
rect -1871 -1051 -1859 -275
rect -1917 -1063 -1859 -1051
rect -1803 -275 -1745 -263
rect -1803 -1051 -1791 -275
rect -1757 -1051 -1745 -275
rect -1803 -1063 -1745 -1051
rect -1345 -275 -1287 -263
rect -1345 -1051 -1333 -275
rect -1299 -1051 -1287 -275
rect -1345 -1063 -1287 -1051
rect -1231 -275 -1173 -263
rect -1231 -1051 -1219 -275
rect -1185 -1051 -1173 -275
rect -1231 -1063 -1173 -1051
rect -773 -275 -715 -263
rect -773 -1051 -761 -275
rect -727 -1051 -715 -275
rect -773 -1063 -715 -1051
rect -659 -275 -601 -263
rect -659 -1051 -647 -275
rect -613 -1051 -601 -275
rect -659 -1063 -601 -1051
rect -201 -275 -143 -263
rect -201 -1051 -189 -275
rect -155 -1051 -143 -275
rect -201 -1063 -143 -1051
rect -87 -275 -29 -263
rect -87 -1051 -75 -275
rect -41 -1051 -29 -275
rect -87 -1063 -29 -1051
rect 371 -275 429 -263
rect 371 -1051 383 -275
rect 417 -1051 429 -275
rect 371 -1063 429 -1051
rect 485 -275 543 -263
rect 485 -1051 497 -275
rect 531 -1051 543 -275
rect 485 -1063 543 -1051
rect 943 -275 1001 -263
rect 943 -1051 955 -275
rect 989 -1051 1001 -275
rect 943 -1063 1001 -1051
rect 1057 -275 1115 -263
rect 1057 -1051 1069 -275
rect 1103 -1051 1115 -275
rect 1057 -1063 1115 -1051
rect 1515 -275 1573 -263
rect 1515 -1051 1527 -275
rect 1561 -1051 1573 -275
rect 1515 -1063 1573 -1051
rect 1629 -275 1687 -263
rect 1629 -1051 1641 -275
rect 1675 -1051 1687 -275
rect 1629 -1063 1687 -1051
rect 2087 -275 2145 -263
rect 2087 -1051 2099 -275
rect 2133 -1051 2145 -275
rect 2087 -1063 2145 -1051
rect 2201 -275 2259 -263
rect 2201 -1051 2213 -275
rect 2247 -1051 2259 -275
rect 2201 -1063 2259 -1051
rect 2659 -275 2717 -263
rect 2659 -1051 2671 -275
rect 2705 -1051 2717 -275
rect 2659 -1063 2717 -1051
rect 2773 -275 2831 -263
rect 2773 -1051 2785 -275
rect 2819 -1051 2831 -275
rect 2773 -1063 2831 -1051
rect 3231 -275 3289 -263
rect 3231 -1051 3243 -275
rect 3277 -1051 3289 -275
rect 3231 -1063 3289 -1051
rect 3345 -275 3403 -263
rect 3345 -1051 3357 -275
rect 3391 -1051 3403 -275
rect 3345 -1063 3403 -1051
rect 3803 -275 3861 -263
rect 3803 -1051 3815 -275
rect 3849 -1051 3861 -275
rect 3803 -1063 3861 -1051
rect 3917 -275 3975 -263
rect 3917 -1051 3929 -275
rect 3963 -1051 3975 -275
rect 3917 -1063 3975 -1051
rect 4375 -275 4433 -263
rect 4375 -1051 4387 -275
rect 4421 -1051 4433 -275
rect 4375 -1063 4433 -1051
rect 4489 -275 4547 -263
rect 4489 -1051 4501 -275
rect 4535 -1051 4547 -275
rect 4489 -1063 4547 -1051
rect 4947 -275 5005 -263
rect 4947 -1051 4959 -275
rect 4993 -1051 5005 -275
rect 4947 -1063 5005 -1051
rect 5061 -275 5119 -263
rect 5061 -1051 5073 -275
rect 5107 -1051 5119 -275
rect 5061 -1063 5119 -1051
rect 5519 -275 5577 -263
rect 5519 -1051 5531 -275
rect 5565 -1051 5577 -275
rect 5519 -1063 5577 -1051
rect -4663 -1293 -4605 -1281
rect -4663 -2069 -4651 -1293
rect -4617 -2069 -4605 -1293
rect -4663 -2081 -4605 -2069
rect -4205 -1293 -4147 -1281
rect -4205 -2069 -4193 -1293
rect -4159 -2069 -4147 -1293
rect -4205 -2081 -4147 -2069
rect -4091 -1293 -4033 -1281
rect -4091 -2069 -4079 -1293
rect -4045 -2069 -4033 -1293
rect -4091 -2081 -4033 -2069
rect -3633 -1293 -3575 -1281
rect -3633 -2069 -3621 -1293
rect -3587 -2069 -3575 -1293
rect -3633 -2081 -3575 -2069
rect -3519 -1293 -3461 -1281
rect -3519 -2069 -3507 -1293
rect -3473 -2069 -3461 -1293
rect -3519 -2081 -3461 -2069
rect -3061 -1293 -3003 -1281
rect -3061 -2069 -3049 -1293
rect -3015 -2069 -3003 -1293
rect -3061 -2081 -3003 -2069
rect -2947 -1293 -2889 -1281
rect -2947 -2069 -2935 -1293
rect -2901 -2069 -2889 -1293
rect -2947 -2081 -2889 -2069
rect -2489 -1293 -2431 -1281
rect -2489 -2069 -2477 -1293
rect -2443 -2069 -2431 -1293
rect -2489 -2081 -2431 -2069
rect -2375 -1293 -2317 -1281
rect -2375 -2069 -2363 -1293
rect -2329 -2069 -2317 -1293
rect -2375 -2081 -2317 -2069
rect -1917 -1293 -1859 -1281
rect -1917 -2069 -1905 -1293
rect -1871 -2069 -1859 -1293
rect -1917 -2081 -1859 -2069
rect -1803 -1293 -1745 -1281
rect -1803 -2069 -1791 -1293
rect -1757 -2069 -1745 -1293
rect -1803 -2081 -1745 -2069
rect -1345 -1293 -1287 -1281
rect -1345 -2069 -1333 -1293
rect -1299 -2069 -1287 -1293
rect -1345 -2081 -1287 -2069
rect -1231 -1293 -1173 -1281
rect -1231 -2069 -1219 -1293
rect -1185 -2069 -1173 -1293
rect -1231 -2081 -1173 -2069
rect -773 -1293 -715 -1281
rect -773 -2069 -761 -1293
rect -727 -2069 -715 -1293
rect -773 -2081 -715 -2069
rect -659 -1293 -601 -1281
rect -659 -2069 -647 -1293
rect -613 -2069 -601 -1293
rect -659 -2081 -601 -2069
rect -201 -1293 -143 -1281
rect -201 -2069 -189 -1293
rect -155 -2069 -143 -1293
rect -201 -2081 -143 -2069
rect -87 -1293 -29 -1281
rect -87 -2069 -75 -1293
rect -41 -2069 -29 -1293
rect -87 -2081 -29 -2069
rect 371 -1293 429 -1281
rect 371 -2069 383 -1293
rect 417 -2069 429 -1293
rect 371 -2081 429 -2069
rect 485 -1293 543 -1281
rect 485 -2069 497 -1293
rect 531 -2069 543 -1293
rect 485 -2081 543 -2069
rect 943 -1293 1001 -1281
rect 943 -2069 955 -1293
rect 989 -2069 1001 -1293
rect 943 -2081 1001 -2069
rect 1057 -1293 1115 -1281
rect 1057 -2069 1069 -1293
rect 1103 -2069 1115 -1293
rect 1057 -2081 1115 -2069
rect 1515 -1293 1573 -1281
rect 1515 -2069 1527 -1293
rect 1561 -2069 1573 -1293
rect 1515 -2081 1573 -2069
rect 1629 -1293 1687 -1281
rect 1629 -2069 1641 -1293
rect 1675 -2069 1687 -1293
rect 1629 -2081 1687 -2069
rect 2087 -1293 2145 -1281
rect 2087 -2069 2099 -1293
rect 2133 -2069 2145 -1293
rect 2087 -2081 2145 -2069
rect 2201 -1293 2259 -1281
rect 2201 -2069 2213 -1293
rect 2247 -2069 2259 -1293
rect 2201 -2081 2259 -2069
rect 2659 -1293 2717 -1281
rect 2659 -2069 2671 -1293
rect 2705 -2069 2717 -1293
rect 2659 -2081 2717 -2069
rect 2773 -1293 2831 -1281
rect 2773 -2069 2785 -1293
rect 2819 -2069 2831 -1293
rect 2773 -2081 2831 -2069
rect 3231 -1293 3289 -1281
rect 3231 -2069 3243 -1293
rect 3277 -2069 3289 -1293
rect 3231 -2081 3289 -2069
rect 3345 -1293 3403 -1281
rect 3345 -2069 3357 -1293
rect 3391 -2069 3403 -1293
rect 3345 -2081 3403 -2069
rect 3803 -1293 3861 -1281
rect 3803 -2069 3815 -1293
rect 3849 -2069 3861 -1293
rect 3803 -2081 3861 -2069
rect 3917 -1293 3975 -1281
rect 3917 -2069 3929 -1293
rect 3963 -2069 3975 -1293
rect 3917 -2081 3975 -2069
rect 4375 -1293 4433 -1281
rect 4375 -2069 4387 -1293
rect 4421 -2069 4433 -1293
rect 4375 -2081 4433 -2069
rect 4489 -1293 4547 -1281
rect 4489 -2069 4501 -1293
rect 4535 -2069 4547 -1293
rect 4489 -2081 4547 -2069
rect 4947 -1293 5005 -1281
rect 4947 -2069 4959 -1293
rect 4993 -2069 5005 -1293
rect 4947 -2081 5005 -2069
rect 5061 -1293 5119 -1281
rect 5061 -2069 5073 -1293
rect 5107 -2069 5119 -1293
rect 5061 -2081 5119 -2069
rect 5519 -1293 5577 -1281
rect 5519 -2069 5531 -1293
rect 5565 -2069 5577 -1293
rect 5519 -2081 5577 -2069
rect -4663 -2311 -4605 -2299
rect -4663 -3087 -4651 -2311
rect -4617 -3087 -4605 -2311
rect -4663 -3099 -4605 -3087
rect -4205 -2311 -4147 -2299
rect -4205 -3087 -4193 -2311
rect -4159 -3087 -4147 -2311
rect -4205 -3099 -4147 -3087
rect -4091 -2311 -4033 -2299
rect -4091 -3087 -4079 -2311
rect -4045 -3087 -4033 -2311
rect -4091 -3099 -4033 -3087
rect -3633 -2311 -3575 -2299
rect -3633 -3087 -3621 -2311
rect -3587 -3087 -3575 -2311
rect -3633 -3099 -3575 -3087
rect -3519 -2311 -3461 -2299
rect -3519 -3087 -3507 -2311
rect -3473 -3087 -3461 -2311
rect -3519 -3099 -3461 -3087
rect -3061 -2311 -3003 -2299
rect -3061 -3087 -3049 -2311
rect -3015 -3087 -3003 -2311
rect -3061 -3099 -3003 -3087
rect -2947 -2311 -2889 -2299
rect -2947 -3087 -2935 -2311
rect -2901 -3087 -2889 -2311
rect -2947 -3099 -2889 -3087
rect -2489 -2311 -2431 -2299
rect -2489 -3087 -2477 -2311
rect -2443 -3087 -2431 -2311
rect -2489 -3099 -2431 -3087
rect -2375 -2311 -2317 -2299
rect -2375 -3087 -2363 -2311
rect -2329 -3087 -2317 -2311
rect -2375 -3099 -2317 -3087
rect -1917 -2311 -1859 -2299
rect -1917 -3087 -1905 -2311
rect -1871 -3087 -1859 -2311
rect -1917 -3099 -1859 -3087
rect -1803 -2311 -1745 -2299
rect -1803 -3087 -1791 -2311
rect -1757 -3087 -1745 -2311
rect -1803 -3099 -1745 -3087
rect -1345 -2311 -1287 -2299
rect -1345 -3087 -1333 -2311
rect -1299 -3087 -1287 -2311
rect -1345 -3099 -1287 -3087
rect -1231 -2311 -1173 -2299
rect -1231 -3087 -1219 -2311
rect -1185 -3087 -1173 -2311
rect -1231 -3099 -1173 -3087
rect -773 -2311 -715 -2299
rect -773 -3087 -761 -2311
rect -727 -3087 -715 -2311
rect -773 -3099 -715 -3087
rect -659 -2311 -601 -2299
rect -659 -3087 -647 -2311
rect -613 -3087 -601 -2311
rect -659 -3099 -601 -3087
rect -201 -2311 -143 -2299
rect -201 -3087 -189 -2311
rect -155 -3087 -143 -2311
rect -201 -3099 -143 -3087
rect -87 -2311 -29 -2299
rect -87 -3087 -75 -2311
rect -41 -3087 -29 -2311
rect -87 -3099 -29 -3087
rect 371 -2311 429 -2299
rect 371 -3087 383 -2311
rect 417 -3087 429 -2311
rect 371 -3099 429 -3087
rect 485 -2311 543 -2299
rect 485 -3087 497 -2311
rect 531 -3087 543 -2311
rect 485 -3099 543 -3087
rect 943 -2311 1001 -2299
rect 943 -3087 955 -2311
rect 989 -3087 1001 -2311
rect 943 -3099 1001 -3087
rect 1057 -2311 1115 -2299
rect 1057 -3087 1069 -2311
rect 1103 -3087 1115 -2311
rect 1057 -3099 1115 -3087
rect 1515 -2311 1573 -2299
rect 1515 -3087 1527 -2311
rect 1561 -3087 1573 -2311
rect 1515 -3099 1573 -3087
rect 1629 -2311 1687 -2299
rect 1629 -3087 1641 -2311
rect 1675 -3087 1687 -2311
rect 1629 -3099 1687 -3087
rect 2087 -2311 2145 -2299
rect 2087 -3087 2099 -2311
rect 2133 -3087 2145 -2311
rect 2087 -3099 2145 -3087
rect 2201 -2311 2259 -2299
rect 2201 -3087 2213 -2311
rect 2247 -3087 2259 -2311
rect 2201 -3099 2259 -3087
rect 2659 -2311 2717 -2299
rect 2659 -3087 2671 -2311
rect 2705 -3087 2717 -2311
rect 2659 -3099 2717 -3087
rect 2773 -2311 2831 -2299
rect 2773 -3087 2785 -2311
rect 2819 -3087 2831 -2311
rect 2773 -3099 2831 -3087
rect 3231 -2311 3289 -2299
rect 3231 -3087 3243 -2311
rect 3277 -3087 3289 -2311
rect 3231 -3099 3289 -3087
rect 3345 -2311 3403 -2299
rect 3345 -3087 3357 -2311
rect 3391 -3087 3403 -2311
rect 3345 -3099 3403 -3087
rect 3803 -2311 3861 -2299
rect 3803 -3087 3815 -2311
rect 3849 -3087 3861 -2311
rect 3803 -3099 3861 -3087
rect 3917 -2311 3975 -2299
rect 3917 -3087 3929 -2311
rect 3963 -3087 3975 -2311
rect 3917 -3099 3975 -3087
rect 4375 -2311 4433 -2299
rect 4375 -3087 4387 -2311
rect 4421 -3087 4433 -2311
rect 4375 -3099 4433 -3087
rect 4489 -2311 4547 -2299
rect 4489 -3087 4501 -2311
rect 4535 -3087 4547 -2311
rect 4489 -3099 4547 -3087
rect 4947 -2311 5005 -2299
rect 4947 -3087 4959 -2311
rect 4993 -3087 5005 -2311
rect 4947 -3099 5005 -3087
rect 5061 -2311 5119 -2299
rect 5061 -3087 5073 -2311
rect 5107 -3087 5119 -2311
rect 5061 -3099 5119 -3087
rect 5519 -2311 5577 -2299
rect 5519 -3087 5531 -2311
rect 5565 -3087 5577 -2311
rect 5519 -3099 5577 -3087
<< ndiffc >>
rect -4651 -33 -4617 743
rect -4193 -33 -4159 743
rect -4079 -33 -4045 743
rect -3621 -33 -3587 743
rect -3507 -33 -3473 743
rect -3049 -33 -3015 743
rect -2935 -33 -2901 743
rect -2477 -33 -2443 743
rect -2363 -33 -2329 743
rect -1905 -33 -1871 743
rect -1791 -33 -1757 743
rect -1333 -33 -1299 743
rect -1219 -33 -1185 743
rect -761 -33 -727 743
rect -647 -33 -613 743
rect -189 -33 -155 743
rect -75 -33 -41 743
rect 383 -33 417 743
rect 497 -33 531 743
rect 955 -33 989 743
rect 1069 -33 1103 743
rect 1527 -33 1561 743
rect 1641 -33 1675 743
rect 2099 -33 2133 743
rect 2213 -33 2247 743
rect 2671 -33 2705 743
rect 2785 -33 2819 743
rect 3243 -33 3277 743
rect 3357 -33 3391 743
rect 3815 -33 3849 743
rect 3929 -33 3963 743
rect 4387 -33 4421 743
rect 4501 -33 4535 743
rect 4959 -33 4993 743
rect 5073 -33 5107 743
rect 5531 -33 5565 743
rect -4651 -1051 -4617 -275
rect -4193 -1051 -4159 -275
rect -4079 -1051 -4045 -275
rect -3621 -1051 -3587 -275
rect -3507 -1051 -3473 -275
rect -3049 -1051 -3015 -275
rect -2935 -1051 -2901 -275
rect -2477 -1051 -2443 -275
rect -2363 -1051 -2329 -275
rect -1905 -1051 -1871 -275
rect -1791 -1051 -1757 -275
rect -1333 -1051 -1299 -275
rect -1219 -1051 -1185 -275
rect -761 -1051 -727 -275
rect -647 -1051 -613 -275
rect -189 -1051 -155 -275
rect -75 -1051 -41 -275
rect 383 -1051 417 -275
rect 497 -1051 531 -275
rect 955 -1051 989 -275
rect 1069 -1051 1103 -275
rect 1527 -1051 1561 -275
rect 1641 -1051 1675 -275
rect 2099 -1051 2133 -275
rect 2213 -1051 2247 -275
rect 2671 -1051 2705 -275
rect 2785 -1051 2819 -275
rect 3243 -1051 3277 -275
rect 3357 -1051 3391 -275
rect 3815 -1051 3849 -275
rect 3929 -1051 3963 -275
rect 4387 -1051 4421 -275
rect 4501 -1051 4535 -275
rect 4959 -1051 4993 -275
rect 5073 -1051 5107 -275
rect 5531 -1051 5565 -275
rect -4651 -2069 -4617 -1293
rect -4193 -2069 -4159 -1293
rect -4079 -2069 -4045 -1293
rect -3621 -2069 -3587 -1293
rect -3507 -2069 -3473 -1293
rect -3049 -2069 -3015 -1293
rect -2935 -2069 -2901 -1293
rect -2477 -2069 -2443 -1293
rect -2363 -2069 -2329 -1293
rect -1905 -2069 -1871 -1293
rect -1791 -2069 -1757 -1293
rect -1333 -2069 -1299 -1293
rect -1219 -2069 -1185 -1293
rect -761 -2069 -727 -1293
rect -647 -2069 -613 -1293
rect -189 -2069 -155 -1293
rect -75 -2069 -41 -1293
rect 383 -2069 417 -1293
rect 497 -2069 531 -1293
rect 955 -2069 989 -1293
rect 1069 -2069 1103 -1293
rect 1527 -2069 1561 -1293
rect 1641 -2069 1675 -1293
rect 2099 -2069 2133 -1293
rect 2213 -2069 2247 -1293
rect 2671 -2069 2705 -1293
rect 2785 -2069 2819 -1293
rect 3243 -2069 3277 -1293
rect 3357 -2069 3391 -1293
rect 3815 -2069 3849 -1293
rect 3929 -2069 3963 -1293
rect 4387 -2069 4421 -1293
rect 4501 -2069 4535 -1293
rect 4959 -2069 4993 -1293
rect 5073 -2069 5107 -1293
rect 5531 -2069 5565 -1293
rect -4651 -3087 -4617 -2311
rect -4193 -3087 -4159 -2311
rect -4079 -3087 -4045 -2311
rect -3621 -3087 -3587 -2311
rect -3507 -3087 -3473 -2311
rect -3049 -3087 -3015 -2311
rect -2935 -3087 -2901 -2311
rect -2477 -3087 -2443 -2311
rect -2363 -3087 -2329 -2311
rect -1905 -3087 -1871 -2311
rect -1791 -3087 -1757 -2311
rect -1333 -3087 -1299 -2311
rect -1219 -3087 -1185 -2311
rect -761 -3087 -727 -2311
rect -647 -3087 -613 -2311
rect -189 -3087 -155 -2311
rect -75 -3087 -41 -2311
rect 383 -3087 417 -2311
rect 497 -3087 531 -2311
rect 955 -3087 989 -2311
rect 1069 -3087 1103 -2311
rect 1527 -3087 1561 -2311
rect 1641 -3087 1675 -2311
rect 2099 -3087 2133 -2311
rect 2213 -3087 2247 -2311
rect 2671 -3087 2705 -2311
rect 2785 -3087 2819 -2311
rect 3243 -3087 3277 -2311
rect 3357 -3087 3391 -2311
rect 3815 -3087 3849 -2311
rect 3929 -3087 3963 -2311
rect 4387 -3087 4421 -2311
rect 4501 -3087 4535 -2311
rect 4959 -3087 4993 -2311
rect 5073 -3087 5107 -2311
rect 5531 -3087 5565 -2311
<< psubdiff >>
rect -4765 895 -4669 929
rect 5583 895 5679 929
rect -4765 833 -4731 895
rect 5645 833 5679 895
rect -4765 -3239 -4731 -3177
rect 5645 -3239 5679 -3177
rect -4765 -3273 -4669 -3239
rect 5583 -3273 5679 -3239
<< psubdiffcont >>
rect -4669 895 5583 929
rect -4765 -3177 -4731 833
rect 5645 -3177 5679 833
rect -4669 -3273 5583 -3239
<< poly >>
rect -4605 827 -4205 843
rect -4605 793 -4589 827
rect -4221 793 -4205 827
rect -4605 755 -4205 793
rect -4033 827 -3633 843
rect -4033 793 -4017 827
rect -3649 793 -3633 827
rect -4033 755 -3633 793
rect -3461 827 -3061 843
rect -3461 793 -3445 827
rect -3077 793 -3061 827
rect -3461 755 -3061 793
rect -2889 827 -2489 843
rect -2889 793 -2873 827
rect -2505 793 -2489 827
rect -2889 755 -2489 793
rect -2317 827 -1917 843
rect -2317 793 -2301 827
rect -1933 793 -1917 827
rect -2317 755 -1917 793
rect -1745 827 -1345 843
rect -1745 793 -1729 827
rect -1361 793 -1345 827
rect -1745 755 -1345 793
rect -1173 827 -773 843
rect -1173 793 -1157 827
rect -789 793 -773 827
rect -1173 755 -773 793
rect -601 827 -201 843
rect -601 793 -585 827
rect -217 793 -201 827
rect -601 755 -201 793
rect -29 827 371 843
rect -29 793 -13 827
rect 355 793 371 827
rect -29 755 371 793
rect 543 827 943 843
rect 543 793 559 827
rect 927 793 943 827
rect 543 755 943 793
rect 1115 827 1515 843
rect 1115 793 1131 827
rect 1499 793 1515 827
rect 1115 755 1515 793
rect 1687 827 2087 843
rect 1687 793 1703 827
rect 2071 793 2087 827
rect 1687 755 2087 793
rect 2259 827 2659 843
rect 2259 793 2275 827
rect 2643 793 2659 827
rect 2259 755 2659 793
rect 2831 827 3231 843
rect 2831 793 2847 827
rect 3215 793 3231 827
rect 2831 755 3231 793
rect 3403 827 3803 843
rect 3403 793 3419 827
rect 3787 793 3803 827
rect 3403 755 3803 793
rect 3975 827 4375 843
rect 3975 793 3991 827
rect 4359 793 4375 827
rect 3975 755 4375 793
rect 4547 827 4947 843
rect 4547 793 4563 827
rect 4931 793 4947 827
rect 4547 755 4947 793
rect 5119 827 5519 843
rect 5119 793 5135 827
rect 5503 793 5519 827
rect 5119 755 5519 793
rect -4605 -83 -4205 -45
rect -4605 -117 -4589 -83
rect -4221 -117 -4205 -83
rect -4605 -133 -4205 -117
rect -4033 -83 -3633 -45
rect -4033 -117 -4017 -83
rect -3649 -117 -3633 -83
rect -4033 -133 -3633 -117
rect -3461 -83 -3061 -45
rect -3461 -117 -3445 -83
rect -3077 -117 -3061 -83
rect -3461 -133 -3061 -117
rect -2889 -83 -2489 -45
rect -2889 -117 -2873 -83
rect -2505 -117 -2489 -83
rect -2889 -133 -2489 -117
rect -2317 -83 -1917 -45
rect -2317 -117 -2301 -83
rect -1933 -117 -1917 -83
rect -2317 -133 -1917 -117
rect -1745 -83 -1345 -45
rect -1745 -117 -1729 -83
rect -1361 -117 -1345 -83
rect -1745 -133 -1345 -117
rect -1173 -83 -773 -45
rect -1173 -117 -1157 -83
rect -789 -117 -773 -83
rect -1173 -133 -773 -117
rect -601 -83 -201 -45
rect -601 -117 -585 -83
rect -217 -117 -201 -83
rect -601 -133 -201 -117
rect -29 -83 371 -45
rect -29 -117 -13 -83
rect 355 -117 371 -83
rect -29 -133 371 -117
rect 543 -83 943 -45
rect 543 -117 559 -83
rect 927 -117 943 -83
rect 543 -133 943 -117
rect 1115 -83 1515 -45
rect 1115 -117 1131 -83
rect 1499 -117 1515 -83
rect 1115 -133 1515 -117
rect 1687 -83 2087 -45
rect 1687 -117 1703 -83
rect 2071 -117 2087 -83
rect 1687 -133 2087 -117
rect 2259 -83 2659 -45
rect 2259 -117 2275 -83
rect 2643 -117 2659 -83
rect 2259 -133 2659 -117
rect 2831 -83 3231 -45
rect 2831 -117 2847 -83
rect 3215 -117 3231 -83
rect 2831 -133 3231 -117
rect 3403 -83 3803 -45
rect 3403 -117 3419 -83
rect 3787 -117 3803 -83
rect 3403 -133 3803 -117
rect 3975 -83 4375 -45
rect 3975 -117 3991 -83
rect 4359 -117 4375 -83
rect 3975 -133 4375 -117
rect 4547 -83 4947 -45
rect 4547 -117 4563 -83
rect 4931 -117 4947 -83
rect 4547 -133 4947 -117
rect 5119 -83 5519 -45
rect 5119 -117 5135 -83
rect 5503 -117 5519 -83
rect 5119 -133 5519 -117
rect -4605 -191 -4205 -175
rect -4605 -225 -4589 -191
rect -4221 -225 -4205 -191
rect -4605 -263 -4205 -225
rect -4033 -191 -3633 -175
rect -4033 -225 -4017 -191
rect -3649 -225 -3633 -191
rect -4033 -263 -3633 -225
rect -3461 -191 -3061 -175
rect -3461 -225 -3445 -191
rect -3077 -225 -3061 -191
rect -3461 -263 -3061 -225
rect -2889 -191 -2489 -175
rect -2889 -225 -2873 -191
rect -2505 -225 -2489 -191
rect -2889 -263 -2489 -225
rect -2317 -191 -1917 -175
rect -2317 -225 -2301 -191
rect -1933 -225 -1917 -191
rect -2317 -263 -1917 -225
rect -1745 -191 -1345 -175
rect -1745 -225 -1729 -191
rect -1361 -225 -1345 -191
rect -1745 -263 -1345 -225
rect -1173 -191 -773 -175
rect -1173 -225 -1157 -191
rect -789 -225 -773 -191
rect -1173 -263 -773 -225
rect -601 -191 -201 -175
rect -601 -225 -585 -191
rect -217 -225 -201 -191
rect -601 -263 -201 -225
rect -29 -191 371 -175
rect -29 -225 -13 -191
rect 355 -225 371 -191
rect -29 -263 371 -225
rect 543 -191 943 -175
rect 543 -225 559 -191
rect 927 -225 943 -191
rect 543 -263 943 -225
rect 1115 -191 1515 -175
rect 1115 -225 1131 -191
rect 1499 -225 1515 -191
rect 1115 -263 1515 -225
rect 1687 -191 2087 -175
rect 1687 -225 1703 -191
rect 2071 -225 2087 -191
rect 1687 -263 2087 -225
rect 2259 -191 2659 -175
rect 2259 -225 2275 -191
rect 2643 -225 2659 -191
rect 2259 -263 2659 -225
rect 2831 -191 3231 -175
rect 2831 -225 2847 -191
rect 3215 -225 3231 -191
rect 2831 -263 3231 -225
rect 3403 -191 3803 -175
rect 3403 -225 3419 -191
rect 3787 -225 3803 -191
rect 3403 -263 3803 -225
rect 3975 -191 4375 -175
rect 3975 -225 3991 -191
rect 4359 -225 4375 -191
rect 3975 -263 4375 -225
rect 4547 -191 4947 -175
rect 4547 -225 4563 -191
rect 4931 -225 4947 -191
rect 4547 -263 4947 -225
rect 5119 -191 5519 -175
rect 5119 -225 5135 -191
rect 5503 -225 5519 -191
rect 5119 -263 5519 -225
rect -4605 -1101 -4205 -1063
rect -4605 -1135 -4589 -1101
rect -4221 -1135 -4205 -1101
rect -4605 -1151 -4205 -1135
rect -4033 -1101 -3633 -1063
rect -4033 -1135 -4017 -1101
rect -3649 -1135 -3633 -1101
rect -4033 -1151 -3633 -1135
rect -3461 -1101 -3061 -1063
rect -3461 -1135 -3445 -1101
rect -3077 -1135 -3061 -1101
rect -3461 -1151 -3061 -1135
rect -2889 -1101 -2489 -1063
rect -2889 -1135 -2873 -1101
rect -2505 -1135 -2489 -1101
rect -2889 -1151 -2489 -1135
rect -2317 -1101 -1917 -1063
rect -2317 -1135 -2301 -1101
rect -1933 -1135 -1917 -1101
rect -2317 -1151 -1917 -1135
rect -1745 -1101 -1345 -1063
rect -1745 -1135 -1729 -1101
rect -1361 -1135 -1345 -1101
rect -1745 -1151 -1345 -1135
rect -1173 -1101 -773 -1063
rect -1173 -1135 -1157 -1101
rect -789 -1135 -773 -1101
rect -1173 -1151 -773 -1135
rect -601 -1101 -201 -1063
rect -601 -1135 -585 -1101
rect -217 -1135 -201 -1101
rect -601 -1151 -201 -1135
rect -29 -1101 371 -1063
rect -29 -1135 -13 -1101
rect 355 -1135 371 -1101
rect -29 -1151 371 -1135
rect 543 -1101 943 -1063
rect 543 -1135 559 -1101
rect 927 -1135 943 -1101
rect 543 -1151 943 -1135
rect 1115 -1101 1515 -1063
rect 1115 -1135 1131 -1101
rect 1499 -1135 1515 -1101
rect 1115 -1151 1515 -1135
rect 1687 -1101 2087 -1063
rect 1687 -1135 1703 -1101
rect 2071 -1135 2087 -1101
rect 1687 -1151 2087 -1135
rect 2259 -1101 2659 -1063
rect 2259 -1135 2275 -1101
rect 2643 -1135 2659 -1101
rect 2259 -1151 2659 -1135
rect 2831 -1101 3231 -1063
rect 2831 -1135 2847 -1101
rect 3215 -1135 3231 -1101
rect 2831 -1151 3231 -1135
rect 3403 -1101 3803 -1063
rect 3403 -1135 3419 -1101
rect 3787 -1135 3803 -1101
rect 3403 -1151 3803 -1135
rect 3975 -1101 4375 -1063
rect 3975 -1135 3991 -1101
rect 4359 -1135 4375 -1101
rect 3975 -1151 4375 -1135
rect 4547 -1101 4947 -1063
rect 4547 -1135 4563 -1101
rect 4931 -1135 4947 -1101
rect 4547 -1151 4947 -1135
rect 5119 -1101 5519 -1063
rect 5119 -1135 5135 -1101
rect 5503 -1135 5519 -1101
rect 5119 -1151 5519 -1135
rect -4605 -1209 -4205 -1193
rect -4605 -1243 -4589 -1209
rect -4221 -1243 -4205 -1209
rect -4605 -1281 -4205 -1243
rect -4033 -1209 -3633 -1193
rect -4033 -1243 -4017 -1209
rect -3649 -1243 -3633 -1209
rect -4033 -1281 -3633 -1243
rect -3461 -1209 -3061 -1193
rect -3461 -1243 -3445 -1209
rect -3077 -1243 -3061 -1209
rect -3461 -1281 -3061 -1243
rect -2889 -1209 -2489 -1193
rect -2889 -1243 -2873 -1209
rect -2505 -1243 -2489 -1209
rect -2889 -1281 -2489 -1243
rect -2317 -1209 -1917 -1193
rect -2317 -1243 -2301 -1209
rect -1933 -1243 -1917 -1209
rect -2317 -1281 -1917 -1243
rect -1745 -1209 -1345 -1193
rect -1745 -1243 -1729 -1209
rect -1361 -1243 -1345 -1209
rect -1745 -1281 -1345 -1243
rect -1173 -1209 -773 -1193
rect -1173 -1243 -1157 -1209
rect -789 -1243 -773 -1209
rect -1173 -1281 -773 -1243
rect -601 -1209 -201 -1193
rect -601 -1243 -585 -1209
rect -217 -1243 -201 -1209
rect -601 -1281 -201 -1243
rect -29 -1209 371 -1193
rect -29 -1243 -13 -1209
rect 355 -1243 371 -1209
rect -29 -1281 371 -1243
rect 543 -1209 943 -1193
rect 543 -1243 559 -1209
rect 927 -1243 943 -1209
rect 543 -1281 943 -1243
rect 1115 -1209 1515 -1193
rect 1115 -1243 1131 -1209
rect 1499 -1243 1515 -1209
rect 1115 -1281 1515 -1243
rect 1687 -1209 2087 -1193
rect 1687 -1243 1703 -1209
rect 2071 -1243 2087 -1209
rect 1687 -1281 2087 -1243
rect 2259 -1209 2659 -1193
rect 2259 -1243 2275 -1209
rect 2643 -1243 2659 -1209
rect 2259 -1281 2659 -1243
rect 2831 -1209 3231 -1193
rect 2831 -1243 2847 -1209
rect 3215 -1243 3231 -1209
rect 2831 -1281 3231 -1243
rect 3403 -1209 3803 -1193
rect 3403 -1243 3419 -1209
rect 3787 -1243 3803 -1209
rect 3403 -1281 3803 -1243
rect 3975 -1209 4375 -1193
rect 3975 -1243 3991 -1209
rect 4359 -1243 4375 -1209
rect 3975 -1281 4375 -1243
rect 4547 -1209 4947 -1193
rect 4547 -1243 4563 -1209
rect 4931 -1243 4947 -1209
rect 4547 -1281 4947 -1243
rect 5119 -1209 5519 -1193
rect 5119 -1243 5135 -1209
rect 5503 -1243 5519 -1209
rect 5119 -1281 5519 -1243
rect -4605 -2119 -4205 -2081
rect -4605 -2153 -4589 -2119
rect -4221 -2153 -4205 -2119
rect -4605 -2169 -4205 -2153
rect -4033 -2119 -3633 -2081
rect -4033 -2153 -4017 -2119
rect -3649 -2153 -3633 -2119
rect -4033 -2169 -3633 -2153
rect -3461 -2119 -3061 -2081
rect -3461 -2153 -3445 -2119
rect -3077 -2153 -3061 -2119
rect -3461 -2169 -3061 -2153
rect -2889 -2119 -2489 -2081
rect -2889 -2153 -2873 -2119
rect -2505 -2153 -2489 -2119
rect -2889 -2169 -2489 -2153
rect -2317 -2119 -1917 -2081
rect -2317 -2153 -2301 -2119
rect -1933 -2153 -1917 -2119
rect -2317 -2169 -1917 -2153
rect -1745 -2119 -1345 -2081
rect -1745 -2153 -1729 -2119
rect -1361 -2153 -1345 -2119
rect -1745 -2169 -1345 -2153
rect -1173 -2119 -773 -2081
rect -1173 -2153 -1157 -2119
rect -789 -2153 -773 -2119
rect -1173 -2169 -773 -2153
rect -601 -2119 -201 -2081
rect -601 -2153 -585 -2119
rect -217 -2153 -201 -2119
rect -601 -2169 -201 -2153
rect -29 -2119 371 -2081
rect -29 -2153 -13 -2119
rect 355 -2153 371 -2119
rect -29 -2169 371 -2153
rect 543 -2119 943 -2081
rect 543 -2153 559 -2119
rect 927 -2153 943 -2119
rect 543 -2169 943 -2153
rect 1115 -2119 1515 -2081
rect 1115 -2153 1131 -2119
rect 1499 -2153 1515 -2119
rect 1115 -2169 1515 -2153
rect 1687 -2119 2087 -2081
rect 1687 -2153 1703 -2119
rect 2071 -2153 2087 -2119
rect 1687 -2169 2087 -2153
rect 2259 -2119 2659 -2081
rect 2259 -2153 2275 -2119
rect 2643 -2153 2659 -2119
rect 2259 -2169 2659 -2153
rect 2831 -2119 3231 -2081
rect 2831 -2153 2847 -2119
rect 3215 -2153 3231 -2119
rect 2831 -2169 3231 -2153
rect 3403 -2119 3803 -2081
rect 3403 -2153 3419 -2119
rect 3787 -2153 3803 -2119
rect 3403 -2169 3803 -2153
rect 3975 -2119 4375 -2081
rect 3975 -2153 3991 -2119
rect 4359 -2153 4375 -2119
rect 3975 -2169 4375 -2153
rect 4547 -2119 4947 -2081
rect 4547 -2153 4563 -2119
rect 4931 -2153 4947 -2119
rect 4547 -2169 4947 -2153
rect 5119 -2119 5519 -2081
rect 5119 -2153 5135 -2119
rect 5503 -2153 5519 -2119
rect 5119 -2169 5519 -2153
rect -4605 -2227 -4205 -2211
rect -4605 -2261 -4589 -2227
rect -4221 -2261 -4205 -2227
rect -4605 -2299 -4205 -2261
rect -4033 -2227 -3633 -2211
rect -4033 -2261 -4017 -2227
rect -3649 -2261 -3633 -2227
rect -4033 -2299 -3633 -2261
rect -3461 -2227 -3061 -2211
rect -3461 -2261 -3445 -2227
rect -3077 -2261 -3061 -2227
rect -3461 -2299 -3061 -2261
rect -2889 -2227 -2489 -2211
rect -2889 -2261 -2873 -2227
rect -2505 -2261 -2489 -2227
rect -2889 -2299 -2489 -2261
rect -2317 -2227 -1917 -2211
rect -2317 -2261 -2301 -2227
rect -1933 -2261 -1917 -2227
rect -2317 -2299 -1917 -2261
rect -1745 -2227 -1345 -2211
rect -1745 -2261 -1729 -2227
rect -1361 -2261 -1345 -2227
rect -1745 -2299 -1345 -2261
rect -1173 -2227 -773 -2211
rect -1173 -2261 -1157 -2227
rect -789 -2261 -773 -2227
rect -1173 -2299 -773 -2261
rect -601 -2227 -201 -2211
rect -601 -2261 -585 -2227
rect -217 -2261 -201 -2227
rect -601 -2299 -201 -2261
rect -29 -2227 371 -2211
rect -29 -2261 -13 -2227
rect 355 -2261 371 -2227
rect -29 -2299 371 -2261
rect 543 -2227 943 -2211
rect 543 -2261 559 -2227
rect 927 -2261 943 -2227
rect 543 -2299 943 -2261
rect 1115 -2227 1515 -2211
rect 1115 -2261 1131 -2227
rect 1499 -2261 1515 -2227
rect 1115 -2299 1515 -2261
rect 1687 -2227 2087 -2211
rect 1687 -2261 1703 -2227
rect 2071 -2261 2087 -2227
rect 1687 -2299 2087 -2261
rect 2259 -2227 2659 -2211
rect 2259 -2261 2275 -2227
rect 2643 -2261 2659 -2227
rect 2259 -2299 2659 -2261
rect 2831 -2227 3231 -2211
rect 2831 -2261 2847 -2227
rect 3215 -2261 3231 -2227
rect 2831 -2299 3231 -2261
rect 3403 -2227 3803 -2211
rect 3403 -2261 3419 -2227
rect 3787 -2261 3803 -2227
rect 3403 -2299 3803 -2261
rect 3975 -2227 4375 -2211
rect 3975 -2261 3991 -2227
rect 4359 -2261 4375 -2227
rect 3975 -2299 4375 -2261
rect 4547 -2227 4947 -2211
rect 4547 -2261 4563 -2227
rect 4931 -2261 4947 -2227
rect 4547 -2299 4947 -2261
rect 5119 -2227 5519 -2211
rect 5119 -2261 5135 -2227
rect 5503 -2261 5519 -2227
rect 5119 -2299 5519 -2261
rect -4605 -3137 -4205 -3099
rect -4605 -3171 -4589 -3137
rect -4221 -3171 -4205 -3137
rect -4605 -3187 -4205 -3171
rect -4033 -3137 -3633 -3099
rect -4033 -3171 -4017 -3137
rect -3649 -3171 -3633 -3137
rect -4033 -3187 -3633 -3171
rect -3461 -3137 -3061 -3099
rect -3461 -3171 -3445 -3137
rect -3077 -3171 -3061 -3137
rect -3461 -3187 -3061 -3171
rect -2889 -3137 -2489 -3099
rect -2889 -3171 -2873 -3137
rect -2505 -3171 -2489 -3137
rect -2889 -3187 -2489 -3171
rect -2317 -3137 -1917 -3099
rect -2317 -3171 -2301 -3137
rect -1933 -3171 -1917 -3137
rect -2317 -3187 -1917 -3171
rect -1745 -3137 -1345 -3099
rect -1745 -3171 -1729 -3137
rect -1361 -3171 -1345 -3137
rect -1745 -3187 -1345 -3171
rect -1173 -3137 -773 -3099
rect -1173 -3171 -1157 -3137
rect -789 -3171 -773 -3137
rect -1173 -3187 -773 -3171
rect -601 -3137 -201 -3099
rect -601 -3171 -585 -3137
rect -217 -3171 -201 -3137
rect -601 -3187 -201 -3171
rect -29 -3137 371 -3099
rect -29 -3171 -13 -3137
rect 355 -3171 371 -3137
rect -29 -3187 371 -3171
rect 543 -3137 943 -3099
rect 543 -3171 559 -3137
rect 927 -3171 943 -3137
rect 543 -3187 943 -3171
rect 1115 -3137 1515 -3099
rect 1115 -3171 1131 -3137
rect 1499 -3171 1515 -3137
rect 1115 -3187 1515 -3171
rect 1687 -3137 2087 -3099
rect 1687 -3171 1703 -3137
rect 2071 -3171 2087 -3137
rect 1687 -3187 2087 -3171
rect 2259 -3137 2659 -3099
rect 2259 -3171 2275 -3137
rect 2643 -3171 2659 -3137
rect 2259 -3187 2659 -3171
rect 2831 -3137 3231 -3099
rect 2831 -3171 2847 -3137
rect 3215 -3171 3231 -3137
rect 2831 -3187 3231 -3171
rect 3403 -3137 3803 -3099
rect 3403 -3171 3419 -3137
rect 3787 -3171 3803 -3137
rect 3403 -3187 3803 -3171
rect 3975 -3137 4375 -3099
rect 3975 -3171 3991 -3137
rect 4359 -3171 4375 -3137
rect 3975 -3187 4375 -3171
rect 4547 -3137 4947 -3099
rect 4547 -3171 4563 -3137
rect 4931 -3171 4947 -3137
rect 4547 -3187 4947 -3171
rect 5119 -3137 5519 -3099
rect 5119 -3171 5135 -3137
rect 5503 -3171 5519 -3137
rect 5119 -3187 5519 -3171
<< polycont >>
rect -4589 793 -4221 827
rect -4017 793 -3649 827
rect -3445 793 -3077 827
rect -2873 793 -2505 827
rect -2301 793 -1933 827
rect -1729 793 -1361 827
rect -1157 793 -789 827
rect -585 793 -217 827
rect -13 793 355 827
rect 559 793 927 827
rect 1131 793 1499 827
rect 1703 793 2071 827
rect 2275 793 2643 827
rect 2847 793 3215 827
rect 3419 793 3787 827
rect 3991 793 4359 827
rect 4563 793 4931 827
rect 5135 793 5503 827
rect -4589 -117 -4221 -83
rect -4017 -117 -3649 -83
rect -3445 -117 -3077 -83
rect -2873 -117 -2505 -83
rect -2301 -117 -1933 -83
rect -1729 -117 -1361 -83
rect -1157 -117 -789 -83
rect -585 -117 -217 -83
rect -13 -117 355 -83
rect 559 -117 927 -83
rect 1131 -117 1499 -83
rect 1703 -117 2071 -83
rect 2275 -117 2643 -83
rect 2847 -117 3215 -83
rect 3419 -117 3787 -83
rect 3991 -117 4359 -83
rect 4563 -117 4931 -83
rect 5135 -117 5503 -83
rect -4589 -225 -4221 -191
rect -4017 -225 -3649 -191
rect -3445 -225 -3077 -191
rect -2873 -225 -2505 -191
rect -2301 -225 -1933 -191
rect -1729 -225 -1361 -191
rect -1157 -225 -789 -191
rect -585 -225 -217 -191
rect -13 -225 355 -191
rect 559 -225 927 -191
rect 1131 -225 1499 -191
rect 1703 -225 2071 -191
rect 2275 -225 2643 -191
rect 2847 -225 3215 -191
rect 3419 -225 3787 -191
rect 3991 -225 4359 -191
rect 4563 -225 4931 -191
rect 5135 -225 5503 -191
rect -4589 -1135 -4221 -1101
rect -4017 -1135 -3649 -1101
rect -3445 -1135 -3077 -1101
rect -2873 -1135 -2505 -1101
rect -2301 -1135 -1933 -1101
rect -1729 -1135 -1361 -1101
rect -1157 -1135 -789 -1101
rect -585 -1135 -217 -1101
rect -13 -1135 355 -1101
rect 559 -1135 927 -1101
rect 1131 -1135 1499 -1101
rect 1703 -1135 2071 -1101
rect 2275 -1135 2643 -1101
rect 2847 -1135 3215 -1101
rect 3419 -1135 3787 -1101
rect 3991 -1135 4359 -1101
rect 4563 -1135 4931 -1101
rect 5135 -1135 5503 -1101
rect -4589 -1243 -4221 -1209
rect -4017 -1243 -3649 -1209
rect -3445 -1243 -3077 -1209
rect -2873 -1243 -2505 -1209
rect -2301 -1243 -1933 -1209
rect -1729 -1243 -1361 -1209
rect -1157 -1243 -789 -1209
rect -585 -1243 -217 -1209
rect -13 -1243 355 -1209
rect 559 -1243 927 -1209
rect 1131 -1243 1499 -1209
rect 1703 -1243 2071 -1209
rect 2275 -1243 2643 -1209
rect 2847 -1243 3215 -1209
rect 3419 -1243 3787 -1209
rect 3991 -1243 4359 -1209
rect 4563 -1243 4931 -1209
rect 5135 -1243 5503 -1209
rect -4589 -2153 -4221 -2119
rect -4017 -2153 -3649 -2119
rect -3445 -2153 -3077 -2119
rect -2873 -2153 -2505 -2119
rect -2301 -2153 -1933 -2119
rect -1729 -2153 -1361 -2119
rect -1157 -2153 -789 -2119
rect -585 -2153 -217 -2119
rect -13 -2153 355 -2119
rect 559 -2153 927 -2119
rect 1131 -2153 1499 -2119
rect 1703 -2153 2071 -2119
rect 2275 -2153 2643 -2119
rect 2847 -2153 3215 -2119
rect 3419 -2153 3787 -2119
rect 3991 -2153 4359 -2119
rect 4563 -2153 4931 -2119
rect 5135 -2153 5503 -2119
rect -4589 -2261 -4221 -2227
rect -4017 -2261 -3649 -2227
rect -3445 -2261 -3077 -2227
rect -2873 -2261 -2505 -2227
rect -2301 -2261 -1933 -2227
rect -1729 -2261 -1361 -2227
rect -1157 -2261 -789 -2227
rect -585 -2261 -217 -2227
rect -13 -2261 355 -2227
rect 559 -2261 927 -2227
rect 1131 -2261 1499 -2227
rect 1703 -2261 2071 -2227
rect 2275 -2261 2643 -2227
rect 2847 -2261 3215 -2227
rect 3419 -2261 3787 -2227
rect 3991 -2261 4359 -2227
rect 4563 -2261 4931 -2227
rect 5135 -2261 5503 -2227
rect -4589 -3171 -4221 -3137
rect -4017 -3171 -3649 -3137
rect -3445 -3171 -3077 -3137
rect -2873 -3171 -2505 -3137
rect -2301 -3171 -1933 -3137
rect -1729 -3171 -1361 -3137
rect -1157 -3171 -789 -3137
rect -585 -3171 -217 -3137
rect -13 -3171 355 -3137
rect 559 -3171 927 -3137
rect 1131 -3171 1499 -3137
rect 1703 -3171 2071 -3137
rect 2275 -3171 2643 -3137
rect 2847 -3171 3215 -3137
rect 3419 -3171 3787 -3137
rect 3991 -3171 4359 -3137
rect 4563 -3171 4931 -3137
rect 5135 -3171 5503 -3137
<< locali >>
rect -4765 895 -4669 929
rect 5583 895 5679 929
rect -4765 833 -4731 895
rect 5645 833 5679 895
rect -4605 793 -4589 827
rect -4221 793 -4205 827
rect -4033 793 -4017 827
rect -3649 793 -3633 827
rect -3461 793 -3445 827
rect -3077 793 -3061 827
rect -2889 793 -2873 827
rect -2505 793 -2489 827
rect -2317 793 -2301 827
rect -1933 793 -1917 827
rect -1745 793 -1729 827
rect -1361 793 -1345 827
rect -1173 793 -1157 827
rect -789 793 -773 827
rect -601 793 -585 827
rect -217 793 -201 827
rect -29 793 -13 827
rect 355 793 371 827
rect 543 793 559 827
rect 927 793 943 827
rect 1115 793 1131 827
rect 1499 793 1515 827
rect 1687 793 1703 827
rect 2071 793 2087 827
rect 2259 793 2275 827
rect 2643 793 2659 827
rect 2831 793 2847 827
rect 3215 793 3231 827
rect 3403 793 3419 827
rect 3787 793 3803 827
rect 3975 793 3991 827
rect 4359 793 4375 827
rect 4547 793 4563 827
rect 4931 793 4947 827
rect 5119 793 5135 827
rect 5503 793 5519 827
rect -4651 743 -4617 759
rect -4651 -49 -4617 -33
rect -4193 743 -4159 759
rect -4193 -49 -4159 -33
rect -4079 743 -4045 759
rect -4079 -49 -4045 -33
rect -3621 743 -3587 759
rect -3621 -49 -3587 -33
rect -3507 743 -3473 759
rect -3507 -49 -3473 -33
rect -3049 743 -3015 759
rect -3049 -49 -3015 -33
rect -2935 743 -2901 759
rect -2935 -49 -2901 -33
rect -2477 743 -2443 759
rect -2477 -49 -2443 -33
rect -2363 743 -2329 759
rect -2363 -49 -2329 -33
rect -1905 743 -1871 759
rect -1905 -49 -1871 -33
rect -1791 743 -1757 759
rect -1791 -49 -1757 -33
rect -1333 743 -1299 759
rect -1333 -49 -1299 -33
rect -1219 743 -1185 759
rect -1219 -49 -1185 -33
rect -761 743 -727 759
rect -761 -49 -727 -33
rect -647 743 -613 759
rect -647 -49 -613 -33
rect -189 743 -155 759
rect -189 -49 -155 -33
rect -75 743 -41 759
rect -75 -49 -41 -33
rect 383 743 417 759
rect 383 -49 417 -33
rect 497 743 531 759
rect 497 -49 531 -33
rect 955 743 989 759
rect 955 -49 989 -33
rect 1069 743 1103 759
rect 1069 -49 1103 -33
rect 1527 743 1561 759
rect 1527 -49 1561 -33
rect 1641 743 1675 759
rect 1641 -49 1675 -33
rect 2099 743 2133 759
rect 2099 -49 2133 -33
rect 2213 743 2247 759
rect 2213 -49 2247 -33
rect 2671 743 2705 759
rect 2671 -49 2705 -33
rect 2785 743 2819 759
rect 2785 -49 2819 -33
rect 3243 743 3277 759
rect 3243 -49 3277 -33
rect 3357 743 3391 759
rect 3357 -49 3391 -33
rect 3815 743 3849 759
rect 3815 -49 3849 -33
rect 3929 743 3963 759
rect 3929 -49 3963 -33
rect 4387 743 4421 759
rect 4387 -49 4421 -33
rect 4501 743 4535 759
rect 4501 -49 4535 -33
rect 4959 743 4993 759
rect 4959 -49 4993 -33
rect 5073 743 5107 759
rect 5073 -49 5107 -33
rect 5531 743 5565 759
rect 5531 -49 5565 -33
rect -4605 -117 -4589 -83
rect -4221 -117 -4205 -83
rect -4033 -117 -4017 -83
rect -3649 -117 -3633 -83
rect -3461 -117 -3445 -83
rect -3077 -117 -3061 -83
rect -2889 -117 -2873 -83
rect -2505 -117 -2489 -83
rect -2317 -117 -2301 -83
rect -1933 -117 -1917 -83
rect -1745 -117 -1729 -83
rect -1361 -117 -1345 -83
rect -1173 -117 -1157 -83
rect -789 -117 -773 -83
rect -601 -117 -585 -83
rect -217 -117 -201 -83
rect -29 -117 -13 -83
rect 355 -117 371 -83
rect 543 -117 559 -83
rect 927 -117 943 -83
rect 1115 -117 1131 -83
rect 1499 -117 1515 -83
rect 1687 -117 1703 -83
rect 2071 -117 2087 -83
rect 2259 -117 2275 -83
rect 2643 -117 2659 -83
rect 2831 -117 2847 -83
rect 3215 -117 3231 -83
rect 3403 -117 3419 -83
rect 3787 -117 3803 -83
rect 3975 -117 3991 -83
rect 4359 -117 4375 -83
rect 4547 -117 4563 -83
rect 4931 -117 4947 -83
rect 5119 -117 5135 -83
rect 5503 -117 5519 -83
rect -4605 -225 -4589 -191
rect -4221 -225 -4205 -191
rect -4033 -225 -4017 -191
rect -3649 -225 -3633 -191
rect -3461 -225 -3445 -191
rect -3077 -225 -3061 -191
rect -2889 -225 -2873 -191
rect -2505 -225 -2489 -191
rect -2317 -225 -2301 -191
rect -1933 -225 -1917 -191
rect -1745 -225 -1729 -191
rect -1361 -225 -1345 -191
rect -1173 -225 -1157 -191
rect -789 -225 -773 -191
rect -601 -225 -585 -191
rect -217 -225 -201 -191
rect -29 -225 -13 -191
rect 355 -225 371 -191
rect 543 -225 559 -191
rect 927 -225 943 -191
rect 1115 -225 1131 -191
rect 1499 -225 1515 -191
rect 1687 -225 1703 -191
rect 2071 -225 2087 -191
rect 2259 -225 2275 -191
rect 2643 -225 2659 -191
rect 2831 -225 2847 -191
rect 3215 -225 3231 -191
rect 3403 -225 3419 -191
rect 3787 -225 3803 -191
rect 3975 -225 3991 -191
rect 4359 -225 4375 -191
rect 4547 -225 4563 -191
rect 4931 -225 4947 -191
rect 5119 -225 5135 -191
rect 5503 -225 5519 -191
rect -4651 -275 -4617 -259
rect -4651 -1067 -4617 -1051
rect -4193 -275 -4159 -259
rect -4193 -1067 -4159 -1051
rect -4079 -275 -4045 -259
rect -4079 -1067 -4045 -1051
rect -3621 -275 -3587 -259
rect -3621 -1067 -3587 -1051
rect -3507 -275 -3473 -259
rect -3507 -1067 -3473 -1051
rect -3049 -275 -3015 -259
rect -3049 -1067 -3015 -1051
rect -2935 -275 -2901 -259
rect -2935 -1067 -2901 -1051
rect -2477 -275 -2443 -259
rect -2477 -1067 -2443 -1051
rect -2363 -275 -2329 -259
rect -2363 -1067 -2329 -1051
rect -1905 -275 -1871 -259
rect -1905 -1067 -1871 -1051
rect -1791 -275 -1757 -259
rect -1791 -1067 -1757 -1051
rect -1333 -275 -1299 -259
rect -1333 -1067 -1299 -1051
rect -1219 -275 -1185 -259
rect -1219 -1067 -1185 -1051
rect -761 -275 -727 -259
rect -761 -1067 -727 -1051
rect -647 -275 -613 -259
rect -647 -1067 -613 -1051
rect -189 -275 -155 -259
rect -189 -1067 -155 -1051
rect -75 -275 -41 -259
rect -75 -1067 -41 -1051
rect 383 -275 417 -259
rect 383 -1067 417 -1051
rect 497 -275 531 -259
rect 497 -1067 531 -1051
rect 955 -275 989 -259
rect 955 -1067 989 -1051
rect 1069 -275 1103 -259
rect 1069 -1067 1103 -1051
rect 1527 -275 1561 -259
rect 1527 -1067 1561 -1051
rect 1641 -275 1675 -259
rect 1641 -1067 1675 -1051
rect 2099 -275 2133 -259
rect 2099 -1067 2133 -1051
rect 2213 -275 2247 -259
rect 2213 -1067 2247 -1051
rect 2671 -275 2705 -259
rect 2671 -1067 2705 -1051
rect 2785 -275 2819 -259
rect 2785 -1067 2819 -1051
rect 3243 -275 3277 -259
rect 3243 -1067 3277 -1051
rect 3357 -275 3391 -259
rect 3357 -1067 3391 -1051
rect 3815 -275 3849 -259
rect 3815 -1067 3849 -1051
rect 3929 -275 3963 -259
rect 3929 -1067 3963 -1051
rect 4387 -275 4421 -259
rect 4387 -1067 4421 -1051
rect 4501 -275 4535 -259
rect 4501 -1067 4535 -1051
rect 4959 -275 4993 -259
rect 4959 -1067 4993 -1051
rect 5073 -275 5107 -259
rect 5073 -1067 5107 -1051
rect 5531 -275 5565 -259
rect 5531 -1067 5565 -1051
rect -4605 -1135 -4589 -1101
rect -4221 -1135 -4205 -1101
rect -4033 -1135 -4017 -1101
rect -3649 -1135 -3633 -1101
rect -3461 -1135 -3445 -1101
rect -3077 -1135 -3061 -1101
rect -2889 -1135 -2873 -1101
rect -2505 -1135 -2489 -1101
rect -2317 -1135 -2301 -1101
rect -1933 -1135 -1917 -1101
rect -1745 -1135 -1729 -1101
rect -1361 -1135 -1345 -1101
rect -1173 -1135 -1157 -1101
rect -789 -1135 -773 -1101
rect -601 -1135 -585 -1101
rect -217 -1135 -201 -1101
rect -29 -1135 -13 -1101
rect 355 -1135 371 -1101
rect 543 -1135 559 -1101
rect 927 -1135 943 -1101
rect 1115 -1135 1131 -1101
rect 1499 -1135 1515 -1101
rect 1687 -1135 1703 -1101
rect 2071 -1135 2087 -1101
rect 2259 -1135 2275 -1101
rect 2643 -1135 2659 -1101
rect 2831 -1135 2847 -1101
rect 3215 -1135 3231 -1101
rect 3403 -1135 3419 -1101
rect 3787 -1135 3803 -1101
rect 3975 -1135 3991 -1101
rect 4359 -1135 4375 -1101
rect 4547 -1135 4563 -1101
rect 4931 -1135 4947 -1101
rect 5119 -1135 5135 -1101
rect 5503 -1135 5519 -1101
rect -4605 -1243 -4589 -1209
rect -4221 -1243 -4205 -1209
rect -4033 -1243 -4017 -1209
rect -3649 -1243 -3633 -1209
rect -3461 -1243 -3445 -1209
rect -3077 -1243 -3061 -1209
rect -2889 -1243 -2873 -1209
rect -2505 -1243 -2489 -1209
rect -2317 -1243 -2301 -1209
rect -1933 -1243 -1917 -1209
rect -1745 -1243 -1729 -1209
rect -1361 -1243 -1345 -1209
rect -1173 -1243 -1157 -1209
rect -789 -1243 -773 -1209
rect -601 -1243 -585 -1209
rect -217 -1243 -201 -1209
rect -29 -1243 -13 -1209
rect 355 -1243 371 -1209
rect 543 -1243 559 -1209
rect 927 -1243 943 -1209
rect 1115 -1243 1131 -1209
rect 1499 -1243 1515 -1209
rect 1687 -1243 1703 -1209
rect 2071 -1243 2087 -1209
rect 2259 -1243 2275 -1209
rect 2643 -1243 2659 -1209
rect 2831 -1243 2847 -1209
rect 3215 -1243 3231 -1209
rect 3403 -1243 3419 -1209
rect 3787 -1243 3803 -1209
rect 3975 -1243 3991 -1209
rect 4359 -1243 4375 -1209
rect 4547 -1243 4563 -1209
rect 4931 -1243 4947 -1209
rect 5119 -1243 5135 -1209
rect 5503 -1243 5519 -1209
rect -4651 -1293 -4617 -1277
rect -4651 -2085 -4617 -2069
rect -4193 -1293 -4159 -1277
rect -4193 -2085 -4159 -2069
rect -4079 -1293 -4045 -1277
rect -4079 -2085 -4045 -2069
rect -3621 -1293 -3587 -1277
rect -3621 -2085 -3587 -2069
rect -3507 -1293 -3473 -1277
rect -3507 -2085 -3473 -2069
rect -3049 -1293 -3015 -1277
rect -3049 -2085 -3015 -2069
rect -2935 -1293 -2901 -1277
rect -2935 -2085 -2901 -2069
rect -2477 -1293 -2443 -1277
rect -2477 -2085 -2443 -2069
rect -2363 -1293 -2329 -1277
rect -2363 -2085 -2329 -2069
rect -1905 -1293 -1871 -1277
rect -1905 -2085 -1871 -2069
rect -1791 -1293 -1757 -1277
rect -1791 -2085 -1757 -2069
rect -1333 -1293 -1299 -1277
rect -1333 -2085 -1299 -2069
rect -1219 -1293 -1185 -1277
rect -1219 -2085 -1185 -2069
rect -761 -1293 -727 -1277
rect -761 -2085 -727 -2069
rect -647 -1293 -613 -1277
rect -647 -2085 -613 -2069
rect -189 -1293 -155 -1277
rect -189 -2085 -155 -2069
rect -75 -1293 -41 -1277
rect -75 -2085 -41 -2069
rect 383 -1293 417 -1277
rect 383 -2085 417 -2069
rect 497 -1293 531 -1277
rect 497 -2085 531 -2069
rect 955 -1293 989 -1277
rect 955 -2085 989 -2069
rect 1069 -1293 1103 -1277
rect 1069 -2085 1103 -2069
rect 1527 -1293 1561 -1277
rect 1527 -2085 1561 -2069
rect 1641 -1293 1675 -1277
rect 1641 -2085 1675 -2069
rect 2099 -1293 2133 -1277
rect 2099 -2085 2133 -2069
rect 2213 -1293 2247 -1277
rect 2213 -2085 2247 -2069
rect 2671 -1293 2705 -1277
rect 2671 -2085 2705 -2069
rect 2785 -1293 2819 -1277
rect 2785 -2085 2819 -2069
rect 3243 -1293 3277 -1277
rect 3243 -2085 3277 -2069
rect 3357 -1293 3391 -1277
rect 3357 -2085 3391 -2069
rect 3815 -1293 3849 -1277
rect 3815 -2085 3849 -2069
rect 3929 -1293 3963 -1277
rect 3929 -2085 3963 -2069
rect 4387 -1293 4421 -1277
rect 4387 -2085 4421 -2069
rect 4501 -1293 4535 -1277
rect 4501 -2085 4535 -2069
rect 4959 -1293 4993 -1277
rect 4959 -2085 4993 -2069
rect 5073 -1293 5107 -1277
rect 5073 -2085 5107 -2069
rect 5531 -1293 5565 -1277
rect 5531 -2085 5565 -2069
rect -4605 -2153 -4589 -2119
rect -4221 -2153 -4205 -2119
rect -4033 -2153 -4017 -2119
rect -3649 -2153 -3633 -2119
rect -3461 -2153 -3445 -2119
rect -3077 -2153 -3061 -2119
rect -2889 -2153 -2873 -2119
rect -2505 -2153 -2489 -2119
rect -2317 -2153 -2301 -2119
rect -1933 -2153 -1917 -2119
rect -1745 -2153 -1729 -2119
rect -1361 -2153 -1345 -2119
rect -1173 -2153 -1157 -2119
rect -789 -2153 -773 -2119
rect -601 -2153 -585 -2119
rect -217 -2153 -201 -2119
rect -29 -2153 -13 -2119
rect 355 -2153 371 -2119
rect 543 -2153 559 -2119
rect 927 -2153 943 -2119
rect 1115 -2153 1131 -2119
rect 1499 -2153 1515 -2119
rect 1687 -2153 1703 -2119
rect 2071 -2153 2087 -2119
rect 2259 -2153 2275 -2119
rect 2643 -2153 2659 -2119
rect 2831 -2153 2847 -2119
rect 3215 -2153 3231 -2119
rect 3403 -2153 3419 -2119
rect 3787 -2153 3803 -2119
rect 3975 -2153 3991 -2119
rect 4359 -2153 4375 -2119
rect 4547 -2153 4563 -2119
rect 4931 -2153 4947 -2119
rect 5119 -2153 5135 -2119
rect 5503 -2153 5519 -2119
rect -4605 -2261 -4589 -2227
rect -4221 -2261 -4205 -2227
rect -4033 -2261 -4017 -2227
rect -3649 -2261 -3633 -2227
rect -3461 -2261 -3445 -2227
rect -3077 -2261 -3061 -2227
rect -2889 -2261 -2873 -2227
rect -2505 -2261 -2489 -2227
rect -2317 -2261 -2301 -2227
rect -1933 -2261 -1917 -2227
rect -1745 -2261 -1729 -2227
rect -1361 -2261 -1345 -2227
rect -1173 -2261 -1157 -2227
rect -789 -2261 -773 -2227
rect -601 -2261 -585 -2227
rect -217 -2261 -201 -2227
rect -29 -2261 -13 -2227
rect 355 -2261 371 -2227
rect 543 -2261 559 -2227
rect 927 -2261 943 -2227
rect 1115 -2261 1131 -2227
rect 1499 -2261 1515 -2227
rect 1687 -2261 1703 -2227
rect 2071 -2261 2087 -2227
rect 2259 -2261 2275 -2227
rect 2643 -2261 2659 -2227
rect 2831 -2261 2847 -2227
rect 3215 -2261 3231 -2227
rect 3403 -2261 3419 -2227
rect 3787 -2261 3803 -2227
rect 3975 -2261 3991 -2227
rect 4359 -2261 4375 -2227
rect 4547 -2261 4563 -2227
rect 4931 -2261 4947 -2227
rect 5119 -2261 5135 -2227
rect 5503 -2261 5519 -2227
rect -4651 -2311 -4617 -2295
rect -4651 -3103 -4617 -3087
rect -4193 -2311 -4159 -2295
rect -4193 -3103 -4159 -3087
rect -4079 -2311 -4045 -2295
rect -4079 -3103 -4045 -3087
rect -3621 -2311 -3587 -2295
rect -3621 -3103 -3587 -3087
rect -3507 -2311 -3473 -2295
rect -3507 -3103 -3473 -3087
rect -3049 -2311 -3015 -2295
rect -3049 -3103 -3015 -3087
rect -2935 -2311 -2901 -2295
rect -2935 -3103 -2901 -3087
rect -2477 -2311 -2443 -2295
rect -2477 -3103 -2443 -3087
rect -2363 -2311 -2329 -2295
rect -2363 -3103 -2329 -3087
rect -1905 -2311 -1871 -2295
rect -1905 -3103 -1871 -3087
rect -1791 -2311 -1757 -2295
rect -1791 -3103 -1757 -3087
rect -1333 -2311 -1299 -2295
rect -1333 -3103 -1299 -3087
rect -1219 -2311 -1185 -2295
rect -1219 -3103 -1185 -3087
rect -761 -2311 -727 -2295
rect -761 -3103 -727 -3087
rect -647 -2311 -613 -2295
rect -647 -3103 -613 -3087
rect -189 -2311 -155 -2295
rect -189 -3103 -155 -3087
rect -75 -2311 -41 -2295
rect -75 -3103 -41 -3087
rect 383 -2311 417 -2295
rect 383 -3103 417 -3087
rect 497 -2311 531 -2295
rect 497 -3103 531 -3087
rect 955 -2311 989 -2295
rect 955 -3103 989 -3087
rect 1069 -2311 1103 -2295
rect 1069 -3103 1103 -3087
rect 1527 -2311 1561 -2295
rect 1527 -3103 1561 -3087
rect 1641 -2311 1675 -2295
rect 1641 -3103 1675 -3087
rect 2099 -2311 2133 -2295
rect 2099 -3103 2133 -3087
rect 2213 -2311 2247 -2295
rect 2213 -3103 2247 -3087
rect 2671 -2311 2705 -2295
rect 2671 -3103 2705 -3087
rect 2785 -2311 2819 -2295
rect 2785 -3103 2819 -3087
rect 3243 -2311 3277 -2295
rect 3243 -3103 3277 -3087
rect 3357 -2311 3391 -2295
rect 3357 -3103 3391 -3087
rect 3815 -2311 3849 -2295
rect 3815 -3103 3849 -3087
rect 3929 -2311 3963 -2295
rect 3929 -3103 3963 -3087
rect 4387 -2311 4421 -2295
rect 4387 -3103 4421 -3087
rect 4501 -2311 4535 -2295
rect 4501 -3103 4535 -3087
rect 4959 -2311 4993 -2295
rect 4959 -3103 4993 -3087
rect 5073 -2311 5107 -2295
rect 5073 -3103 5107 -3087
rect 5531 -2311 5565 -2295
rect 5531 -3103 5565 -3087
rect -4605 -3171 -4589 -3137
rect -4221 -3171 -4205 -3137
rect -4033 -3171 -4017 -3137
rect -3649 -3171 -3633 -3137
rect -3461 -3171 -3445 -3137
rect -3077 -3171 -3061 -3137
rect -2889 -3171 -2873 -3137
rect -2505 -3171 -2489 -3137
rect -2317 -3171 -2301 -3137
rect -1933 -3171 -1917 -3137
rect -1745 -3171 -1729 -3137
rect -1361 -3171 -1345 -3137
rect -1173 -3171 -1157 -3137
rect -789 -3171 -773 -3137
rect -601 -3171 -585 -3137
rect -217 -3171 -201 -3137
rect -29 -3171 -13 -3137
rect 355 -3171 371 -3137
rect 543 -3171 559 -3137
rect 927 -3171 943 -3137
rect 1115 -3171 1131 -3137
rect 1499 -3171 1515 -3137
rect 1687 -3171 1703 -3137
rect 2071 -3171 2087 -3137
rect 2259 -3171 2275 -3137
rect 2643 -3171 2659 -3137
rect 2831 -3171 2847 -3137
rect 3215 -3171 3231 -3137
rect 3403 -3171 3419 -3137
rect 3787 -3171 3803 -3137
rect 3975 -3171 3991 -3137
rect 4359 -3171 4375 -3137
rect 4547 -3171 4563 -3137
rect 4931 -3171 4947 -3137
rect 5119 -3171 5135 -3137
rect 5503 -3171 5519 -3137
rect -4765 -3239 -4731 -3177
rect 5645 -3239 5679 -3177
rect -4765 -3273 -4669 -3239
rect 5598 -3273 5679 -3239
<< viali >>
rect -4589 793 -4221 827
rect -4017 793 -3649 827
rect -3445 793 -3077 827
rect -2873 793 -2505 827
rect -2301 793 -1933 827
rect -1729 793 -1361 827
rect -1157 793 -789 827
rect -585 793 -217 827
rect -13 793 355 827
rect 559 793 927 827
rect 1131 793 1499 827
rect 1703 793 2071 827
rect 2275 793 2643 827
rect 2847 793 3215 827
rect 3419 793 3787 827
rect 3991 793 4359 827
rect 4563 793 4931 827
rect 5135 793 5503 827
rect -4651 -33 -4617 743
rect -4193 -33 -4159 743
rect -4079 -33 -4045 743
rect -3621 -33 -3587 743
rect -3507 -33 -3473 743
rect -3049 -33 -3015 743
rect -2935 -33 -2901 743
rect -2477 -33 -2443 743
rect -2363 -33 -2329 743
rect -1905 -33 -1871 743
rect -1791 -33 -1757 743
rect -1333 -33 -1299 743
rect -1219 -33 -1185 743
rect -761 -33 -727 743
rect -647 -33 -613 743
rect -189 -33 -155 743
rect -75 -33 -41 743
rect 383 -33 417 743
rect 497 -33 531 743
rect 955 -33 989 743
rect 1069 -33 1103 743
rect 1527 -33 1561 743
rect 1641 -33 1675 743
rect 2099 -33 2133 743
rect 2213 -33 2247 743
rect 2671 -33 2705 743
rect 2785 -33 2819 743
rect 3243 -33 3277 743
rect 3357 -33 3391 743
rect 3815 -33 3849 743
rect 3929 -33 3963 743
rect 4387 -33 4421 743
rect 4501 -33 4535 743
rect 4959 -33 4993 743
rect 5073 -33 5107 743
rect 5531 -33 5565 743
rect -4589 -117 -4221 -83
rect -4017 -117 -3649 -83
rect -3445 -117 -3077 -83
rect -2873 -117 -2505 -83
rect -2301 -117 -1933 -83
rect -1729 -117 -1361 -83
rect -1157 -117 -789 -83
rect -585 -117 -217 -83
rect -13 -117 355 -83
rect 559 -117 927 -83
rect 1131 -117 1499 -83
rect 1703 -117 2071 -83
rect 2275 -117 2643 -83
rect 2847 -117 3215 -83
rect 3419 -117 3787 -83
rect 3991 -117 4359 -83
rect 4563 -117 4931 -83
rect 5135 -117 5503 -83
rect -4589 -225 -4221 -191
rect -4017 -225 -3649 -191
rect -3445 -225 -3077 -191
rect -2873 -225 -2505 -191
rect -2301 -225 -1933 -191
rect -1729 -225 -1361 -191
rect -1157 -225 -789 -191
rect -585 -225 -217 -191
rect -13 -225 355 -191
rect 559 -225 927 -191
rect 1131 -225 1499 -191
rect 1703 -225 2071 -191
rect 2275 -225 2643 -191
rect 2847 -225 3215 -191
rect 3419 -225 3787 -191
rect 3991 -225 4359 -191
rect 4563 -225 4931 -191
rect 5135 -225 5503 -191
rect -4651 -1051 -4617 -275
rect -4193 -1051 -4159 -275
rect -4079 -1051 -4045 -275
rect -3621 -1051 -3587 -275
rect -3507 -1051 -3473 -275
rect -3049 -1051 -3015 -275
rect -2935 -1051 -2901 -275
rect -2477 -1051 -2443 -275
rect -2363 -1051 -2329 -275
rect -1905 -1051 -1871 -275
rect -1791 -1051 -1757 -275
rect -1333 -1051 -1299 -275
rect -1219 -1051 -1185 -275
rect -761 -1051 -727 -275
rect -647 -1051 -613 -275
rect -189 -1051 -155 -275
rect -75 -1051 -41 -275
rect 383 -1051 417 -275
rect 497 -1051 531 -275
rect 955 -1051 989 -275
rect 1069 -1051 1103 -275
rect 1527 -1051 1561 -275
rect 1641 -1051 1675 -275
rect 2099 -1051 2133 -275
rect 2213 -1051 2247 -275
rect 2671 -1051 2705 -275
rect 2785 -1051 2819 -275
rect 3243 -1051 3277 -275
rect 3357 -1051 3391 -275
rect 3815 -1051 3849 -275
rect 3929 -1051 3963 -275
rect 4387 -1051 4421 -275
rect 4501 -1051 4535 -275
rect 4959 -1051 4993 -275
rect 5073 -1051 5107 -275
rect 5531 -1051 5565 -275
rect -4589 -1135 -4221 -1101
rect -4017 -1135 -3649 -1101
rect -3445 -1135 -3077 -1101
rect -2873 -1135 -2505 -1101
rect -2301 -1135 -1933 -1101
rect -1729 -1135 -1361 -1101
rect -1157 -1135 -789 -1101
rect -585 -1135 -217 -1101
rect -13 -1135 355 -1101
rect 559 -1135 927 -1101
rect 1131 -1135 1499 -1101
rect 1703 -1135 2071 -1101
rect 2275 -1135 2643 -1101
rect 2847 -1135 3215 -1101
rect 3419 -1135 3787 -1101
rect 3991 -1135 4359 -1101
rect 4563 -1135 4931 -1101
rect 5135 -1135 5503 -1101
rect -4589 -1243 -4221 -1209
rect -4017 -1243 -3649 -1209
rect -3445 -1243 -3077 -1209
rect -2873 -1243 -2505 -1209
rect -2301 -1243 -1933 -1209
rect -1729 -1243 -1361 -1209
rect -1157 -1243 -789 -1209
rect -585 -1243 -217 -1209
rect -13 -1243 355 -1209
rect 559 -1243 927 -1209
rect 1131 -1243 1499 -1209
rect 1703 -1243 2071 -1209
rect 2275 -1243 2643 -1209
rect 2847 -1243 3215 -1209
rect 3419 -1243 3787 -1209
rect 3991 -1243 4359 -1209
rect 4563 -1243 4931 -1209
rect 5135 -1243 5503 -1209
rect -4651 -2069 -4617 -1293
rect -4193 -2069 -4159 -1293
rect -4079 -2069 -4045 -1293
rect -3621 -2069 -3587 -1293
rect -3507 -2069 -3473 -1293
rect -3049 -2069 -3015 -1293
rect -2935 -2069 -2901 -1293
rect -2477 -2069 -2443 -1293
rect -2363 -2069 -2329 -1293
rect -1905 -2069 -1871 -1293
rect -1791 -2069 -1757 -1293
rect -1333 -2069 -1299 -1293
rect -1219 -2069 -1185 -1293
rect -761 -2069 -727 -1293
rect -647 -2069 -613 -1293
rect -189 -2069 -155 -1293
rect -75 -2069 -41 -1293
rect 383 -2069 417 -1293
rect 497 -2069 531 -1293
rect 955 -2069 989 -1293
rect 1069 -2069 1103 -1293
rect 1527 -2069 1561 -1293
rect 1641 -2069 1675 -1293
rect 2099 -2069 2133 -1293
rect 2213 -2069 2247 -1293
rect 2671 -2069 2705 -1293
rect 2785 -2069 2819 -1293
rect 3243 -2069 3277 -1293
rect 3357 -2069 3391 -1293
rect 3815 -2069 3849 -1293
rect 3929 -2069 3963 -1293
rect 4387 -2069 4421 -1293
rect 4501 -2069 4535 -1293
rect 4959 -2069 4993 -1293
rect 5073 -2069 5107 -1293
rect 5531 -2069 5565 -1293
rect -4589 -2153 -4221 -2119
rect -4017 -2153 -3649 -2119
rect -3445 -2153 -3077 -2119
rect -2873 -2153 -2505 -2119
rect -2301 -2153 -1933 -2119
rect -1729 -2153 -1361 -2119
rect -1157 -2153 -789 -2119
rect -585 -2153 -217 -2119
rect -13 -2153 355 -2119
rect 559 -2153 927 -2119
rect 1131 -2153 1499 -2119
rect 1703 -2153 2071 -2119
rect 2275 -2153 2643 -2119
rect 2847 -2153 3215 -2119
rect 3419 -2153 3787 -2119
rect 3991 -2153 4359 -2119
rect 4563 -2153 4931 -2119
rect 5135 -2153 5503 -2119
rect -4589 -2261 -4221 -2227
rect -4017 -2261 -3649 -2227
rect -3445 -2261 -3077 -2227
rect -2873 -2261 -2505 -2227
rect -2301 -2261 -1933 -2227
rect -1729 -2261 -1361 -2227
rect -1157 -2261 -789 -2227
rect -585 -2261 -217 -2227
rect -13 -2261 355 -2227
rect 559 -2261 927 -2227
rect 1131 -2261 1499 -2227
rect 1703 -2261 2071 -2227
rect 2275 -2261 2643 -2227
rect 2847 -2261 3215 -2227
rect 3419 -2261 3787 -2227
rect 3991 -2261 4359 -2227
rect 4563 -2261 4931 -2227
rect 5135 -2261 5503 -2227
rect -4651 -3087 -4617 -2311
rect -4193 -3087 -4159 -2311
rect -4079 -3087 -4045 -2311
rect -3621 -3087 -3587 -2311
rect -3507 -3087 -3473 -2311
rect -3049 -3087 -3015 -2311
rect -2935 -3087 -2901 -2311
rect -2477 -3087 -2443 -2311
rect -2363 -3087 -2329 -2311
rect -1905 -3087 -1871 -2311
rect -1791 -3087 -1757 -2311
rect -1333 -3087 -1299 -2311
rect -1219 -3087 -1185 -2311
rect -761 -3087 -727 -2311
rect -647 -3087 -613 -2311
rect -189 -3087 -155 -2311
rect -75 -3087 -41 -2311
rect 383 -3087 417 -2311
rect 497 -3087 531 -2311
rect 955 -3087 989 -2311
rect 1069 -3087 1103 -2311
rect 1527 -3087 1561 -2311
rect 1641 -3087 1675 -2311
rect 2099 -3087 2133 -2311
rect 2213 -3087 2247 -2311
rect 2671 -3087 2705 -2311
rect 2785 -3087 2819 -2311
rect 3243 -3087 3277 -2311
rect 3357 -3087 3391 -2311
rect 3815 -3087 3849 -2311
rect 3929 -3087 3963 -2311
rect 4387 -3087 4421 -2311
rect 4501 -3087 4535 -2311
rect 4959 -3087 4993 -2311
rect 5073 -3087 5107 -2311
rect 5531 -3087 5565 -2311
rect -4589 -3171 -4221 -3137
rect -4017 -3171 -3649 -3137
rect -3445 -3171 -3077 -3137
rect -2873 -3171 -2505 -3137
rect -2301 -3171 -1933 -3137
rect -1729 -3171 -1361 -3137
rect -1157 -3171 -789 -3137
rect -585 -3171 -217 -3137
rect -13 -3171 355 -3137
rect 559 -3171 927 -3137
rect 1131 -3171 1499 -3137
rect 1703 -3171 2071 -3137
rect 2275 -3171 2643 -3137
rect 2847 -3171 3215 -3137
rect 3419 -3171 3787 -3137
rect 3991 -3171 4359 -3137
rect 4563 -3171 4931 -3137
rect 5135 -3171 5503 -3137
rect -4664 -3239 -4592 -3218
rect -3582 -3239 -3510 -3218
rect -2438 -3239 -2366 -3218
rect -1294 -3239 -1222 -3218
rect -150 -3239 -78 -3218
rect 994 -3239 1066 -3218
rect 2138 -3239 2210 -3218
rect 3282 -3239 3354 -3218
rect 4426 -3239 4498 -3218
rect 5526 -3239 5598 -3218
rect -4664 -3273 -4592 -3239
rect -3582 -3273 -3510 -3239
rect -2438 -3273 -2366 -3239
rect -1294 -3273 -1222 -3239
rect -150 -3273 -78 -3239
rect 994 -3273 1066 -3239
rect 2138 -3273 2210 -3239
rect 3282 -3273 3354 -3239
rect 4426 -3273 4498 -3239
rect 5526 -3273 5583 -3239
rect 5583 -3273 5598 -3239
rect -4664 -3292 -4592 -3273
rect -3582 -3292 -3510 -3273
rect -2438 -3292 -2366 -3273
rect -1294 -3292 -1222 -3273
rect -150 -3292 -78 -3273
rect 994 -3292 1066 -3273
rect 2138 -3292 2210 -3273
rect 3282 -3292 3354 -3273
rect 4426 -3292 4498 -3273
rect 5526 -3292 5598 -3273
<< metal1 >>
rect -4602 827 5516 834
rect -4602 793 -4589 827
rect -4221 793 -4017 827
rect -3649 793 -3445 827
rect -3077 793 -2873 827
rect -2505 793 -2301 827
rect -1933 793 -1729 827
rect -1361 793 -1157 827
rect -789 793 -585 827
rect -217 793 -13 827
rect 355 793 559 827
rect 927 793 1131 827
rect 1499 793 1703 827
rect 2071 793 2275 827
rect 2643 793 2847 827
rect 3215 793 3419 827
rect 3787 793 3991 827
rect 4359 793 4563 827
rect 4931 793 5135 827
rect 5503 793 5516 827
rect -4602 786 5516 793
rect -4702 755 -4654 756
rect -4702 743 -4611 755
rect -4702 -33 -4651 743
rect -4617 -33 -4611 743
rect -4702 -45 -4611 -33
rect -4702 -263 -4654 -45
rect -4210 -46 -4200 756
rect -4038 -46 -4028 756
rect -3638 -46 -3628 756
rect -3466 -46 -3456 756
rect -3066 -46 -3056 756
rect -2894 -46 -2884 756
rect -2494 -46 -2484 756
rect -2322 -46 -2312 756
rect -1922 -46 -1912 756
rect -1750 -46 -1740 756
rect -1350 -46 -1340 756
rect -1178 -46 -1168 756
rect -778 -46 -768 756
rect -606 -46 -596 756
rect -206 -46 -196 756
rect -34 -46 -24 756
rect 366 743 548 786
rect 366 -33 383 743
rect 417 -33 497 743
rect 531 -33 548 743
rect 366 -76 548 -33
rect 938 -46 948 756
rect 1110 -46 1120 756
rect 1510 -46 1520 756
rect 1682 -46 1692 756
rect 2082 -46 2092 756
rect 2254 -46 2264 756
rect 2654 -46 2664 756
rect 2826 -46 2836 756
rect 3226 -46 3236 756
rect 3398 -46 3408 756
rect 3798 -46 3808 756
rect 3970 -46 3980 756
rect 4370 -46 4380 756
rect 4542 -46 4552 756
rect 4942 -46 4952 756
rect 5114 -46 5124 756
rect 5570 755 5618 756
rect 5525 743 5618 755
rect 5525 -33 5531 743
rect 5565 -33 5618 743
rect 5525 -45 5618 -33
rect -4602 -83 5516 -76
rect -4602 -117 -4589 -83
rect -4221 -117 -4017 -83
rect -3649 -117 -3445 -83
rect -3077 -117 -2873 -83
rect -2505 -117 -2301 -83
rect -1933 -117 -1729 -83
rect -1361 -117 -1157 -83
rect -789 -117 -585 -83
rect -217 -117 -13 -83
rect 355 -117 559 -83
rect 927 -117 1131 -83
rect 1499 -117 1703 -83
rect 2071 -117 2275 -83
rect 2643 -117 2847 -83
rect 3215 -117 3419 -83
rect 3787 -117 3991 -83
rect 4359 -117 4563 -83
rect 4931 -117 5135 -83
rect 5503 -117 5516 -83
rect -4602 -191 5516 -117
rect -4602 -225 -4589 -191
rect -4221 -225 -4017 -191
rect -3649 -225 -3445 -191
rect -3077 -225 -2873 -191
rect -2505 -225 -2301 -191
rect -1933 -225 -1729 -191
rect -1361 -225 -1157 -191
rect -789 -225 -585 -191
rect -217 -225 -13 -191
rect 355 -225 559 -191
rect 927 -225 1131 -191
rect 1499 -225 1703 -191
rect 2071 -225 2275 -191
rect 2643 -225 2847 -191
rect 3215 -225 3419 -191
rect 3787 -225 3991 -191
rect 4359 -225 4563 -191
rect 4931 -225 5135 -191
rect 5503 -225 5516 -191
rect -4602 -232 5516 -225
rect -4702 -275 -4611 -263
rect -4702 -1051 -4651 -275
rect -4617 -1051 -4611 -275
rect -4702 -1063 -4611 -1051
rect -4702 -1281 -4654 -1063
rect -4210 -1064 -4200 -262
rect -4038 -1064 -4028 -262
rect -3638 -1064 -3628 -262
rect -3466 -1064 -3456 -262
rect -3066 -1064 -3056 -262
rect -2894 -1064 -2884 -262
rect -2494 -1064 -2484 -262
rect -2322 -1064 -2312 -262
rect -1922 -1064 -1912 -262
rect -1750 -1064 -1740 -262
rect -1350 -1064 -1340 -262
rect -1178 -1064 -1168 -262
rect -778 -1064 -768 -262
rect -606 -1064 -596 -262
rect -206 -1064 -196 -262
rect -34 -1064 -24 -262
rect 366 -275 548 -232
rect 366 -1051 383 -275
rect 417 -1051 497 -275
rect 531 -1051 548 -275
rect 366 -1094 548 -1051
rect 938 -1064 948 -262
rect 1110 -1064 1120 -262
rect 1510 -1064 1520 -262
rect 1682 -1064 1692 -262
rect 2082 -1064 2092 -262
rect 2254 -1064 2264 -262
rect 2654 -1064 2664 -262
rect 2826 -1064 2836 -262
rect 3226 -1064 3236 -262
rect 3398 -1064 3408 -262
rect 3798 -1064 3808 -262
rect 3970 -1064 3980 -262
rect 4370 -1064 4380 -262
rect 4542 -1064 4552 -262
rect 4942 -1064 4952 -262
rect 5114 -1064 5124 -262
rect 5570 -263 5618 -45
rect 5525 -275 5618 -263
rect 5525 -1051 5531 -275
rect 5565 -1051 5618 -275
rect 5525 -1063 5618 -1051
rect -4602 -1101 5516 -1094
rect -4602 -1135 -4589 -1101
rect -4221 -1135 -4017 -1101
rect -3649 -1135 -3445 -1101
rect -3077 -1135 -2873 -1101
rect -2505 -1135 -2301 -1101
rect -1933 -1135 -1729 -1101
rect -1361 -1135 -1157 -1101
rect -789 -1135 -585 -1101
rect -217 -1135 -13 -1101
rect 355 -1135 559 -1101
rect 927 -1135 1131 -1101
rect 1499 -1135 1703 -1101
rect 2071 -1135 2275 -1101
rect 2643 -1135 2847 -1101
rect 3215 -1135 3419 -1101
rect 3787 -1135 3991 -1101
rect 4359 -1135 4563 -1101
rect 4931 -1135 5135 -1101
rect 5503 -1135 5516 -1101
rect -4602 -1209 5516 -1135
rect -4602 -1243 -4589 -1209
rect -4221 -1243 -4017 -1209
rect -3649 -1243 -3445 -1209
rect -3077 -1243 -2873 -1209
rect -2505 -1243 -2301 -1209
rect -1933 -1243 -1729 -1209
rect -1361 -1243 -1157 -1209
rect -789 -1243 -585 -1209
rect -217 -1243 -13 -1209
rect 355 -1243 559 -1209
rect 927 -1243 1131 -1209
rect 1499 -1243 1703 -1209
rect 2071 -1243 2275 -1209
rect 2643 -1243 2847 -1209
rect 3215 -1243 3419 -1209
rect 3787 -1243 3991 -1209
rect 4359 -1243 4563 -1209
rect 4931 -1243 5135 -1209
rect 5503 -1243 5516 -1209
rect -4602 -1250 5516 -1243
rect -4702 -1293 -4611 -1281
rect -4702 -2069 -4651 -1293
rect -4617 -2069 -4611 -1293
rect -4702 -2081 -4611 -2069
rect -4702 -2299 -4654 -2081
rect -4210 -2082 -4200 -1280
rect -4038 -2082 -4028 -1280
rect -3638 -2082 -3628 -1280
rect -3466 -2082 -3456 -1280
rect -3066 -2082 -3056 -1280
rect -2894 -2082 -2884 -1280
rect -2494 -2082 -2484 -1280
rect -2322 -2082 -2312 -1280
rect -1922 -2082 -1912 -1280
rect -1750 -2082 -1740 -1280
rect -1350 -2082 -1340 -1280
rect -1178 -2082 -1168 -1280
rect -778 -2082 -768 -1280
rect -606 -2082 -596 -1280
rect -206 -2082 -196 -1280
rect -34 -2082 -24 -1280
rect 366 -1293 548 -1250
rect 366 -2069 383 -1293
rect 417 -2069 497 -1293
rect 531 -2069 548 -1293
rect 366 -2112 548 -2069
rect 938 -2082 948 -1280
rect 1110 -2082 1120 -1280
rect 1510 -2082 1520 -1280
rect 1682 -2082 1692 -1280
rect 2082 -2082 2092 -1280
rect 2254 -2082 2264 -1280
rect 2654 -2082 2664 -1280
rect 2826 -2082 2836 -1280
rect 3226 -2082 3236 -1280
rect 3398 -2082 3408 -1280
rect 3798 -2082 3808 -1280
rect 3970 -2082 3980 -1280
rect 4370 -2082 4380 -1280
rect 4542 -2082 4552 -1280
rect 4942 -2082 4952 -1280
rect 5114 -2082 5124 -1280
rect 5570 -1281 5618 -1063
rect 5525 -1293 5618 -1281
rect 5525 -2069 5531 -1293
rect 5565 -2069 5618 -1293
rect 5525 -2081 5618 -2069
rect -4602 -2119 5516 -2112
rect -4602 -2153 -4589 -2119
rect -4221 -2153 -4017 -2119
rect -3649 -2153 -3445 -2119
rect -3077 -2153 -2873 -2119
rect -2505 -2153 -2301 -2119
rect -1933 -2153 -1729 -2119
rect -1361 -2153 -1157 -2119
rect -789 -2153 -585 -2119
rect -217 -2153 -13 -2119
rect 355 -2153 559 -2119
rect 927 -2153 1131 -2119
rect 1499 -2153 1703 -2119
rect 2071 -2153 2275 -2119
rect 2643 -2153 2847 -2119
rect 3215 -2153 3419 -2119
rect 3787 -2153 3991 -2119
rect 4359 -2153 4563 -2119
rect 4931 -2153 5135 -2119
rect 5503 -2153 5516 -2119
rect -4602 -2227 5516 -2153
rect -4602 -2261 -4589 -2227
rect -4221 -2261 -4017 -2227
rect -3649 -2261 -3445 -2227
rect -3077 -2261 -2873 -2227
rect -2505 -2261 -2301 -2227
rect -1933 -2261 -1729 -2227
rect -1361 -2261 -1157 -2227
rect -789 -2261 -585 -2227
rect -217 -2261 -13 -2227
rect 355 -2261 559 -2227
rect 927 -2261 1131 -2227
rect 1499 -2261 1703 -2227
rect 2071 -2261 2275 -2227
rect 2643 -2261 2847 -2227
rect 3215 -2261 3419 -2227
rect 3787 -2261 3991 -2227
rect 4359 -2261 4563 -2227
rect 4931 -2261 5135 -2227
rect 5503 -2261 5516 -2227
rect -4602 -2268 5516 -2261
rect -4702 -2311 -4611 -2299
rect -4702 -3087 -4651 -2311
rect -4617 -3087 -4611 -2311
rect -4702 -3099 -4611 -3087
rect -4702 -3206 -4654 -3099
rect -4210 -3100 -4200 -2298
rect -4038 -3100 -4028 -2298
rect -3638 -3100 -3628 -2298
rect -3466 -3100 -3456 -2298
rect -3066 -3100 -3056 -2298
rect -2894 -3100 -2884 -2298
rect -2494 -3100 -2484 -2298
rect -2322 -3100 -2312 -2298
rect -1922 -3100 -1912 -2298
rect -1750 -3100 -1740 -2298
rect -1350 -3100 -1340 -2298
rect -1178 -3100 -1168 -2298
rect -778 -3100 -768 -2298
rect -606 -3100 -596 -2298
rect -206 -3100 -196 -2298
rect -34 -3100 -24 -2298
rect 366 -2311 548 -2268
rect 366 -3087 383 -2311
rect 417 -3087 497 -2311
rect 531 -3087 548 -2311
rect 366 -3130 548 -3087
rect 938 -3100 948 -2298
rect 1110 -3100 1120 -2298
rect 1510 -3100 1520 -2298
rect 1682 -3100 1692 -2298
rect 2082 -3100 2092 -2298
rect 2254 -3100 2264 -2298
rect 2654 -3100 2664 -2298
rect 2826 -3100 2836 -2298
rect 3226 -3100 3236 -2298
rect 3398 -3100 3408 -2298
rect 3798 -3100 3808 -2298
rect 3970 -3100 3980 -2298
rect 4370 -3100 4380 -2298
rect 4542 -3100 4552 -2298
rect 4942 -3100 4952 -2298
rect 5114 -3100 5124 -2298
rect 5570 -2299 5618 -2081
rect 5525 -2311 5618 -2299
rect 5525 -3087 5531 -2311
rect 5565 -3087 5618 -2311
rect 5525 -3099 5618 -3087
rect -4602 -3137 5516 -3130
rect -4602 -3171 -4589 -3137
rect -4221 -3171 -4017 -3137
rect -3649 -3171 -3445 -3137
rect -3077 -3171 -2873 -3137
rect -2505 -3171 -2301 -3137
rect -1933 -3171 -1729 -3137
rect -1361 -3171 -1157 -3137
rect -789 -3171 -585 -3137
rect -217 -3171 -13 -3137
rect 355 -3171 559 -3137
rect 927 -3171 1131 -3137
rect 1499 -3171 1703 -3137
rect 2071 -3171 2275 -3137
rect 2643 -3171 2847 -3137
rect 3215 -3171 3419 -3137
rect 3787 -3171 3991 -3137
rect 4359 -3171 4563 -3137
rect 4931 -3171 5135 -3137
rect 5503 -3171 5516 -3137
rect -4602 -3178 5516 -3171
rect -4702 -3218 -4586 -3206
rect -4702 -3292 -4664 -3218
rect -4592 -3292 -4586 -3218
rect -4702 -3304 -4586 -3292
rect -3588 -3218 -3504 -3206
rect -3588 -3292 -3582 -3218
rect -3510 -3292 -3504 -3218
rect -4702 -3476 -4654 -3304
rect -4738 -3688 -4728 -3476
rect -4506 -3688 -4496 -3476
rect -3588 -3482 -3504 -3292
rect -2444 -3218 -2360 -3206
rect -2444 -3292 -2438 -3218
rect -2366 -3292 -2360 -3218
rect -2444 -3482 -2360 -3292
rect -1300 -3218 -1216 -3206
rect -1300 -3292 -1294 -3218
rect -1222 -3292 -1216 -3218
rect -1300 -3482 -1216 -3292
rect -156 -3218 -72 -3206
rect -156 -3292 -150 -3218
rect -78 -3292 -72 -3218
rect -156 -3482 -72 -3292
rect -3668 -3694 -3658 -3482
rect -3436 -3694 -3426 -3482
rect -2524 -3694 -2514 -3482
rect -2292 -3694 -2282 -3482
rect -1380 -3694 -1370 -3482
rect -1148 -3694 -1138 -3482
rect -236 -3694 -226 -3482
rect -4 -3694 6 -3482
rect 366 -4684 548 -3178
rect 5570 -3206 5618 -3099
rect 988 -3218 1072 -3206
rect 988 -3292 994 -3218
rect 1066 -3292 1072 -3218
rect 988 -3482 1072 -3292
rect 2132 -3218 2216 -3206
rect 2132 -3292 2138 -3218
rect 2210 -3292 2216 -3218
rect 2132 -3482 2216 -3292
rect 3276 -3218 3360 -3206
rect 3276 -3292 3282 -3218
rect 3354 -3292 3360 -3218
rect 3276 -3482 3360 -3292
rect 4420 -3218 4504 -3206
rect 4420 -3292 4426 -3218
rect 4498 -3292 4504 -3218
rect 4420 -3482 4504 -3292
rect 5520 -3218 5618 -3206
rect 5520 -3292 5526 -3218
rect 5598 -3292 5618 -3218
rect 5520 -3304 5618 -3292
rect 908 -3694 918 -3482
rect 1140 -3694 1150 -3482
rect 2052 -3694 2062 -3482
rect 2284 -3694 2294 -3482
rect 3196 -3694 3206 -3482
rect 3428 -3694 3438 -3482
rect 4340 -3694 4350 -3482
rect 4572 -3694 4582 -3482
rect 5570 -3596 5618 -3304
<< via1 >>
rect -4200 743 -4038 756
rect -4200 -33 -4193 743
rect -4193 -33 -4159 743
rect -4159 -33 -4079 743
rect -4079 -33 -4045 743
rect -4045 -33 -4038 743
rect -4200 -46 -4038 -33
rect -3628 743 -3466 756
rect -3628 -33 -3621 743
rect -3621 -33 -3587 743
rect -3587 -33 -3507 743
rect -3507 -33 -3473 743
rect -3473 -33 -3466 743
rect -3628 -46 -3466 -33
rect -3056 743 -2894 756
rect -3056 -33 -3049 743
rect -3049 -33 -3015 743
rect -3015 -33 -2935 743
rect -2935 -33 -2901 743
rect -2901 -33 -2894 743
rect -3056 -46 -2894 -33
rect -2484 743 -2322 756
rect -2484 -33 -2477 743
rect -2477 -33 -2443 743
rect -2443 -33 -2363 743
rect -2363 -33 -2329 743
rect -2329 -33 -2322 743
rect -2484 -46 -2322 -33
rect -1912 743 -1750 756
rect -1912 -33 -1905 743
rect -1905 -33 -1871 743
rect -1871 -33 -1791 743
rect -1791 -33 -1757 743
rect -1757 -33 -1750 743
rect -1912 -46 -1750 -33
rect -1340 743 -1178 756
rect -1340 -33 -1333 743
rect -1333 -33 -1299 743
rect -1299 -33 -1219 743
rect -1219 -33 -1185 743
rect -1185 -33 -1178 743
rect -1340 -46 -1178 -33
rect -768 743 -606 756
rect -768 -33 -761 743
rect -761 -33 -727 743
rect -727 -33 -647 743
rect -647 -33 -613 743
rect -613 -33 -606 743
rect -768 -46 -606 -33
rect -196 743 -34 756
rect -196 -33 -189 743
rect -189 -33 -155 743
rect -155 -33 -75 743
rect -75 -33 -41 743
rect -41 -33 -34 743
rect -196 -46 -34 -33
rect 948 743 1110 756
rect 948 -33 955 743
rect 955 -33 989 743
rect 989 -33 1069 743
rect 1069 -33 1103 743
rect 1103 -33 1110 743
rect 948 -46 1110 -33
rect 1520 743 1682 756
rect 1520 -33 1527 743
rect 1527 -33 1561 743
rect 1561 -33 1641 743
rect 1641 -33 1675 743
rect 1675 -33 1682 743
rect 1520 -46 1682 -33
rect 2092 743 2254 756
rect 2092 -33 2099 743
rect 2099 -33 2133 743
rect 2133 -33 2213 743
rect 2213 -33 2247 743
rect 2247 -33 2254 743
rect 2092 -46 2254 -33
rect 2664 743 2826 756
rect 2664 -33 2671 743
rect 2671 -33 2705 743
rect 2705 -33 2785 743
rect 2785 -33 2819 743
rect 2819 -33 2826 743
rect 2664 -46 2826 -33
rect 3236 743 3398 756
rect 3236 -33 3243 743
rect 3243 -33 3277 743
rect 3277 -33 3357 743
rect 3357 -33 3391 743
rect 3391 -33 3398 743
rect 3236 -46 3398 -33
rect 3808 743 3970 756
rect 3808 -33 3815 743
rect 3815 -33 3849 743
rect 3849 -33 3929 743
rect 3929 -33 3963 743
rect 3963 -33 3970 743
rect 3808 -46 3970 -33
rect 4380 743 4542 756
rect 4380 -33 4387 743
rect 4387 -33 4421 743
rect 4421 -33 4501 743
rect 4501 -33 4535 743
rect 4535 -33 4542 743
rect 4380 -46 4542 -33
rect 4952 743 5114 756
rect 4952 -33 4959 743
rect 4959 -33 4993 743
rect 4993 -33 5073 743
rect 5073 -33 5107 743
rect 5107 -33 5114 743
rect 4952 -46 5114 -33
rect -4200 -275 -4038 -262
rect -4200 -1051 -4193 -275
rect -4193 -1051 -4159 -275
rect -4159 -1051 -4079 -275
rect -4079 -1051 -4045 -275
rect -4045 -1051 -4038 -275
rect -4200 -1064 -4038 -1051
rect -3628 -275 -3466 -262
rect -3628 -1051 -3621 -275
rect -3621 -1051 -3587 -275
rect -3587 -1051 -3507 -275
rect -3507 -1051 -3473 -275
rect -3473 -1051 -3466 -275
rect -3628 -1064 -3466 -1051
rect -3056 -275 -2894 -262
rect -3056 -1051 -3049 -275
rect -3049 -1051 -3015 -275
rect -3015 -1051 -2935 -275
rect -2935 -1051 -2901 -275
rect -2901 -1051 -2894 -275
rect -3056 -1064 -2894 -1051
rect -2484 -275 -2322 -262
rect -2484 -1051 -2477 -275
rect -2477 -1051 -2443 -275
rect -2443 -1051 -2363 -275
rect -2363 -1051 -2329 -275
rect -2329 -1051 -2322 -275
rect -2484 -1064 -2322 -1051
rect -1912 -275 -1750 -262
rect -1912 -1051 -1905 -275
rect -1905 -1051 -1871 -275
rect -1871 -1051 -1791 -275
rect -1791 -1051 -1757 -275
rect -1757 -1051 -1750 -275
rect -1912 -1064 -1750 -1051
rect -1340 -275 -1178 -262
rect -1340 -1051 -1333 -275
rect -1333 -1051 -1299 -275
rect -1299 -1051 -1219 -275
rect -1219 -1051 -1185 -275
rect -1185 -1051 -1178 -275
rect -1340 -1064 -1178 -1051
rect -768 -275 -606 -262
rect -768 -1051 -761 -275
rect -761 -1051 -727 -275
rect -727 -1051 -647 -275
rect -647 -1051 -613 -275
rect -613 -1051 -606 -275
rect -768 -1064 -606 -1051
rect -196 -275 -34 -262
rect -196 -1051 -189 -275
rect -189 -1051 -155 -275
rect -155 -1051 -75 -275
rect -75 -1051 -41 -275
rect -41 -1051 -34 -275
rect -196 -1064 -34 -1051
rect 948 -275 1110 -262
rect 948 -1051 955 -275
rect 955 -1051 989 -275
rect 989 -1051 1069 -275
rect 1069 -1051 1103 -275
rect 1103 -1051 1110 -275
rect 948 -1064 1110 -1051
rect 1520 -275 1682 -262
rect 1520 -1051 1527 -275
rect 1527 -1051 1561 -275
rect 1561 -1051 1641 -275
rect 1641 -1051 1675 -275
rect 1675 -1051 1682 -275
rect 1520 -1064 1682 -1051
rect 2092 -275 2254 -262
rect 2092 -1051 2099 -275
rect 2099 -1051 2133 -275
rect 2133 -1051 2213 -275
rect 2213 -1051 2247 -275
rect 2247 -1051 2254 -275
rect 2092 -1064 2254 -1051
rect 2664 -275 2826 -262
rect 2664 -1051 2671 -275
rect 2671 -1051 2705 -275
rect 2705 -1051 2785 -275
rect 2785 -1051 2819 -275
rect 2819 -1051 2826 -275
rect 2664 -1064 2826 -1051
rect 3236 -275 3398 -262
rect 3236 -1051 3243 -275
rect 3243 -1051 3277 -275
rect 3277 -1051 3357 -275
rect 3357 -1051 3391 -275
rect 3391 -1051 3398 -275
rect 3236 -1064 3398 -1051
rect 3808 -275 3970 -262
rect 3808 -1051 3815 -275
rect 3815 -1051 3849 -275
rect 3849 -1051 3929 -275
rect 3929 -1051 3963 -275
rect 3963 -1051 3970 -275
rect 3808 -1064 3970 -1051
rect 4380 -275 4542 -262
rect 4380 -1051 4387 -275
rect 4387 -1051 4421 -275
rect 4421 -1051 4501 -275
rect 4501 -1051 4535 -275
rect 4535 -1051 4542 -275
rect 4380 -1064 4542 -1051
rect 4952 -275 5114 -262
rect 4952 -1051 4959 -275
rect 4959 -1051 4993 -275
rect 4993 -1051 5073 -275
rect 5073 -1051 5107 -275
rect 5107 -1051 5114 -275
rect 4952 -1064 5114 -1051
rect -4200 -1293 -4038 -1280
rect -4200 -2069 -4193 -1293
rect -4193 -2069 -4159 -1293
rect -4159 -2069 -4079 -1293
rect -4079 -2069 -4045 -1293
rect -4045 -2069 -4038 -1293
rect -4200 -2082 -4038 -2069
rect -3628 -1293 -3466 -1280
rect -3628 -2069 -3621 -1293
rect -3621 -2069 -3587 -1293
rect -3587 -2069 -3507 -1293
rect -3507 -2069 -3473 -1293
rect -3473 -2069 -3466 -1293
rect -3628 -2082 -3466 -2069
rect -3056 -1293 -2894 -1280
rect -3056 -2069 -3049 -1293
rect -3049 -2069 -3015 -1293
rect -3015 -2069 -2935 -1293
rect -2935 -2069 -2901 -1293
rect -2901 -2069 -2894 -1293
rect -3056 -2082 -2894 -2069
rect -2484 -1293 -2322 -1280
rect -2484 -2069 -2477 -1293
rect -2477 -2069 -2443 -1293
rect -2443 -2069 -2363 -1293
rect -2363 -2069 -2329 -1293
rect -2329 -2069 -2322 -1293
rect -2484 -2082 -2322 -2069
rect -1912 -1293 -1750 -1280
rect -1912 -2069 -1905 -1293
rect -1905 -2069 -1871 -1293
rect -1871 -2069 -1791 -1293
rect -1791 -2069 -1757 -1293
rect -1757 -2069 -1750 -1293
rect -1912 -2082 -1750 -2069
rect -1340 -1293 -1178 -1280
rect -1340 -2069 -1333 -1293
rect -1333 -2069 -1299 -1293
rect -1299 -2069 -1219 -1293
rect -1219 -2069 -1185 -1293
rect -1185 -2069 -1178 -1293
rect -1340 -2082 -1178 -2069
rect -768 -1293 -606 -1280
rect -768 -2069 -761 -1293
rect -761 -2069 -727 -1293
rect -727 -2069 -647 -1293
rect -647 -2069 -613 -1293
rect -613 -2069 -606 -1293
rect -768 -2082 -606 -2069
rect -196 -1293 -34 -1280
rect -196 -2069 -189 -1293
rect -189 -2069 -155 -1293
rect -155 -2069 -75 -1293
rect -75 -2069 -41 -1293
rect -41 -2069 -34 -1293
rect -196 -2082 -34 -2069
rect 948 -1293 1110 -1280
rect 948 -2069 955 -1293
rect 955 -2069 989 -1293
rect 989 -2069 1069 -1293
rect 1069 -2069 1103 -1293
rect 1103 -2069 1110 -1293
rect 948 -2082 1110 -2069
rect 1520 -1293 1682 -1280
rect 1520 -2069 1527 -1293
rect 1527 -2069 1561 -1293
rect 1561 -2069 1641 -1293
rect 1641 -2069 1675 -1293
rect 1675 -2069 1682 -1293
rect 1520 -2082 1682 -2069
rect 2092 -1293 2254 -1280
rect 2092 -2069 2099 -1293
rect 2099 -2069 2133 -1293
rect 2133 -2069 2213 -1293
rect 2213 -2069 2247 -1293
rect 2247 -2069 2254 -1293
rect 2092 -2082 2254 -2069
rect 2664 -1293 2826 -1280
rect 2664 -2069 2671 -1293
rect 2671 -2069 2705 -1293
rect 2705 -2069 2785 -1293
rect 2785 -2069 2819 -1293
rect 2819 -2069 2826 -1293
rect 2664 -2082 2826 -2069
rect 3236 -1293 3398 -1280
rect 3236 -2069 3243 -1293
rect 3243 -2069 3277 -1293
rect 3277 -2069 3357 -1293
rect 3357 -2069 3391 -1293
rect 3391 -2069 3398 -1293
rect 3236 -2082 3398 -2069
rect 3808 -1293 3970 -1280
rect 3808 -2069 3815 -1293
rect 3815 -2069 3849 -1293
rect 3849 -2069 3929 -1293
rect 3929 -2069 3963 -1293
rect 3963 -2069 3970 -1293
rect 3808 -2082 3970 -2069
rect 4380 -1293 4542 -1280
rect 4380 -2069 4387 -1293
rect 4387 -2069 4421 -1293
rect 4421 -2069 4501 -1293
rect 4501 -2069 4535 -1293
rect 4535 -2069 4542 -1293
rect 4380 -2082 4542 -2069
rect 4952 -1293 5114 -1280
rect 4952 -2069 4959 -1293
rect 4959 -2069 4993 -1293
rect 4993 -2069 5073 -1293
rect 5073 -2069 5107 -1293
rect 5107 -2069 5114 -1293
rect 4952 -2082 5114 -2069
rect -4200 -2311 -4038 -2298
rect -4200 -3087 -4193 -2311
rect -4193 -3087 -4159 -2311
rect -4159 -3087 -4079 -2311
rect -4079 -3087 -4045 -2311
rect -4045 -3087 -4038 -2311
rect -4200 -3100 -4038 -3087
rect -3628 -2311 -3466 -2298
rect -3628 -3087 -3621 -2311
rect -3621 -3087 -3587 -2311
rect -3587 -3087 -3507 -2311
rect -3507 -3087 -3473 -2311
rect -3473 -3087 -3466 -2311
rect -3628 -3100 -3466 -3087
rect -3056 -2311 -2894 -2298
rect -3056 -3087 -3049 -2311
rect -3049 -3087 -3015 -2311
rect -3015 -3087 -2935 -2311
rect -2935 -3087 -2901 -2311
rect -2901 -3087 -2894 -2311
rect -3056 -3100 -2894 -3087
rect -2484 -2311 -2322 -2298
rect -2484 -3087 -2477 -2311
rect -2477 -3087 -2443 -2311
rect -2443 -3087 -2363 -2311
rect -2363 -3087 -2329 -2311
rect -2329 -3087 -2322 -2311
rect -2484 -3100 -2322 -3087
rect -1912 -2311 -1750 -2298
rect -1912 -3087 -1905 -2311
rect -1905 -3087 -1871 -2311
rect -1871 -3087 -1791 -2311
rect -1791 -3087 -1757 -2311
rect -1757 -3087 -1750 -2311
rect -1912 -3100 -1750 -3087
rect -1340 -2311 -1178 -2298
rect -1340 -3087 -1333 -2311
rect -1333 -3087 -1299 -2311
rect -1299 -3087 -1219 -2311
rect -1219 -3087 -1185 -2311
rect -1185 -3087 -1178 -2311
rect -1340 -3100 -1178 -3087
rect -768 -2311 -606 -2298
rect -768 -3087 -761 -2311
rect -761 -3087 -727 -2311
rect -727 -3087 -647 -2311
rect -647 -3087 -613 -2311
rect -613 -3087 -606 -2311
rect -768 -3100 -606 -3087
rect -196 -2311 -34 -2298
rect -196 -3087 -189 -2311
rect -189 -3087 -155 -2311
rect -155 -3087 -75 -2311
rect -75 -3087 -41 -2311
rect -41 -3087 -34 -2311
rect -196 -3100 -34 -3087
rect 948 -2311 1110 -2298
rect 948 -3087 955 -2311
rect 955 -3087 989 -2311
rect 989 -3087 1069 -2311
rect 1069 -3087 1103 -2311
rect 1103 -3087 1110 -2311
rect 948 -3100 1110 -3087
rect 1520 -2311 1682 -2298
rect 1520 -3087 1527 -2311
rect 1527 -3087 1561 -2311
rect 1561 -3087 1641 -2311
rect 1641 -3087 1675 -2311
rect 1675 -3087 1682 -2311
rect 1520 -3100 1682 -3087
rect 2092 -2311 2254 -2298
rect 2092 -3087 2099 -2311
rect 2099 -3087 2133 -2311
rect 2133 -3087 2213 -2311
rect 2213 -3087 2247 -2311
rect 2247 -3087 2254 -2311
rect 2092 -3100 2254 -3087
rect 2664 -2311 2826 -2298
rect 2664 -3087 2671 -2311
rect 2671 -3087 2705 -2311
rect 2705 -3087 2785 -2311
rect 2785 -3087 2819 -2311
rect 2819 -3087 2826 -2311
rect 2664 -3100 2826 -3087
rect 3236 -2311 3398 -2298
rect 3236 -3087 3243 -2311
rect 3243 -3087 3277 -2311
rect 3277 -3087 3357 -2311
rect 3357 -3087 3391 -2311
rect 3391 -3087 3398 -2311
rect 3236 -3100 3398 -3087
rect 3808 -2311 3970 -2298
rect 3808 -3087 3815 -2311
rect 3815 -3087 3849 -2311
rect 3849 -3087 3929 -2311
rect 3929 -3087 3963 -2311
rect 3963 -3087 3970 -2311
rect 3808 -3100 3970 -3087
rect 4380 -2311 4542 -2298
rect 4380 -3087 4387 -2311
rect 4387 -3087 4421 -2311
rect 4421 -3087 4501 -2311
rect 4501 -3087 4535 -2311
rect 4535 -3087 4542 -2311
rect 4380 -3100 4542 -3087
rect 4952 -2311 5114 -2298
rect 4952 -3087 4959 -2311
rect 4959 -3087 4993 -2311
rect 4993 -3087 5073 -2311
rect 5073 -3087 5107 -2311
rect 5107 -3087 5114 -2311
rect 4952 -3100 5114 -3087
rect -4728 -3688 -4506 -3476
rect -3658 -3694 -3436 -3482
rect -2514 -3694 -2292 -3482
rect -1370 -3694 -1148 -3482
rect -226 -3694 -4 -3482
rect 918 -3694 1140 -3482
rect 2062 -3694 2284 -3482
rect 3206 -3694 3428 -3482
rect 4350 -3694 4572 -3482
<< metal2 >>
rect -4210 756 -4028 1016
rect -4210 -46 -4200 756
rect -4038 -46 -4028 756
rect -4210 -262 -4028 -46
rect -4210 -1064 -4200 -262
rect -4038 -1064 -4028 -262
rect -4210 -1280 -4028 -1064
rect -4210 -2082 -4200 -1280
rect -4038 -2082 -4028 -1280
rect -4210 -2298 -4028 -2082
rect -4210 -3100 -4200 -2298
rect -4038 -3100 -4028 -2298
rect -4210 -3110 -4028 -3100
rect -3638 756 -3456 766
rect -3638 -46 -3628 756
rect -3466 -46 -3456 756
rect -3638 -262 -3456 -46
rect -3638 -1064 -3628 -262
rect -3466 -1064 -3456 -262
rect -3638 -1280 -3456 -1064
rect -3638 -2082 -3628 -1280
rect -3466 -2082 -3456 -1280
rect -3638 -2298 -3456 -2082
rect -3638 -3100 -3628 -2298
rect -3466 -3100 -3456 -2298
rect -4728 -3476 -4506 -3466
rect -3638 -3472 -3456 -3100
rect -3066 756 -2884 1016
rect -3066 -46 -3056 756
rect -2894 -46 -2884 756
rect -3066 -262 -2884 -46
rect -3066 -1064 -3056 -262
rect -2894 -1064 -2884 -262
rect -3066 -1280 -2884 -1064
rect -3066 -2082 -3056 -1280
rect -2894 -2082 -2884 -1280
rect -3066 -2298 -2884 -2082
rect -3066 -3100 -3056 -2298
rect -2894 -3100 -2884 -2298
rect -3066 -3110 -2884 -3100
rect -2494 756 -2312 766
rect -2494 -46 -2484 756
rect -2322 -46 -2312 756
rect -2494 -262 -2312 -46
rect -2494 -1064 -2484 -262
rect -2322 -1064 -2312 -262
rect -2494 -1280 -2312 -1064
rect -2494 -2082 -2484 -1280
rect -2322 -2082 -2312 -1280
rect -2494 -2298 -2312 -2082
rect -2494 -3100 -2484 -2298
rect -2322 -3100 -2312 -2298
rect -2494 -3472 -2312 -3100
rect -1922 756 -1740 1016
rect -1922 -46 -1912 756
rect -1750 -46 -1740 756
rect -1922 -262 -1740 -46
rect -1922 -1064 -1912 -262
rect -1750 -1064 -1740 -262
rect -1922 -1280 -1740 -1064
rect -1922 -2082 -1912 -1280
rect -1750 -2082 -1740 -1280
rect -1922 -2298 -1740 -2082
rect -1922 -3100 -1912 -2298
rect -1750 -3100 -1740 -2298
rect -1922 -3110 -1740 -3100
rect -1350 756 -1168 766
rect -1350 -46 -1340 756
rect -1178 -46 -1168 756
rect -1350 -262 -1168 -46
rect -1350 -1064 -1340 -262
rect -1178 -1064 -1168 -262
rect -1350 -1280 -1168 -1064
rect -1350 -2082 -1340 -1280
rect -1178 -2082 -1168 -1280
rect -1350 -2298 -1168 -2082
rect -1350 -3100 -1340 -2298
rect -1178 -3100 -1168 -2298
rect -1350 -3472 -1168 -3100
rect -778 756 -596 1016
rect -778 -46 -768 756
rect -606 -46 -596 756
rect -778 -262 -596 -46
rect -778 -1064 -768 -262
rect -606 -1064 -596 -262
rect -778 -1280 -596 -1064
rect -778 -2082 -768 -1280
rect -606 -2082 -596 -1280
rect -778 -2298 -596 -2082
rect -778 -3100 -768 -2298
rect -606 -3100 -596 -2298
rect -778 -3110 -596 -3100
rect -206 756 -24 766
rect -206 -46 -196 756
rect -34 -46 -24 756
rect -206 -262 -24 -46
rect -206 -1064 -196 -262
rect -34 -1064 -24 -262
rect -206 -1280 -24 -1064
rect -206 -2082 -196 -1280
rect -34 -2082 -24 -1280
rect -206 -2298 -24 -2082
rect -206 -3100 -196 -2298
rect -34 -3100 -24 -2298
rect -206 -3472 -24 -3100
rect 938 756 1120 766
rect 938 -46 948 756
rect 1110 -46 1120 756
rect 938 -262 1120 -46
rect 938 -1064 948 -262
rect 1110 -1064 1120 -262
rect 938 -1280 1120 -1064
rect 938 -2082 948 -1280
rect 1110 -2082 1120 -1280
rect 938 -2298 1120 -2082
rect 938 -3100 948 -2298
rect 1110 -3100 1120 -2298
rect 938 -3472 1120 -3100
rect 1510 756 1692 1016
rect 1510 -46 1520 756
rect 1682 -46 1692 756
rect 1510 -262 1692 -46
rect 1510 -1064 1520 -262
rect 1682 -1064 1692 -262
rect 1510 -1280 1692 -1064
rect 1510 -2082 1520 -1280
rect 1682 -2082 1692 -1280
rect 1510 -2298 1692 -2082
rect 1510 -3100 1520 -2298
rect 1682 -3100 1692 -2298
rect 1510 -3110 1692 -3100
rect 2082 756 2264 766
rect 2082 -46 2092 756
rect 2254 -46 2264 756
rect 2082 -262 2264 -46
rect 2082 -1064 2092 -262
rect 2254 -1064 2264 -262
rect 2082 -1280 2264 -1064
rect 2082 -2082 2092 -1280
rect 2254 -2082 2264 -1280
rect 2082 -2298 2264 -2082
rect 2082 -3100 2092 -2298
rect 2254 -3100 2264 -2298
rect 2082 -3472 2264 -3100
rect 2654 756 2836 1016
rect 2654 -46 2664 756
rect 2826 -46 2836 756
rect 2654 -262 2836 -46
rect 2654 -1064 2664 -262
rect 2826 -1064 2836 -262
rect 2654 -1280 2836 -1064
rect 2654 -2082 2664 -1280
rect 2826 -2082 2836 -1280
rect 2654 -2298 2836 -2082
rect 2654 -3100 2664 -2298
rect 2826 -3100 2836 -2298
rect 2654 -3110 2836 -3100
rect 3226 756 3408 766
rect 3226 -46 3236 756
rect 3398 -46 3408 756
rect 3226 -262 3408 -46
rect 3226 -1064 3236 -262
rect 3398 -1064 3408 -262
rect 3226 -1280 3408 -1064
rect 3226 -2082 3236 -1280
rect 3398 -2082 3408 -1280
rect 3226 -2298 3408 -2082
rect 3226 -3100 3236 -2298
rect 3398 -3100 3408 -2298
rect 3226 -3472 3408 -3100
rect 3798 756 3980 1016
rect 3798 -46 3808 756
rect 3970 -46 3980 756
rect 3798 -262 3980 -46
rect 3798 -1064 3808 -262
rect 3970 -1064 3980 -262
rect 3798 -1280 3980 -1064
rect 3798 -2082 3808 -1280
rect 3970 -2082 3980 -1280
rect 3798 -2298 3980 -2082
rect 3798 -3100 3808 -2298
rect 3970 -3100 3980 -2298
rect 3798 -3110 3980 -3100
rect 4370 756 4552 766
rect 4370 -46 4380 756
rect 4542 -46 4552 756
rect 4370 -262 4552 -46
rect 4370 -1064 4380 -262
rect 4542 -1064 4552 -262
rect 4370 -1280 4552 -1064
rect 4370 -2082 4380 -1280
rect 4542 -2082 4552 -1280
rect 4370 -2298 4552 -2082
rect 4370 -3100 4380 -2298
rect 4542 -3100 4552 -2298
rect 4370 -3472 4552 -3100
rect 4942 756 5124 1016
rect 4942 -46 4952 756
rect 5114 -46 5124 756
rect 4942 -262 5124 -46
rect 4942 -1064 4952 -262
rect 5114 -1064 5124 -262
rect 4942 -1280 5124 -1064
rect 4942 -2082 4952 -1280
rect 5114 -2082 5124 -1280
rect 4942 -2298 5124 -2082
rect 4942 -3100 4952 -2298
rect 5114 -3100 5124 -2298
rect 4942 -3110 5124 -3100
rect 5514 -3472 5696 -3466
rect -4728 -3698 -4506 -3688
rect -3658 -3482 -3436 -3472
rect -3658 -3704 -3436 -3694
rect -2514 -3482 -2292 -3472
rect -2514 -3704 -2292 -3694
rect -1370 -3482 -1148 -3472
rect -1370 -3704 -1148 -3694
rect -226 -3482 -4 -3472
rect -226 -3704 -4 -3694
rect 918 -3482 1140 -3472
rect 918 -3704 1140 -3694
rect 2062 -3482 2284 -3472
rect 2062 -3704 2284 -3694
rect 3206 -3482 3428 -3472
rect 3206 -3704 3428 -3694
rect 4350 -3482 4572 -3472
rect 4350 -3704 4572 -3694
rect 5494 -3482 5716 -3472
rect 5494 -3704 5716 -3694
<< via2 >>
rect -4728 -3688 -4506 -3476
rect -3658 -3694 -3436 -3482
rect -2514 -3694 -2292 -3482
rect -1370 -3694 -1148 -3482
rect -226 -3694 -4 -3482
rect 918 -3694 1140 -3482
rect 2062 -3694 2284 -3482
rect 3206 -3694 3428 -3482
rect 4350 -3694 4572 -3482
rect 5494 -3694 5716 -3482
<< metal3 >>
rect -4758 -3476 5802 -3406
rect -4758 -3688 -4728 -3476
rect -4506 -3482 5802 -3476
rect -4506 -3688 -3658 -3482
rect -4758 -3694 -3658 -3688
rect -3436 -3694 -2514 -3482
rect -2292 -3694 -1370 -3482
rect -1148 -3694 -226 -3482
rect -4 -3694 918 -3482
rect 1140 -3694 2062 -3482
rect 2284 -3694 3206 -3482
rect 3428 -3694 4350 -3482
rect 4572 -3694 5494 -3482
rect 5716 -3694 5802 -3482
rect -4758 -4296 5802 -3694
<< labels >>
flabel metal2 -4130 990 -4130 990 0 FreeSans 1600 0 0 0 vbias1
port 1 nsew
flabel metal2 -2968 990 -2968 990 0 FreeSans 1600 0 0 0 vbias2
port 2 nsew
flabel metal2 -1836 998 -1836 998 0 FreeSans 1600 0 0 0 vbias3
port 3 nsew
flabel metal2 -702 982 -702 982 0 FreeSans 1600 0 0 0 vbias4
port 4 nsew
flabel metal2 1608 992 1608 992 0 FreeSans 1600 0 0 0 vbias5
port 5 nsew
flabel metal2 2760 986 2760 986 0 FreeSans 1600 0 0 0 vbias6
port 6 nsew
flabel metal2 3884 992 3884 992 0 FreeSans 1600 0 0 0 vbias7
port 7 nsew
flabel metal2 5042 1000 5042 1000 0 FreeSans 1600 0 0 0 vbias8
port 8 nsew
flabel metal1 462 -4564 462 -4564 0 FreeSans 1600 0 0 0 iin
port 0 nsew
flabel metal3 -1680 -3950 -1680 -3950 0 FreeSans 1600 0 0 0 vss
port 9 nsew
<< end >>
