magic
tech sky130A
magscale 1 2
timestamp 1629189639
<< isosubstrate >>
rect 54142 8686 55900 11460
<< nwell >>
rect 37859 7151 49983 9261
rect 39347 2527 42543 6873
<< pwell >>
rect 42973 3203 43375 4959
rect 39347 305 48495 2179
<< pmoslvt >>
rect 38055 8642 38255 9042
rect 38427 8642 38627 9042
rect 38799 8642 38999 9042
rect 39171 8642 39371 9042
rect 39543 8642 39743 9042
rect 39915 8642 40115 9042
rect 40287 8642 40487 9042
rect 40659 8642 40859 9042
rect 41031 8642 41231 9042
rect 41403 8642 41603 9042
rect 41775 8642 41975 9042
rect 42147 8642 42347 9042
rect 42519 8642 42719 9042
rect 42891 8642 43091 9042
rect 43263 8642 43463 9042
rect 43635 8642 43835 9042
rect 44007 8642 44207 9042
rect 44379 8642 44579 9042
rect 44751 8642 44951 9042
rect 45123 8642 45323 9042
rect 45495 8642 45695 9042
rect 45867 8642 46067 9042
rect 46239 8642 46439 9042
rect 46611 8642 46811 9042
rect 46983 8642 47183 9042
rect 47355 8642 47555 9042
rect 47727 8642 47927 9042
rect 48099 8642 48299 9042
rect 48471 8642 48671 9042
rect 48843 8642 49043 9042
rect 49215 8642 49415 9042
rect 49587 8642 49787 9042
rect 38055 8006 38255 8406
rect 38427 8006 38627 8406
rect 38799 8006 38999 8406
rect 39171 8006 39371 8406
rect 39543 8006 39743 8406
rect 39915 8006 40115 8406
rect 40287 8006 40487 8406
rect 40659 8006 40859 8406
rect 41031 8006 41231 8406
rect 41403 8006 41603 8406
rect 41775 8006 41975 8406
rect 42147 8006 42347 8406
rect 42519 8006 42719 8406
rect 42891 8006 43091 8406
rect 43263 8006 43463 8406
rect 43635 8006 43835 8406
rect 44007 8006 44207 8406
rect 44379 8006 44579 8406
rect 44751 8006 44951 8406
rect 45123 8006 45323 8406
rect 45495 8006 45695 8406
rect 45867 8006 46067 8406
rect 46239 8006 46439 8406
rect 46611 8006 46811 8406
rect 46983 8006 47183 8406
rect 47355 8006 47555 8406
rect 47727 8006 47927 8406
rect 48099 8006 48299 8406
rect 48471 8006 48671 8406
rect 48843 8006 49043 8406
rect 49215 8006 49415 8406
rect 49587 8006 49787 8406
rect 38055 7370 38255 7770
rect 38427 7370 38627 7770
rect 38799 7370 38999 7770
rect 39171 7370 39371 7770
rect 39543 7370 39743 7770
rect 39915 7370 40115 7770
rect 40287 7370 40487 7770
rect 40659 7370 40859 7770
rect 41031 7370 41231 7770
rect 41403 7370 41603 7770
rect 41775 7370 41975 7770
rect 42147 7370 42347 7770
rect 42519 7370 42719 7770
rect 42891 7370 43091 7770
rect 43263 7370 43463 7770
rect 43635 7370 43835 7770
rect 44007 7370 44207 7770
rect 44379 7370 44579 7770
rect 44751 7370 44951 7770
rect 45123 7370 45323 7770
rect 45495 7370 45695 7770
rect 45867 7370 46067 7770
rect 46239 7370 46439 7770
rect 46611 7370 46811 7770
rect 46983 7370 47183 7770
rect 47355 7370 47555 7770
rect 47727 7370 47927 7770
rect 48099 7370 48299 7770
rect 48471 7370 48671 7770
rect 48843 7370 49043 7770
rect 49215 7370 49415 7770
rect 49587 7370 49787 7770
rect 39543 5854 39743 6654
rect 39915 5854 40115 6654
rect 40287 5854 40487 6654
rect 40659 5854 40859 6654
rect 41031 5854 41231 6654
rect 41403 5854 41603 6654
rect 41775 5854 41975 6654
rect 42147 5854 42347 6654
rect 39543 4818 39743 5618
rect 39915 4818 40115 5618
rect 40287 4818 40487 5618
rect 40659 4818 40859 5618
rect 41031 4818 41231 5618
rect 41403 4818 41603 5618
rect 41775 4818 41975 5618
rect 42147 4818 42347 5618
rect 39543 3782 39743 4582
rect 39915 3782 40115 4582
rect 40287 3782 40487 4582
rect 40659 3782 40859 4582
rect 41031 3782 41231 4582
rect 41403 3782 41603 4582
rect 41775 3782 41975 4582
rect 42147 3782 42347 4582
rect 39543 2746 39743 3546
rect 39915 2746 40115 3546
rect 40287 2746 40487 3546
rect 40659 2746 40859 3546
rect 41031 2746 41231 3546
rect 41403 2746 41603 3546
rect 41775 2746 41975 3546
rect 42147 2746 42347 3546
<< nmoslvt >>
rect 39543 1769 39743 1969
rect 39915 1769 40115 1969
rect 40287 1769 40487 1969
rect 40659 1769 40859 1969
rect 41031 1769 41231 1969
rect 41403 1769 41603 1969
rect 41775 1769 41975 1969
rect 42147 1769 42347 1969
rect 42519 1769 42719 1969
rect 42891 1769 43091 1969
rect 43263 1769 43463 1969
rect 43635 1769 43835 1969
rect 44007 1769 44207 1969
rect 44379 1769 44579 1969
rect 44751 1769 44951 1969
rect 45123 1769 45323 1969
rect 45495 1769 45695 1969
rect 45867 1769 46067 1969
rect 46239 1769 46439 1969
rect 46611 1769 46811 1969
rect 46983 1769 47183 1969
rect 47355 1769 47555 1969
rect 47727 1769 47927 1969
rect 48099 1769 48299 1969
rect 39543 1351 39743 1551
rect 39915 1351 40115 1551
rect 40287 1351 40487 1551
rect 40659 1351 40859 1551
rect 41031 1351 41231 1551
rect 41403 1351 41603 1551
rect 41775 1351 41975 1551
rect 42147 1351 42347 1551
rect 42519 1351 42719 1551
rect 42891 1351 43091 1551
rect 43263 1351 43463 1551
rect 43635 1351 43835 1551
rect 44007 1351 44207 1551
rect 44379 1351 44579 1551
rect 44751 1351 44951 1551
rect 45123 1351 45323 1551
rect 45495 1351 45695 1551
rect 45867 1351 46067 1551
rect 46239 1351 46439 1551
rect 46611 1351 46811 1551
rect 46983 1351 47183 1551
rect 47355 1351 47555 1551
rect 47727 1351 47927 1551
rect 48099 1351 48299 1551
rect 39543 933 39743 1133
rect 39915 933 40115 1133
rect 40287 933 40487 1133
rect 40659 933 40859 1133
rect 41031 933 41231 1133
rect 41403 933 41603 1133
rect 41775 933 41975 1133
rect 42147 933 42347 1133
rect 42519 933 42719 1133
rect 42891 933 43091 1133
rect 43263 933 43463 1133
rect 43635 933 43835 1133
rect 44007 933 44207 1133
rect 44379 933 44579 1133
rect 44751 933 44951 1133
rect 45123 933 45323 1133
rect 45495 933 45695 1133
rect 45867 933 46067 1133
rect 46239 933 46439 1133
rect 46611 933 46811 1133
rect 46983 933 47183 1133
rect 47355 933 47555 1133
rect 47727 933 47927 1133
rect 48099 933 48299 1133
rect 39543 515 39743 715
rect 39915 515 40115 715
rect 40287 515 40487 715
rect 40659 515 40859 715
rect 41031 515 41231 715
rect 41403 515 41603 715
rect 41775 515 41975 715
rect 42147 515 42347 715
rect 42519 515 42719 715
rect 42891 515 43091 715
rect 43263 515 43463 715
rect 43635 515 43835 715
rect 44007 515 44207 715
rect 44379 515 44579 715
rect 44751 515 44951 715
rect 45123 515 45323 715
rect 45495 515 45695 715
rect 45867 515 46067 715
rect 46239 515 46439 715
rect 46611 515 46811 715
rect 46983 515 47183 715
rect 47355 515 47555 715
rect 47727 515 47927 715
rect 48099 515 48299 715
<< ndiff >>
rect 39485 1957 39543 1969
rect 39485 1781 39497 1957
rect 39531 1781 39543 1957
rect 39485 1769 39543 1781
rect 39743 1957 39801 1969
rect 39743 1781 39755 1957
rect 39789 1781 39801 1957
rect 39743 1769 39801 1781
rect 39857 1957 39915 1969
rect 39857 1781 39869 1957
rect 39903 1781 39915 1957
rect 39857 1769 39915 1781
rect 40115 1957 40173 1969
rect 40115 1781 40127 1957
rect 40161 1781 40173 1957
rect 40115 1769 40173 1781
rect 40229 1957 40287 1969
rect 40229 1781 40241 1957
rect 40275 1781 40287 1957
rect 40229 1769 40287 1781
rect 40487 1957 40545 1969
rect 40487 1781 40499 1957
rect 40533 1781 40545 1957
rect 40487 1769 40545 1781
rect 40601 1957 40659 1969
rect 40601 1781 40613 1957
rect 40647 1781 40659 1957
rect 40601 1769 40659 1781
rect 40859 1957 40917 1969
rect 40859 1781 40871 1957
rect 40905 1781 40917 1957
rect 40859 1769 40917 1781
rect 40973 1957 41031 1969
rect 40973 1781 40985 1957
rect 41019 1781 41031 1957
rect 40973 1769 41031 1781
rect 41231 1957 41289 1969
rect 41231 1781 41243 1957
rect 41277 1781 41289 1957
rect 41231 1769 41289 1781
rect 41345 1957 41403 1969
rect 41345 1781 41357 1957
rect 41391 1781 41403 1957
rect 41345 1769 41403 1781
rect 41603 1957 41661 1969
rect 41603 1781 41615 1957
rect 41649 1781 41661 1957
rect 41603 1769 41661 1781
rect 41717 1957 41775 1969
rect 41717 1781 41729 1957
rect 41763 1781 41775 1957
rect 41717 1769 41775 1781
rect 41975 1957 42033 1969
rect 41975 1781 41987 1957
rect 42021 1781 42033 1957
rect 41975 1769 42033 1781
rect 42089 1957 42147 1969
rect 42089 1781 42101 1957
rect 42135 1781 42147 1957
rect 42089 1769 42147 1781
rect 42347 1957 42405 1969
rect 42347 1781 42359 1957
rect 42393 1781 42405 1957
rect 42347 1769 42405 1781
rect 42461 1957 42519 1969
rect 42461 1781 42473 1957
rect 42507 1781 42519 1957
rect 42461 1769 42519 1781
rect 42719 1957 42777 1969
rect 42719 1781 42731 1957
rect 42765 1781 42777 1957
rect 42719 1769 42777 1781
rect 42833 1957 42891 1969
rect 42833 1781 42845 1957
rect 42879 1781 42891 1957
rect 42833 1769 42891 1781
rect 43091 1957 43149 1969
rect 43091 1781 43103 1957
rect 43137 1781 43149 1957
rect 43091 1769 43149 1781
rect 43205 1957 43263 1969
rect 43205 1781 43217 1957
rect 43251 1781 43263 1957
rect 43205 1769 43263 1781
rect 43463 1957 43521 1969
rect 43463 1781 43475 1957
rect 43509 1781 43521 1957
rect 43463 1769 43521 1781
rect 43577 1957 43635 1969
rect 43577 1781 43589 1957
rect 43623 1781 43635 1957
rect 43577 1769 43635 1781
rect 43835 1957 43893 1969
rect 43835 1781 43847 1957
rect 43881 1781 43893 1957
rect 43835 1769 43893 1781
rect 43949 1957 44007 1969
rect 43949 1781 43961 1957
rect 43995 1781 44007 1957
rect 43949 1769 44007 1781
rect 44207 1957 44265 1969
rect 44207 1781 44219 1957
rect 44253 1781 44265 1957
rect 44207 1769 44265 1781
rect 44321 1957 44379 1969
rect 44321 1781 44333 1957
rect 44367 1781 44379 1957
rect 44321 1769 44379 1781
rect 44579 1957 44637 1969
rect 44579 1781 44591 1957
rect 44625 1781 44637 1957
rect 44579 1769 44637 1781
rect 44693 1957 44751 1969
rect 44693 1781 44705 1957
rect 44739 1781 44751 1957
rect 44693 1769 44751 1781
rect 44951 1957 45009 1969
rect 44951 1781 44963 1957
rect 44997 1781 45009 1957
rect 44951 1769 45009 1781
rect 45065 1957 45123 1969
rect 45065 1781 45077 1957
rect 45111 1781 45123 1957
rect 45065 1769 45123 1781
rect 45323 1957 45381 1969
rect 45323 1781 45335 1957
rect 45369 1781 45381 1957
rect 45323 1769 45381 1781
rect 45437 1957 45495 1969
rect 45437 1781 45449 1957
rect 45483 1781 45495 1957
rect 45437 1769 45495 1781
rect 45695 1957 45753 1969
rect 45695 1781 45707 1957
rect 45741 1781 45753 1957
rect 45695 1769 45753 1781
rect 45809 1957 45867 1969
rect 45809 1781 45821 1957
rect 45855 1781 45867 1957
rect 45809 1769 45867 1781
rect 46067 1957 46125 1969
rect 46067 1781 46079 1957
rect 46113 1781 46125 1957
rect 46067 1769 46125 1781
rect 46181 1957 46239 1969
rect 46181 1781 46193 1957
rect 46227 1781 46239 1957
rect 46181 1769 46239 1781
rect 46439 1957 46497 1969
rect 46439 1781 46451 1957
rect 46485 1781 46497 1957
rect 46439 1769 46497 1781
rect 46553 1957 46611 1969
rect 46553 1781 46565 1957
rect 46599 1781 46611 1957
rect 46553 1769 46611 1781
rect 46811 1957 46869 1969
rect 46811 1781 46823 1957
rect 46857 1781 46869 1957
rect 46811 1769 46869 1781
rect 46925 1957 46983 1969
rect 46925 1781 46937 1957
rect 46971 1781 46983 1957
rect 46925 1769 46983 1781
rect 47183 1957 47241 1969
rect 47183 1781 47195 1957
rect 47229 1781 47241 1957
rect 47183 1769 47241 1781
rect 47297 1957 47355 1969
rect 47297 1781 47309 1957
rect 47343 1781 47355 1957
rect 47297 1769 47355 1781
rect 47555 1957 47613 1969
rect 47555 1781 47567 1957
rect 47601 1781 47613 1957
rect 47555 1769 47613 1781
rect 47669 1957 47727 1969
rect 47669 1781 47681 1957
rect 47715 1781 47727 1957
rect 47669 1769 47727 1781
rect 47927 1957 47985 1969
rect 47927 1781 47939 1957
rect 47973 1781 47985 1957
rect 47927 1769 47985 1781
rect 48041 1957 48099 1969
rect 48041 1781 48053 1957
rect 48087 1781 48099 1957
rect 48041 1769 48099 1781
rect 48299 1957 48357 1969
rect 48299 1781 48311 1957
rect 48345 1781 48357 1957
rect 48299 1769 48357 1781
rect 39485 1539 39543 1551
rect 39485 1363 39497 1539
rect 39531 1363 39543 1539
rect 39485 1351 39543 1363
rect 39743 1539 39801 1551
rect 39743 1363 39755 1539
rect 39789 1363 39801 1539
rect 39743 1351 39801 1363
rect 39857 1539 39915 1551
rect 39857 1363 39869 1539
rect 39903 1363 39915 1539
rect 39857 1351 39915 1363
rect 40115 1539 40173 1551
rect 40115 1363 40127 1539
rect 40161 1363 40173 1539
rect 40115 1351 40173 1363
rect 40229 1539 40287 1551
rect 40229 1363 40241 1539
rect 40275 1363 40287 1539
rect 40229 1351 40287 1363
rect 40487 1539 40545 1551
rect 40487 1363 40499 1539
rect 40533 1363 40545 1539
rect 40487 1351 40545 1363
rect 40601 1539 40659 1551
rect 40601 1363 40613 1539
rect 40647 1363 40659 1539
rect 40601 1351 40659 1363
rect 40859 1539 40917 1551
rect 40859 1363 40871 1539
rect 40905 1363 40917 1539
rect 40859 1351 40917 1363
rect 40973 1539 41031 1551
rect 40973 1363 40985 1539
rect 41019 1363 41031 1539
rect 40973 1351 41031 1363
rect 41231 1539 41289 1551
rect 41231 1363 41243 1539
rect 41277 1363 41289 1539
rect 41231 1351 41289 1363
rect 41345 1539 41403 1551
rect 41345 1363 41357 1539
rect 41391 1363 41403 1539
rect 41345 1351 41403 1363
rect 41603 1539 41661 1551
rect 41603 1363 41615 1539
rect 41649 1363 41661 1539
rect 41603 1351 41661 1363
rect 41717 1539 41775 1551
rect 41717 1363 41729 1539
rect 41763 1363 41775 1539
rect 41717 1351 41775 1363
rect 41975 1539 42033 1551
rect 41975 1363 41987 1539
rect 42021 1363 42033 1539
rect 41975 1351 42033 1363
rect 42089 1539 42147 1551
rect 42089 1363 42101 1539
rect 42135 1363 42147 1539
rect 42089 1351 42147 1363
rect 42347 1539 42405 1551
rect 42347 1363 42359 1539
rect 42393 1363 42405 1539
rect 42347 1351 42405 1363
rect 42461 1539 42519 1551
rect 42461 1363 42473 1539
rect 42507 1363 42519 1539
rect 42461 1351 42519 1363
rect 42719 1539 42777 1551
rect 42719 1363 42731 1539
rect 42765 1363 42777 1539
rect 42719 1351 42777 1363
rect 42833 1539 42891 1551
rect 42833 1363 42845 1539
rect 42879 1363 42891 1539
rect 42833 1351 42891 1363
rect 43091 1539 43149 1551
rect 43091 1363 43103 1539
rect 43137 1363 43149 1539
rect 43091 1351 43149 1363
rect 43205 1539 43263 1551
rect 43205 1363 43217 1539
rect 43251 1363 43263 1539
rect 43205 1351 43263 1363
rect 43463 1539 43521 1551
rect 43463 1363 43475 1539
rect 43509 1363 43521 1539
rect 43463 1351 43521 1363
rect 43577 1539 43635 1551
rect 43577 1363 43589 1539
rect 43623 1363 43635 1539
rect 43577 1351 43635 1363
rect 43835 1539 43893 1551
rect 43835 1363 43847 1539
rect 43881 1363 43893 1539
rect 43835 1351 43893 1363
rect 43949 1539 44007 1551
rect 43949 1363 43961 1539
rect 43995 1363 44007 1539
rect 43949 1351 44007 1363
rect 44207 1539 44265 1551
rect 44207 1363 44219 1539
rect 44253 1363 44265 1539
rect 44207 1351 44265 1363
rect 44321 1539 44379 1551
rect 44321 1363 44333 1539
rect 44367 1363 44379 1539
rect 44321 1351 44379 1363
rect 44579 1539 44637 1551
rect 44579 1363 44591 1539
rect 44625 1363 44637 1539
rect 44579 1351 44637 1363
rect 44693 1539 44751 1551
rect 44693 1363 44705 1539
rect 44739 1363 44751 1539
rect 44693 1351 44751 1363
rect 44951 1539 45009 1551
rect 44951 1363 44963 1539
rect 44997 1363 45009 1539
rect 44951 1351 45009 1363
rect 45065 1539 45123 1551
rect 45065 1363 45077 1539
rect 45111 1363 45123 1539
rect 45065 1351 45123 1363
rect 45323 1539 45381 1551
rect 45323 1363 45335 1539
rect 45369 1363 45381 1539
rect 45323 1351 45381 1363
rect 45437 1539 45495 1551
rect 45437 1363 45449 1539
rect 45483 1363 45495 1539
rect 45437 1351 45495 1363
rect 45695 1539 45753 1551
rect 45695 1363 45707 1539
rect 45741 1363 45753 1539
rect 45695 1351 45753 1363
rect 45809 1539 45867 1551
rect 45809 1363 45821 1539
rect 45855 1363 45867 1539
rect 45809 1351 45867 1363
rect 46067 1539 46125 1551
rect 46067 1363 46079 1539
rect 46113 1363 46125 1539
rect 46067 1351 46125 1363
rect 46181 1539 46239 1551
rect 46181 1363 46193 1539
rect 46227 1363 46239 1539
rect 46181 1351 46239 1363
rect 46439 1539 46497 1551
rect 46439 1363 46451 1539
rect 46485 1363 46497 1539
rect 46439 1351 46497 1363
rect 46553 1539 46611 1551
rect 46553 1363 46565 1539
rect 46599 1363 46611 1539
rect 46553 1351 46611 1363
rect 46811 1539 46869 1551
rect 46811 1363 46823 1539
rect 46857 1363 46869 1539
rect 46811 1351 46869 1363
rect 46925 1539 46983 1551
rect 46925 1363 46937 1539
rect 46971 1363 46983 1539
rect 46925 1351 46983 1363
rect 47183 1539 47241 1551
rect 47183 1363 47195 1539
rect 47229 1363 47241 1539
rect 47183 1351 47241 1363
rect 47297 1539 47355 1551
rect 47297 1363 47309 1539
rect 47343 1363 47355 1539
rect 47297 1351 47355 1363
rect 47555 1539 47613 1551
rect 47555 1363 47567 1539
rect 47601 1363 47613 1539
rect 47555 1351 47613 1363
rect 47669 1539 47727 1551
rect 47669 1363 47681 1539
rect 47715 1363 47727 1539
rect 47669 1351 47727 1363
rect 47927 1539 47985 1551
rect 47927 1363 47939 1539
rect 47973 1363 47985 1539
rect 47927 1351 47985 1363
rect 48041 1539 48099 1551
rect 48041 1363 48053 1539
rect 48087 1363 48099 1539
rect 48041 1351 48099 1363
rect 48299 1539 48357 1551
rect 48299 1363 48311 1539
rect 48345 1363 48357 1539
rect 48299 1351 48357 1363
rect 39485 1121 39543 1133
rect 39485 945 39497 1121
rect 39531 945 39543 1121
rect 39485 933 39543 945
rect 39743 1121 39801 1133
rect 39743 945 39755 1121
rect 39789 945 39801 1121
rect 39743 933 39801 945
rect 39857 1121 39915 1133
rect 39857 945 39869 1121
rect 39903 945 39915 1121
rect 39857 933 39915 945
rect 40115 1121 40173 1133
rect 40115 945 40127 1121
rect 40161 945 40173 1121
rect 40115 933 40173 945
rect 40229 1121 40287 1133
rect 40229 945 40241 1121
rect 40275 945 40287 1121
rect 40229 933 40287 945
rect 40487 1121 40545 1133
rect 40487 945 40499 1121
rect 40533 945 40545 1121
rect 40487 933 40545 945
rect 40601 1121 40659 1133
rect 40601 945 40613 1121
rect 40647 945 40659 1121
rect 40601 933 40659 945
rect 40859 1121 40917 1133
rect 40859 945 40871 1121
rect 40905 945 40917 1121
rect 40859 933 40917 945
rect 40973 1121 41031 1133
rect 40973 945 40985 1121
rect 41019 945 41031 1121
rect 40973 933 41031 945
rect 41231 1121 41289 1133
rect 41231 945 41243 1121
rect 41277 945 41289 1121
rect 41231 933 41289 945
rect 41345 1121 41403 1133
rect 41345 945 41357 1121
rect 41391 945 41403 1121
rect 41345 933 41403 945
rect 41603 1121 41661 1133
rect 41603 945 41615 1121
rect 41649 945 41661 1121
rect 41603 933 41661 945
rect 41717 1121 41775 1133
rect 41717 945 41729 1121
rect 41763 945 41775 1121
rect 41717 933 41775 945
rect 41975 1121 42033 1133
rect 41975 945 41987 1121
rect 42021 945 42033 1121
rect 41975 933 42033 945
rect 42089 1121 42147 1133
rect 42089 945 42101 1121
rect 42135 945 42147 1121
rect 42089 933 42147 945
rect 42347 1121 42405 1133
rect 42347 945 42359 1121
rect 42393 945 42405 1121
rect 42347 933 42405 945
rect 42461 1121 42519 1133
rect 42461 945 42473 1121
rect 42507 945 42519 1121
rect 42461 933 42519 945
rect 42719 1121 42777 1133
rect 42719 945 42731 1121
rect 42765 945 42777 1121
rect 42719 933 42777 945
rect 42833 1121 42891 1133
rect 42833 945 42845 1121
rect 42879 945 42891 1121
rect 42833 933 42891 945
rect 43091 1121 43149 1133
rect 43091 945 43103 1121
rect 43137 945 43149 1121
rect 43091 933 43149 945
rect 43205 1121 43263 1133
rect 43205 945 43217 1121
rect 43251 945 43263 1121
rect 43205 933 43263 945
rect 43463 1121 43521 1133
rect 43463 945 43475 1121
rect 43509 945 43521 1121
rect 43463 933 43521 945
rect 43577 1121 43635 1133
rect 43577 945 43589 1121
rect 43623 945 43635 1121
rect 43577 933 43635 945
rect 43835 1121 43893 1133
rect 43835 945 43847 1121
rect 43881 945 43893 1121
rect 43835 933 43893 945
rect 43949 1121 44007 1133
rect 43949 945 43961 1121
rect 43995 945 44007 1121
rect 43949 933 44007 945
rect 44207 1121 44265 1133
rect 44207 945 44219 1121
rect 44253 945 44265 1121
rect 44207 933 44265 945
rect 44321 1121 44379 1133
rect 44321 945 44333 1121
rect 44367 945 44379 1121
rect 44321 933 44379 945
rect 44579 1121 44637 1133
rect 44579 945 44591 1121
rect 44625 945 44637 1121
rect 44579 933 44637 945
rect 44693 1121 44751 1133
rect 44693 945 44705 1121
rect 44739 945 44751 1121
rect 44693 933 44751 945
rect 44951 1121 45009 1133
rect 44951 945 44963 1121
rect 44997 945 45009 1121
rect 44951 933 45009 945
rect 45065 1121 45123 1133
rect 45065 945 45077 1121
rect 45111 945 45123 1121
rect 45065 933 45123 945
rect 45323 1121 45381 1133
rect 45323 945 45335 1121
rect 45369 945 45381 1121
rect 45323 933 45381 945
rect 45437 1121 45495 1133
rect 45437 945 45449 1121
rect 45483 945 45495 1121
rect 45437 933 45495 945
rect 45695 1121 45753 1133
rect 45695 945 45707 1121
rect 45741 945 45753 1121
rect 45695 933 45753 945
rect 45809 1121 45867 1133
rect 45809 945 45821 1121
rect 45855 945 45867 1121
rect 45809 933 45867 945
rect 46067 1121 46125 1133
rect 46067 945 46079 1121
rect 46113 945 46125 1121
rect 46067 933 46125 945
rect 46181 1121 46239 1133
rect 46181 945 46193 1121
rect 46227 945 46239 1121
rect 46181 933 46239 945
rect 46439 1121 46497 1133
rect 46439 945 46451 1121
rect 46485 945 46497 1121
rect 46439 933 46497 945
rect 46553 1121 46611 1133
rect 46553 945 46565 1121
rect 46599 945 46611 1121
rect 46553 933 46611 945
rect 46811 1121 46869 1133
rect 46811 945 46823 1121
rect 46857 945 46869 1121
rect 46811 933 46869 945
rect 46925 1121 46983 1133
rect 46925 945 46937 1121
rect 46971 945 46983 1121
rect 46925 933 46983 945
rect 47183 1121 47241 1133
rect 47183 945 47195 1121
rect 47229 945 47241 1121
rect 47183 933 47241 945
rect 47297 1121 47355 1133
rect 47297 945 47309 1121
rect 47343 945 47355 1121
rect 47297 933 47355 945
rect 47555 1121 47613 1133
rect 47555 945 47567 1121
rect 47601 945 47613 1121
rect 47555 933 47613 945
rect 47669 1121 47727 1133
rect 47669 945 47681 1121
rect 47715 945 47727 1121
rect 47669 933 47727 945
rect 47927 1121 47985 1133
rect 47927 945 47939 1121
rect 47973 945 47985 1121
rect 47927 933 47985 945
rect 48041 1121 48099 1133
rect 48041 945 48053 1121
rect 48087 945 48099 1121
rect 48041 933 48099 945
rect 48299 1121 48357 1133
rect 48299 945 48311 1121
rect 48345 945 48357 1121
rect 48299 933 48357 945
rect 39485 703 39543 715
rect 39485 527 39497 703
rect 39531 527 39543 703
rect 39485 515 39543 527
rect 39743 703 39801 715
rect 39743 527 39755 703
rect 39789 527 39801 703
rect 39743 515 39801 527
rect 39857 703 39915 715
rect 39857 527 39869 703
rect 39903 527 39915 703
rect 39857 515 39915 527
rect 40115 703 40173 715
rect 40115 527 40127 703
rect 40161 527 40173 703
rect 40115 515 40173 527
rect 40229 703 40287 715
rect 40229 527 40241 703
rect 40275 527 40287 703
rect 40229 515 40287 527
rect 40487 703 40545 715
rect 40487 527 40499 703
rect 40533 527 40545 703
rect 40487 515 40545 527
rect 40601 703 40659 715
rect 40601 527 40613 703
rect 40647 527 40659 703
rect 40601 515 40659 527
rect 40859 703 40917 715
rect 40859 527 40871 703
rect 40905 527 40917 703
rect 40859 515 40917 527
rect 40973 703 41031 715
rect 40973 527 40985 703
rect 41019 527 41031 703
rect 40973 515 41031 527
rect 41231 703 41289 715
rect 41231 527 41243 703
rect 41277 527 41289 703
rect 41231 515 41289 527
rect 41345 703 41403 715
rect 41345 527 41357 703
rect 41391 527 41403 703
rect 41345 515 41403 527
rect 41603 703 41661 715
rect 41603 527 41615 703
rect 41649 527 41661 703
rect 41603 515 41661 527
rect 41717 703 41775 715
rect 41717 527 41729 703
rect 41763 527 41775 703
rect 41717 515 41775 527
rect 41975 703 42033 715
rect 41975 527 41987 703
rect 42021 527 42033 703
rect 41975 515 42033 527
rect 42089 703 42147 715
rect 42089 527 42101 703
rect 42135 527 42147 703
rect 42089 515 42147 527
rect 42347 703 42405 715
rect 42347 527 42359 703
rect 42393 527 42405 703
rect 42347 515 42405 527
rect 42461 703 42519 715
rect 42461 527 42473 703
rect 42507 527 42519 703
rect 42461 515 42519 527
rect 42719 703 42777 715
rect 42719 527 42731 703
rect 42765 527 42777 703
rect 42719 515 42777 527
rect 42833 703 42891 715
rect 42833 527 42845 703
rect 42879 527 42891 703
rect 42833 515 42891 527
rect 43091 703 43149 715
rect 43091 527 43103 703
rect 43137 527 43149 703
rect 43091 515 43149 527
rect 43205 703 43263 715
rect 43205 527 43217 703
rect 43251 527 43263 703
rect 43205 515 43263 527
rect 43463 703 43521 715
rect 43463 527 43475 703
rect 43509 527 43521 703
rect 43463 515 43521 527
rect 43577 703 43635 715
rect 43577 527 43589 703
rect 43623 527 43635 703
rect 43577 515 43635 527
rect 43835 703 43893 715
rect 43835 527 43847 703
rect 43881 527 43893 703
rect 43835 515 43893 527
rect 43949 703 44007 715
rect 43949 527 43961 703
rect 43995 527 44007 703
rect 43949 515 44007 527
rect 44207 703 44265 715
rect 44207 527 44219 703
rect 44253 527 44265 703
rect 44207 515 44265 527
rect 44321 703 44379 715
rect 44321 527 44333 703
rect 44367 527 44379 703
rect 44321 515 44379 527
rect 44579 703 44637 715
rect 44579 527 44591 703
rect 44625 527 44637 703
rect 44579 515 44637 527
rect 44693 703 44751 715
rect 44693 527 44705 703
rect 44739 527 44751 703
rect 44693 515 44751 527
rect 44951 703 45009 715
rect 44951 527 44963 703
rect 44997 527 45009 703
rect 44951 515 45009 527
rect 45065 703 45123 715
rect 45065 527 45077 703
rect 45111 527 45123 703
rect 45065 515 45123 527
rect 45323 703 45381 715
rect 45323 527 45335 703
rect 45369 527 45381 703
rect 45323 515 45381 527
rect 45437 703 45495 715
rect 45437 527 45449 703
rect 45483 527 45495 703
rect 45437 515 45495 527
rect 45695 703 45753 715
rect 45695 527 45707 703
rect 45741 527 45753 703
rect 45695 515 45753 527
rect 45809 703 45867 715
rect 45809 527 45821 703
rect 45855 527 45867 703
rect 45809 515 45867 527
rect 46067 703 46125 715
rect 46067 527 46079 703
rect 46113 527 46125 703
rect 46067 515 46125 527
rect 46181 703 46239 715
rect 46181 527 46193 703
rect 46227 527 46239 703
rect 46181 515 46239 527
rect 46439 703 46497 715
rect 46439 527 46451 703
rect 46485 527 46497 703
rect 46439 515 46497 527
rect 46553 703 46611 715
rect 46553 527 46565 703
rect 46599 527 46611 703
rect 46553 515 46611 527
rect 46811 703 46869 715
rect 46811 527 46823 703
rect 46857 527 46869 703
rect 46811 515 46869 527
rect 46925 703 46983 715
rect 46925 527 46937 703
rect 46971 527 46983 703
rect 46925 515 46983 527
rect 47183 703 47241 715
rect 47183 527 47195 703
rect 47229 527 47241 703
rect 47183 515 47241 527
rect 47297 703 47355 715
rect 47297 527 47309 703
rect 47343 527 47355 703
rect 47297 515 47355 527
rect 47555 703 47613 715
rect 47555 527 47567 703
rect 47601 527 47613 703
rect 47555 515 47613 527
rect 47669 703 47727 715
rect 47669 527 47681 703
rect 47715 527 47727 703
rect 47669 515 47727 527
rect 47927 703 47985 715
rect 47927 527 47939 703
rect 47973 527 47985 703
rect 47927 515 47985 527
rect 48041 703 48099 715
rect 48041 527 48053 703
rect 48087 527 48099 703
rect 48041 515 48099 527
rect 48299 703 48357 715
rect 48299 527 48311 703
rect 48345 527 48357 703
rect 48299 515 48357 527
<< pdiff >>
rect 37997 9030 38055 9042
rect 37997 8654 38009 9030
rect 38043 8654 38055 9030
rect 37997 8642 38055 8654
rect 38255 9030 38313 9042
rect 38255 8654 38267 9030
rect 38301 8654 38313 9030
rect 38255 8642 38313 8654
rect 38369 9030 38427 9042
rect 38369 8654 38381 9030
rect 38415 8654 38427 9030
rect 38369 8642 38427 8654
rect 38627 9030 38685 9042
rect 38627 8654 38639 9030
rect 38673 8654 38685 9030
rect 38627 8642 38685 8654
rect 38741 9030 38799 9042
rect 38741 8654 38753 9030
rect 38787 8654 38799 9030
rect 38741 8642 38799 8654
rect 38999 9030 39057 9042
rect 38999 8654 39011 9030
rect 39045 8654 39057 9030
rect 38999 8642 39057 8654
rect 39113 9030 39171 9042
rect 39113 8654 39125 9030
rect 39159 8654 39171 9030
rect 39113 8642 39171 8654
rect 39371 9030 39429 9042
rect 39371 8654 39383 9030
rect 39417 8654 39429 9030
rect 39371 8642 39429 8654
rect 39485 9030 39543 9042
rect 39485 8654 39497 9030
rect 39531 8654 39543 9030
rect 39485 8642 39543 8654
rect 39743 9030 39801 9042
rect 39743 8654 39755 9030
rect 39789 8654 39801 9030
rect 39743 8642 39801 8654
rect 39857 9030 39915 9042
rect 39857 8654 39869 9030
rect 39903 8654 39915 9030
rect 39857 8642 39915 8654
rect 40115 9030 40173 9042
rect 40115 8654 40127 9030
rect 40161 8654 40173 9030
rect 40115 8642 40173 8654
rect 40229 9030 40287 9042
rect 40229 8654 40241 9030
rect 40275 8654 40287 9030
rect 40229 8642 40287 8654
rect 40487 9030 40545 9042
rect 40487 8654 40499 9030
rect 40533 8654 40545 9030
rect 40487 8642 40545 8654
rect 40601 9030 40659 9042
rect 40601 8654 40613 9030
rect 40647 8654 40659 9030
rect 40601 8642 40659 8654
rect 40859 9030 40917 9042
rect 40859 8654 40871 9030
rect 40905 8654 40917 9030
rect 40859 8642 40917 8654
rect 40973 9030 41031 9042
rect 40973 8654 40985 9030
rect 41019 8654 41031 9030
rect 40973 8642 41031 8654
rect 41231 9030 41289 9042
rect 41231 8654 41243 9030
rect 41277 8654 41289 9030
rect 41231 8642 41289 8654
rect 41345 9030 41403 9042
rect 41345 8654 41357 9030
rect 41391 8654 41403 9030
rect 41345 8642 41403 8654
rect 41603 9030 41661 9042
rect 41603 8654 41615 9030
rect 41649 8654 41661 9030
rect 41603 8642 41661 8654
rect 41717 9030 41775 9042
rect 41717 8654 41729 9030
rect 41763 8654 41775 9030
rect 41717 8642 41775 8654
rect 41975 9030 42033 9042
rect 41975 8654 41987 9030
rect 42021 8654 42033 9030
rect 41975 8642 42033 8654
rect 42089 9030 42147 9042
rect 42089 8654 42101 9030
rect 42135 8654 42147 9030
rect 42089 8642 42147 8654
rect 42347 9030 42405 9042
rect 42347 8654 42359 9030
rect 42393 8654 42405 9030
rect 42347 8642 42405 8654
rect 42461 9030 42519 9042
rect 42461 8654 42473 9030
rect 42507 8654 42519 9030
rect 42461 8642 42519 8654
rect 42719 9030 42777 9042
rect 42719 8654 42731 9030
rect 42765 8654 42777 9030
rect 42719 8642 42777 8654
rect 42833 9030 42891 9042
rect 42833 8654 42845 9030
rect 42879 8654 42891 9030
rect 42833 8642 42891 8654
rect 43091 9030 43149 9042
rect 43091 8654 43103 9030
rect 43137 8654 43149 9030
rect 43091 8642 43149 8654
rect 43205 9030 43263 9042
rect 43205 8654 43217 9030
rect 43251 8654 43263 9030
rect 43205 8642 43263 8654
rect 43463 9030 43521 9042
rect 43463 8654 43475 9030
rect 43509 8654 43521 9030
rect 43463 8642 43521 8654
rect 43577 9030 43635 9042
rect 43577 8654 43589 9030
rect 43623 8654 43635 9030
rect 43577 8642 43635 8654
rect 43835 9030 43893 9042
rect 43835 8654 43847 9030
rect 43881 8654 43893 9030
rect 43835 8642 43893 8654
rect 43949 9030 44007 9042
rect 43949 8654 43961 9030
rect 43995 8654 44007 9030
rect 43949 8642 44007 8654
rect 44207 9030 44265 9042
rect 44207 8654 44219 9030
rect 44253 8654 44265 9030
rect 44207 8642 44265 8654
rect 44321 9030 44379 9042
rect 44321 8654 44333 9030
rect 44367 8654 44379 9030
rect 44321 8642 44379 8654
rect 44579 9030 44637 9042
rect 44579 8654 44591 9030
rect 44625 8654 44637 9030
rect 44579 8642 44637 8654
rect 44693 9030 44751 9042
rect 44693 8654 44705 9030
rect 44739 8654 44751 9030
rect 44693 8642 44751 8654
rect 44951 9030 45009 9042
rect 44951 8654 44963 9030
rect 44997 8654 45009 9030
rect 44951 8642 45009 8654
rect 45065 9030 45123 9042
rect 45065 8654 45077 9030
rect 45111 8654 45123 9030
rect 45065 8642 45123 8654
rect 45323 9030 45381 9042
rect 45323 8654 45335 9030
rect 45369 8654 45381 9030
rect 45323 8642 45381 8654
rect 45437 9030 45495 9042
rect 45437 8654 45449 9030
rect 45483 8654 45495 9030
rect 45437 8642 45495 8654
rect 45695 9030 45753 9042
rect 45695 8654 45707 9030
rect 45741 8654 45753 9030
rect 45695 8642 45753 8654
rect 45809 9030 45867 9042
rect 45809 8654 45821 9030
rect 45855 8654 45867 9030
rect 45809 8642 45867 8654
rect 46067 9030 46125 9042
rect 46067 8654 46079 9030
rect 46113 8654 46125 9030
rect 46067 8642 46125 8654
rect 46181 9030 46239 9042
rect 46181 8654 46193 9030
rect 46227 8654 46239 9030
rect 46181 8642 46239 8654
rect 46439 9030 46497 9042
rect 46439 8654 46451 9030
rect 46485 8654 46497 9030
rect 46439 8642 46497 8654
rect 46553 9030 46611 9042
rect 46553 8654 46565 9030
rect 46599 8654 46611 9030
rect 46553 8642 46611 8654
rect 46811 9030 46869 9042
rect 46811 8654 46823 9030
rect 46857 8654 46869 9030
rect 46811 8642 46869 8654
rect 46925 9030 46983 9042
rect 46925 8654 46937 9030
rect 46971 8654 46983 9030
rect 46925 8642 46983 8654
rect 47183 9030 47241 9042
rect 47183 8654 47195 9030
rect 47229 8654 47241 9030
rect 47183 8642 47241 8654
rect 47297 9030 47355 9042
rect 47297 8654 47309 9030
rect 47343 8654 47355 9030
rect 47297 8642 47355 8654
rect 47555 9030 47613 9042
rect 47555 8654 47567 9030
rect 47601 8654 47613 9030
rect 47555 8642 47613 8654
rect 47669 9030 47727 9042
rect 47669 8654 47681 9030
rect 47715 8654 47727 9030
rect 47669 8642 47727 8654
rect 47927 9030 47985 9042
rect 47927 8654 47939 9030
rect 47973 8654 47985 9030
rect 47927 8642 47985 8654
rect 48041 9030 48099 9042
rect 48041 8654 48053 9030
rect 48087 8654 48099 9030
rect 48041 8642 48099 8654
rect 48299 9030 48357 9042
rect 48299 8654 48311 9030
rect 48345 8654 48357 9030
rect 48299 8642 48357 8654
rect 48413 9030 48471 9042
rect 48413 8654 48425 9030
rect 48459 8654 48471 9030
rect 48413 8642 48471 8654
rect 48671 9030 48729 9042
rect 48671 8654 48683 9030
rect 48717 8654 48729 9030
rect 48671 8642 48729 8654
rect 48785 9030 48843 9042
rect 48785 8654 48797 9030
rect 48831 8654 48843 9030
rect 48785 8642 48843 8654
rect 49043 9030 49101 9042
rect 49043 8654 49055 9030
rect 49089 8654 49101 9030
rect 49043 8642 49101 8654
rect 49157 9030 49215 9042
rect 49157 8654 49169 9030
rect 49203 8654 49215 9030
rect 49157 8642 49215 8654
rect 49415 9030 49473 9042
rect 49415 8654 49427 9030
rect 49461 8654 49473 9030
rect 49415 8642 49473 8654
rect 49529 9030 49587 9042
rect 49529 8654 49541 9030
rect 49575 8654 49587 9030
rect 49529 8642 49587 8654
rect 49787 9030 49845 9042
rect 49787 8654 49799 9030
rect 49833 8654 49845 9030
rect 49787 8642 49845 8654
rect 37997 8394 38055 8406
rect 37997 8018 38009 8394
rect 38043 8018 38055 8394
rect 37997 8006 38055 8018
rect 38255 8394 38313 8406
rect 38255 8018 38267 8394
rect 38301 8018 38313 8394
rect 38255 8006 38313 8018
rect 38369 8394 38427 8406
rect 38369 8018 38381 8394
rect 38415 8018 38427 8394
rect 38369 8006 38427 8018
rect 38627 8394 38685 8406
rect 38627 8018 38639 8394
rect 38673 8018 38685 8394
rect 38627 8006 38685 8018
rect 38741 8394 38799 8406
rect 38741 8018 38753 8394
rect 38787 8018 38799 8394
rect 38741 8006 38799 8018
rect 38999 8394 39057 8406
rect 38999 8018 39011 8394
rect 39045 8018 39057 8394
rect 38999 8006 39057 8018
rect 39113 8394 39171 8406
rect 39113 8018 39125 8394
rect 39159 8018 39171 8394
rect 39113 8006 39171 8018
rect 39371 8394 39429 8406
rect 39371 8018 39383 8394
rect 39417 8018 39429 8394
rect 39371 8006 39429 8018
rect 39485 8394 39543 8406
rect 39485 8018 39497 8394
rect 39531 8018 39543 8394
rect 39485 8006 39543 8018
rect 39743 8394 39801 8406
rect 39743 8018 39755 8394
rect 39789 8018 39801 8394
rect 39743 8006 39801 8018
rect 39857 8394 39915 8406
rect 39857 8018 39869 8394
rect 39903 8018 39915 8394
rect 39857 8006 39915 8018
rect 40115 8394 40173 8406
rect 40115 8018 40127 8394
rect 40161 8018 40173 8394
rect 40115 8006 40173 8018
rect 40229 8394 40287 8406
rect 40229 8018 40241 8394
rect 40275 8018 40287 8394
rect 40229 8006 40287 8018
rect 40487 8394 40545 8406
rect 40487 8018 40499 8394
rect 40533 8018 40545 8394
rect 40487 8006 40545 8018
rect 40601 8394 40659 8406
rect 40601 8018 40613 8394
rect 40647 8018 40659 8394
rect 40601 8006 40659 8018
rect 40859 8394 40917 8406
rect 40859 8018 40871 8394
rect 40905 8018 40917 8394
rect 40859 8006 40917 8018
rect 40973 8394 41031 8406
rect 40973 8018 40985 8394
rect 41019 8018 41031 8394
rect 40973 8006 41031 8018
rect 41231 8394 41289 8406
rect 41231 8018 41243 8394
rect 41277 8018 41289 8394
rect 41231 8006 41289 8018
rect 41345 8394 41403 8406
rect 41345 8018 41357 8394
rect 41391 8018 41403 8394
rect 41345 8006 41403 8018
rect 41603 8394 41661 8406
rect 41603 8018 41615 8394
rect 41649 8018 41661 8394
rect 41603 8006 41661 8018
rect 41717 8394 41775 8406
rect 41717 8018 41729 8394
rect 41763 8018 41775 8394
rect 41717 8006 41775 8018
rect 41975 8394 42033 8406
rect 41975 8018 41987 8394
rect 42021 8018 42033 8394
rect 41975 8006 42033 8018
rect 42089 8394 42147 8406
rect 42089 8018 42101 8394
rect 42135 8018 42147 8394
rect 42089 8006 42147 8018
rect 42347 8394 42405 8406
rect 42347 8018 42359 8394
rect 42393 8018 42405 8394
rect 42347 8006 42405 8018
rect 42461 8394 42519 8406
rect 42461 8018 42473 8394
rect 42507 8018 42519 8394
rect 42461 8006 42519 8018
rect 42719 8394 42777 8406
rect 42719 8018 42731 8394
rect 42765 8018 42777 8394
rect 42719 8006 42777 8018
rect 42833 8394 42891 8406
rect 42833 8018 42845 8394
rect 42879 8018 42891 8394
rect 42833 8006 42891 8018
rect 43091 8394 43149 8406
rect 43091 8018 43103 8394
rect 43137 8018 43149 8394
rect 43091 8006 43149 8018
rect 43205 8394 43263 8406
rect 43205 8018 43217 8394
rect 43251 8018 43263 8394
rect 43205 8006 43263 8018
rect 43463 8394 43521 8406
rect 43463 8018 43475 8394
rect 43509 8018 43521 8394
rect 43463 8006 43521 8018
rect 43577 8394 43635 8406
rect 43577 8018 43589 8394
rect 43623 8018 43635 8394
rect 43577 8006 43635 8018
rect 43835 8394 43893 8406
rect 43835 8018 43847 8394
rect 43881 8018 43893 8394
rect 43835 8006 43893 8018
rect 43949 8394 44007 8406
rect 43949 8018 43961 8394
rect 43995 8018 44007 8394
rect 43949 8006 44007 8018
rect 44207 8394 44265 8406
rect 44207 8018 44219 8394
rect 44253 8018 44265 8394
rect 44207 8006 44265 8018
rect 44321 8394 44379 8406
rect 44321 8018 44333 8394
rect 44367 8018 44379 8394
rect 44321 8006 44379 8018
rect 44579 8394 44637 8406
rect 44579 8018 44591 8394
rect 44625 8018 44637 8394
rect 44579 8006 44637 8018
rect 44693 8394 44751 8406
rect 44693 8018 44705 8394
rect 44739 8018 44751 8394
rect 44693 8006 44751 8018
rect 44951 8394 45009 8406
rect 44951 8018 44963 8394
rect 44997 8018 45009 8394
rect 44951 8006 45009 8018
rect 45065 8394 45123 8406
rect 45065 8018 45077 8394
rect 45111 8018 45123 8394
rect 45065 8006 45123 8018
rect 45323 8394 45381 8406
rect 45323 8018 45335 8394
rect 45369 8018 45381 8394
rect 45323 8006 45381 8018
rect 45437 8394 45495 8406
rect 45437 8018 45449 8394
rect 45483 8018 45495 8394
rect 45437 8006 45495 8018
rect 45695 8394 45753 8406
rect 45695 8018 45707 8394
rect 45741 8018 45753 8394
rect 45695 8006 45753 8018
rect 45809 8394 45867 8406
rect 45809 8018 45821 8394
rect 45855 8018 45867 8394
rect 45809 8006 45867 8018
rect 46067 8394 46125 8406
rect 46067 8018 46079 8394
rect 46113 8018 46125 8394
rect 46067 8006 46125 8018
rect 46181 8394 46239 8406
rect 46181 8018 46193 8394
rect 46227 8018 46239 8394
rect 46181 8006 46239 8018
rect 46439 8394 46497 8406
rect 46439 8018 46451 8394
rect 46485 8018 46497 8394
rect 46439 8006 46497 8018
rect 46553 8394 46611 8406
rect 46553 8018 46565 8394
rect 46599 8018 46611 8394
rect 46553 8006 46611 8018
rect 46811 8394 46869 8406
rect 46811 8018 46823 8394
rect 46857 8018 46869 8394
rect 46811 8006 46869 8018
rect 46925 8394 46983 8406
rect 46925 8018 46937 8394
rect 46971 8018 46983 8394
rect 46925 8006 46983 8018
rect 47183 8394 47241 8406
rect 47183 8018 47195 8394
rect 47229 8018 47241 8394
rect 47183 8006 47241 8018
rect 47297 8394 47355 8406
rect 47297 8018 47309 8394
rect 47343 8018 47355 8394
rect 47297 8006 47355 8018
rect 47555 8394 47613 8406
rect 47555 8018 47567 8394
rect 47601 8018 47613 8394
rect 47555 8006 47613 8018
rect 47669 8394 47727 8406
rect 47669 8018 47681 8394
rect 47715 8018 47727 8394
rect 47669 8006 47727 8018
rect 47927 8394 47985 8406
rect 47927 8018 47939 8394
rect 47973 8018 47985 8394
rect 47927 8006 47985 8018
rect 48041 8394 48099 8406
rect 48041 8018 48053 8394
rect 48087 8018 48099 8394
rect 48041 8006 48099 8018
rect 48299 8394 48357 8406
rect 48299 8018 48311 8394
rect 48345 8018 48357 8394
rect 48299 8006 48357 8018
rect 48413 8394 48471 8406
rect 48413 8018 48425 8394
rect 48459 8018 48471 8394
rect 48413 8006 48471 8018
rect 48671 8394 48729 8406
rect 48671 8018 48683 8394
rect 48717 8018 48729 8394
rect 48671 8006 48729 8018
rect 48785 8394 48843 8406
rect 48785 8018 48797 8394
rect 48831 8018 48843 8394
rect 48785 8006 48843 8018
rect 49043 8394 49101 8406
rect 49043 8018 49055 8394
rect 49089 8018 49101 8394
rect 49043 8006 49101 8018
rect 49157 8394 49215 8406
rect 49157 8018 49169 8394
rect 49203 8018 49215 8394
rect 49157 8006 49215 8018
rect 49415 8394 49473 8406
rect 49415 8018 49427 8394
rect 49461 8018 49473 8394
rect 49415 8006 49473 8018
rect 49529 8394 49587 8406
rect 49529 8018 49541 8394
rect 49575 8018 49587 8394
rect 49529 8006 49587 8018
rect 49787 8394 49845 8406
rect 49787 8018 49799 8394
rect 49833 8018 49845 8394
rect 49787 8006 49845 8018
rect 37997 7758 38055 7770
rect 37997 7382 38009 7758
rect 38043 7382 38055 7758
rect 37997 7370 38055 7382
rect 38255 7758 38313 7770
rect 38255 7382 38267 7758
rect 38301 7382 38313 7758
rect 38255 7370 38313 7382
rect 38369 7758 38427 7770
rect 38369 7382 38381 7758
rect 38415 7382 38427 7758
rect 38369 7370 38427 7382
rect 38627 7758 38685 7770
rect 38627 7382 38639 7758
rect 38673 7382 38685 7758
rect 38627 7370 38685 7382
rect 38741 7758 38799 7770
rect 38741 7382 38753 7758
rect 38787 7382 38799 7758
rect 38741 7370 38799 7382
rect 38999 7758 39057 7770
rect 38999 7382 39011 7758
rect 39045 7382 39057 7758
rect 38999 7370 39057 7382
rect 39113 7758 39171 7770
rect 39113 7382 39125 7758
rect 39159 7382 39171 7758
rect 39113 7370 39171 7382
rect 39371 7758 39429 7770
rect 39371 7382 39383 7758
rect 39417 7382 39429 7758
rect 39371 7370 39429 7382
rect 39485 7758 39543 7770
rect 39485 7382 39497 7758
rect 39531 7382 39543 7758
rect 39485 7370 39543 7382
rect 39743 7758 39801 7770
rect 39743 7382 39755 7758
rect 39789 7382 39801 7758
rect 39743 7370 39801 7382
rect 39857 7758 39915 7770
rect 39857 7382 39869 7758
rect 39903 7382 39915 7758
rect 39857 7370 39915 7382
rect 40115 7758 40173 7770
rect 40115 7382 40127 7758
rect 40161 7382 40173 7758
rect 40115 7370 40173 7382
rect 40229 7758 40287 7770
rect 40229 7382 40241 7758
rect 40275 7382 40287 7758
rect 40229 7370 40287 7382
rect 40487 7758 40545 7770
rect 40487 7382 40499 7758
rect 40533 7382 40545 7758
rect 40487 7370 40545 7382
rect 40601 7758 40659 7770
rect 40601 7382 40613 7758
rect 40647 7382 40659 7758
rect 40601 7370 40659 7382
rect 40859 7758 40917 7770
rect 40859 7382 40871 7758
rect 40905 7382 40917 7758
rect 40859 7370 40917 7382
rect 40973 7758 41031 7770
rect 40973 7382 40985 7758
rect 41019 7382 41031 7758
rect 40973 7370 41031 7382
rect 41231 7758 41289 7770
rect 41231 7382 41243 7758
rect 41277 7382 41289 7758
rect 41231 7370 41289 7382
rect 41345 7758 41403 7770
rect 41345 7382 41357 7758
rect 41391 7382 41403 7758
rect 41345 7370 41403 7382
rect 41603 7758 41661 7770
rect 41603 7382 41615 7758
rect 41649 7382 41661 7758
rect 41603 7370 41661 7382
rect 41717 7758 41775 7770
rect 41717 7382 41729 7758
rect 41763 7382 41775 7758
rect 41717 7370 41775 7382
rect 41975 7758 42033 7770
rect 41975 7382 41987 7758
rect 42021 7382 42033 7758
rect 41975 7370 42033 7382
rect 42089 7758 42147 7770
rect 42089 7382 42101 7758
rect 42135 7382 42147 7758
rect 42089 7370 42147 7382
rect 42347 7758 42405 7770
rect 42347 7382 42359 7758
rect 42393 7382 42405 7758
rect 42347 7370 42405 7382
rect 42461 7758 42519 7770
rect 42461 7382 42473 7758
rect 42507 7382 42519 7758
rect 42461 7370 42519 7382
rect 42719 7758 42777 7770
rect 42719 7382 42731 7758
rect 42765 7382 42777 7758
rect 42719 7370 42777 7382
rect 42833 7758 42891 7770
rect 42833 7382 42845 7758
rect 42879 7382 42891 7758
rect 42833 7370 42891 7382
rect 43091 7758 43149 7770
rect 43091 7382 43103 7758
rect 43137 7382 43149 7758
rect 43091 7370 43149 7382
rect 43205 7758 43263 7770
rect 43205 7382 43217 7758
rect 43251 7382 43263 7758
rect 43205 7370 43263 7382
rect 43463 7758 43521 7770
rect 43463 7382 43475 7758
rect 43509 7382 43521 7758
rect 43463 7370 43521 7382
rect 43577 7758 43635 7770
rect 43577 7382 43589 7758
rect 43623 7382 43635 7758
rect 43577 7370 43635 7382
rect 43835 7758 43893 7770
rect 43835 7382 43847 7758
rect 43881 7382 43893 7758
rect 43835 7370 43893 7382
rect 43949 7758 44007 7770
rect 43949 7382 43961 7758
rect 43995 7382 44007 7758
rect 43949 7370 44007 7382
rect 44207 7758 44265 7770
rect 44207 7382 44219 7758
rect 44253 7382 44265 7758
rect 44207 7370 44265 7382
rect 44321 7758 44379 7770
rect 44321 7382 44333 7758
rect 44367 7382 44379 7758
rect 44321 7370 44379 7382
rect 44579 7758 44637 7770
rect 44579 7382 44591 7758
rect 44625 7382 44637 7758
rect 44579 7370 44637 7382
rect 44693 7758 44751 7770
rect 44693 7382 44705 7758
rect 44739 7382 44751 7758
rect 44693 7370 44751 7382
rect 44951 7758 45009 7770
rect 44951 7382 44963 7758
rect 44997 7382 45009 7758
rect 44951 7370 45009 7382
rect 45065 7758 45123 7770
rect 45065 7382 45077 7758
rect 45111 7382 45123 7758
rect 45065 7370 45123 7382
rect 45323 7758 45381 7770
rect 45323 7382 45335 7758
rect 45369 7382 45381 7758
rect 45323 7370 45381 7382
rect 45437 7758 45495 7770
rect 45437 7382 45449 7758
rect 45483 7382 45495 7758
rect 45437 7370 45495 7382
rect 45695 7758 45753 7770
rect 45695 7382 45707 7758
rect 45741 7382 45753 7758
rect 45695 7370 45753 7382
rect 45809 7758 45867 7770
rect 45809 7382 45821 7758
rect 45855 7382 45867 7758
rect 45809 7370 45867 7382
rect 46067 7758 46125 7770
rect 46067 7382 46079 7758
rect 46113 7382 46125 7758
rect 46067 7370 46125 7382
rect 46181 7758 46239 7770
rect 46181 7382 46193 7758
rect 46227 7382 46239 7758
rect 46181 7370 46239 7382
rect 46439 7758 46497 7770
rect 46439 7382 46451 7758
rect 46485 7382 46497 7758
rect 46439 7370 46497 7382
rect 46553 7758 46611 7770
rect 46553 7382 46565 7758
rect 46599 7382 46611 7758
rect 46553 7370 46611 7382
rect 46811 7758 46869 7770
rect 46811 7382 46823 7758
rect 46857 7382 46869 7758
rect 46811 7370 46869 7382
rect 46925 7758 46983 7770
rect 46925 7382 46937 7758
rect 46971 7382 46983 7758
rect 46925 7370 46983 7382
rect 47183 7758 47241 7770
rect 47183 7382 47195 7758
rect 47229 7382 47241 7758
rect 47183 7370 47241 7382
rect 47297 7758 47355 7770
rect 47297 7382 47309 7758
rect 47343 7382 47355 7758
rect 47297 7370 47355 7382
rect 47555 7758 47613 7770
rect 47555 7382 47567 7758
rect 47601 7382 47613 7758
rect 47555 7370 47613 7382
rect 47669 7758 47727 7770
rect 47669 7382 47681 7758
rect 47715 7382 47727 7758
rect 47669 7370 47727 7382
rect 47927 7758 47985 7770
rect 47927 7382 47939 7758
rect 47973 7382 47985 7758
rect 47927 7370 47985 7382
rect 48041 7758 48099 7770
rect 48041 7382 48053 7758
rect 48087 7382 48099 7758
rect 48041 7370 48099 7382
rect 48299 7758 48357 7770
rect 48299 7382 48311 7758
rect 48345 7382 48357 7758
rect 48299 7370 48357 7382
rect 48413 7758 48471 7770
rect 48413 7382 48425 7758
rect 48459 7382 48471 7758
rect 48413 7370 48471 7382
rect 48671 7758 48729 7770
rect 48671 7382 48683 7758
rect 48717 7382 48729 7758
rect 48671 7370 48729 7382
rect 48785 7758 48843 7770
rect 48785 7382 48797 7758
rect 48831 7382 48843 7758
rect 48785 7370 48843 7382
rect 49043 7758 49101 7770
rect 49043 7382 49055 7758
rect 49089 7382 49101 7758
rect 49043 7370 49101 7382
rect 49157 7758 49215 7770
rect 49157 7382 49169 7758
rect 49203 7382 49215 7758
rect 49157 7370 49215 7382
rect 49415 7758 49473 7770
rect 49415 7382 49427 7758
rect 49461 7382 49473 7758
rect 49415 7370 49473 7382
rect 49529 7758 49587 7770
rect 49529 7382 49541 7758
rect 49575 7382 49587 7758
rect 49529 7370 49587 7382
rect 49787 7758 49845 7770
rect 49787 7382 49799 7758
rect 49833 7382 49845 7758
rect 49787 7370 49845 7382
rect 39485 6642 39543 6654
rect 39485 5866 39497 6642
rect 39531 5866 39543 6642
rect 39485 5854 39543 5866
rect 39743 6642 39801 6654
rect 39743 5866 39755 6642
rect 39789 5866 39801 6642
rect 39743 5854 39801 5866
rect 39857 6642 39915 6654
rect 39857 5866 39869 6642
rect 39903 5866 39915 6642
rect 39857 5854 39915 5866
rect 40115 6642 40173 6654
rect 40115 5866 40127 6642
rect 40161 5866 40173 6642
rect 40115 5854 40173 5866
rect 40229 6642 40287 6654
rect 40229 5866 40241 6642
rect 40275 5866 40287 6642
rect 40229 5854 40287 5866
rect 40487 6642 40545 6654
rect 40487 5866 40499 6642
rect 40533 5866 40545 6642
rect 40487 5854 40545 5866
rect 40601 6642 40659 6654
rect 40601 5866 40613 6642
rect 40647 5866 40659 6642
rect 40601 5854 40659 5866
rect 40859 6642 40917 6654
rect 40859 5866 40871 6642
rect 40905 5866 40917 6642
rect 40859 5854 40917 5866
rect 40973 6642 41031 6654
rect 40973 5866 40985 6642
rect 41019 5866 41031 6642
rect 40973 5854 41031 5866
rect 41231 6642 41289 6654
rect 41231 5866 41243 6642
rect 41277 5866 41289 6642
rect 41231 5854 41289 5866
rect 41345 6642 41403 6654
rect 41345 5866 41357 6642
rect 41391 5866 41403 6642
rect 41345 5854 41403 5866
rect 41603 6642 41661 6654
rect 41603 5866 41615 6642
rect 41649 5866 41661 6642
rect 41603 5854 41661 5866
rect 41717 6642 41775 6654
rect 41717 5866 41729 6642
rect 41763 5866 41775 6642
rect 41717 5854 41775 5866
rect 41975 6642 42033 6654
rect 41975 5866 41987 6642
rect 42021 5866 42033 6642
rect 41975 5854 42033 5866
rect 42089 6642 42147 6654
rect 42089 5866 42101 6642
rect 42135 5866 42147 6642
rect 42089 5854 42147 5866
rect 42347 6642 42405 6654
rect 42347 5866 42359 6642
rect 42393 5866 42405 6642
rect 42347 5854 42405 5866
rect 39485 5606 39543 5618
rect 39485 4830 39497 5606
rect 39531 4830 39543 5606
rect 39485 4818 39543 4830
rect 39743 5606 39801 5618
rect 39743 4830 39755 5606
rect 39789 4830 39801 5606
rect 39743 4818 39801 4830
rect 39857 5606 39915 5618
rect 39857 4830 39869 5606
rect 39903 4830 39915 5606
rect 39857 4818 39915 4830
rect 40115 5606 40173 5618
rect 40115 4830 40127 5606
rect 40161 4830 40173 5606
rect 40115 4818 40173 4830
rect 40229 5606 40287 5618
rect 40229 4830 40241 5606
rect 40275 4830 40287 5606
rect 40229 4818 40287 4830
rect 40487 5606 40545 5618
rect 40487 4830 40499 5606
rect 40533 4830 40545 5606
rect 40487 4818 40545 4830
rect 40601 5606 40659 5618
rect 40601 4830 40613 5606
rect 40647 4830 40659 5606
rect 40601 4818 40659 4830
rect 40859 5606 40917 5618
rect 40859 4830 40871 5606
rect 40905 4830 40917 5606
rect 40859 4818 40917 4830
rect 40973 5606 41031 5618
rect 40973 4830 40985 5606
rect 41019 4830 41031 5606
rect 40973 4818 41031 4830
rect 41231 5606 41289 5618
rect 41231 4830 41243 5606
rect 41277 4830 41289 5606
rect 41231 4818 41289 4830
rect 41345 5606 41403 5618
rect 41345 4830 41357 5606
rect 41391 4830 41403 5606
rect 41345 4818 41403 4830
rect 41603 5606 41661 5618
rect 41603 4830 41615 5606
rect 41649 4830 41661 5606
rect 41603 4818 41661 4830
rect 41717 5606 41775 5618
rect 41717 4830 41729 5606
rect 41763 4830 41775 5606
rect 41717 4818 41775 4830
rect 41975 5606 42033 5618
rect 41975 4830 41987 5606
rect 42021 4830 42033 5606
rect 41975 4818 42033 4830
rect 42089 5606 42147 5618
rect 42089 4830 42101 5606
rect 42135 4830 42147 5606
rect 42089 4818 42147 4830
rect 42347 5606 42405 5618
rect 42347 4830 42359 5606
rect 42393 4830 42405 5606
rect 42347 4818 42405 4830
rect 39485 4570 39543 4582
rect 39485 3794 39497 4570
rect 39531 3794 39543 4570
rect 39485 3782 39543 3794
rect 39743 4570 39801 4582
rect 39743 3794 39755 4570
rect 39789 3794 39801 4570
rect 39743 3782 39801 3794
rect 39857 4570 39915 4582
rect 39857 3794 39869 4570
rect 39903 3794 39915 4570
rect 39857 3782 39915 3794
rect 40115 4570 40173 4582
rect 40115 3794 40127 4570
rect 40161 3794 40173 4570
rect 40115 3782 40173 3794
rect 40229 4570 40287 4582
rect 40229 3794 40241 4570
rect 40275 3794 40287 4570
rect 40229 3782 40287 3794
rect 40487 4570 40545 4582
rect 40487 3794 40499 4570
rect 40533 3794 40545 4570
rect 40487 3782 40545 3794
rect 40601 4570 40659 4582
rect 40601 3794 40613 4570
rect 40647 3794 40659 4570
rect 40601 3782 40659 3794
rect 40859 4570 40917 4582
rect 40859 3794 40871 4570
rect 40905 3794 40917 4570
rect 40859 3782 40917 3794
rect 40973 4570 41031 4582
rect 40973 3794 40985 4570
rect 41019 3794 41031 4570
rect 40973 3782 41031 3794
rect 41231 4570 41289 4582
rect 41231 3794 41243 4570
rect 41277 3794 41289 4570
rect 41231 3782 41289 3794
rect 41345 4570 41403 4582
rect 41345 3794 41357 4570
rect 41391 3794 41403 4570
rect 41345 3782 41403 3794
rect 41603 4570 41661 4582
rect 41603 3794 41615 4570
rect 41649 3794 41661 4570
rect 41603 3782 41661 3794
rect 41717 4570 41775 4582
rect 41717 3794 41729 4570
rect 41763 3794 41775 4570
rect 41717 3782 41775 3794
rect 41975 4570 42033 4582
rect 41975 3794 41987 4570
rect 42021 3794 42033 4570
rect 41975 3782 42033 3794
rect 42089 4570 42147 4582
rect 42089 3794 42101 4570
rect 42135 3794 42147 4570
rect 42089 3782 42147 3794
rect 42347 4570 42405 4582
rect 42347 3794 42359 4570
rect 42393 3794 42405 4570
rect 42347 3782 42405 3794
rect 39485 3534 39543 3546
rect 39485 2758 39497 3534
rect 39531 2758 39543 3534
rect 39485 2746 39543 2758
rect 39743 3534 39801 3546
rect 39743 2758 39755 3534
rect 39789 2758 39801 3534
rect 39743 2746 39801 2758
rect 39857 3534 39915 3546
rect 39857 2758 39869 3534
rect 39903 2758 39915 3534
rect 39857 2746 39915 2758
rect 40115 3534 40173 3546
rect 40115 2758 40127 3534
rect 40161 2758 40173 3534
rect 40115 2746 40173 2758
rect 40229 3534 40287 3546
rect 40229 2758 40241 3534
rect 40275 2758 40287 3534
rect 40229 2746 40287 2758
rect 40487 3534 40545 3546
rect 40487 2758 40499 3534
rect 40533 2758 40545 3534
rect 40487 2746 40545 2758
rect 40601 3534 40659 3546
rect 40601 2758 40613 3534
rect 40647 2758 40659 3534
rect 40601 2746 40659 2758
rect 40859 3534 40917 3546
rect 40859 2758 40871 3534
rect 40905 2758 40917 3534
rect 40859 2746 40917 2758
rect 40973 3534 41031 3546
rect 40973 2758 40985 3534
rect 41019 2758 41031 3534
rect 40973 2746 41031 2758
rect 41231 3534 41289 3546
rect 41231 2758 41243 3534
rect 41277 2758 41289 3534
rect 41231 2746 41289 2758
rect 41345 3534 41403 3546
rect 41345 2758 41357 3534
rect 41391 2758 41403 3534
rect 41345 2746 41403 2758
rect 41603 3534 41661 3546
rect 41603 2758 41615 3534
rect 41649 2758 41661 3534
rect 41603 2746 41661 2758
rect 41717 3534 41775 3546
rect 41717 2758 41729 3534
rect 41763 2758 41775 3534
rect 41717 2746 41775 2758
rect 41975 3534 42033 3546
rect 41975 2758 41987 3534
rect 42021 2758 42033 3534
rect 41975 2746 42033 2758
rect 42089 3534 42147 3546
rect 42089 2758 42101 3534
rect 42135 2758 42147 3534
rect 42089 2746 42147 2758
rect 42347 3534 42405 3546
rect 42347 2758 42359 3534
rect 42393 2758 42405 3534
rect 42347 2746 42405 2758
<< ndiffc >>
rect 39497 1781 39531 1957
rect 39755 1781 39789 1957
rect 39869 1781 39903 1957
rect 40127 1781 40161 1957
rect 40241 1781 40275 1957
rect 40499 1781 40533 1957
rect 40613 1781 40647 1957
rect 40871 1781 40905 1957
rect 40985 1781 41019 1957
rect 41243 1781 41277 1957
rect 41357 1781 41391 1957
rect 41615 1781 41649 1957
rect 41729 1781 41763 1957
rect 41987 1781 42021 1957
rect 42101 1781 42135 1957
rect 42359 1781 42393 1957
rect 42473 1781 42507 1957
rect 42731 1781 42765 1957
rect 42845 1781 42879 1957
rect 43103 1781 43137 1957
rect 43217 1781 43251 1957
rect 43475 1781 43509 1957
rect 43589 1781 43623 1957
rect 43847 1781 43881 1957
rect 43961 1781 43995 1957
rect 44219 1781 44253 1957
rect 44333 1781 44367 1957
rect 44591 1781 44625 1957
rect 44705 1781 44739 1957
rect 44963 1781 44997 1957
rect 45077 1781 45111 1957
rect 45335 1781 45369 1957
rect 45449 1781 45483 1957
rect 45707 1781 45741 1957
rect 45821 1781 45855 1957
rect 46079 1781 46113 1957
rect 46193 1781 46227 1957
rect 46451 1781 46485 1957
rect 46565 1781 46599 1957
rect 46823 1781 46857 1957
rect 46937 1781 46971 1957
rect 47195 1781 47229 1957
rect 47309 1781 47343 1957
rect 47567 1781 47601 1957
rect 47681 1781 47715 1957
rect 47939 1781 47973 1957
rect 48053 1781 48087 1957
rect 48311 1781 48345 1957
rect 39497 1363 39531 1539
rect 39755 1363 39789 1539
rect 39869 1363 39903 1539
rect 40127 1363 40161 1539
rect 40241 1363 40275 1539
rect 40499 1363 40533 1539
rect 40613 1363 40647 1539
rect 40871 1363 40905 1539
rect 40985 1363 41019 1539
rect 41243 1363 41277 1539
rect 41357 1363 41391 1539
rect 41615 1363 41649 1539
rect 41729 1363 41763 1539
rect 41987 1363 42021 1539
rect 42101 1363 42135 1539
rect 42359 1363 42393 1539
rect 42473 1363 42507 1539
rect 42731 1363 42765 1539
rect 42845 1363 42879 1539
rect 43103 1363 43137 1539
rect 43217 1363 43251 1539
rect 43475 1363 43509 1539
rect 43589 1363 43623 1539
rect 43847 1363 43881 1539
rect 43961 1363 43995 1539
rect 44219 1363 44253 1539
rect 44333 1363 44367 1539
rect 44591 1363 44625 1539
rect 44705 1363 44739 1539
rect 44963 1363 44997 1539
rect 45077 1363 45111 1539
rect 45335 1363 45369 1539
rect 45449 1363 45483 1539
rect 45707 1363 45741 1539
rect 45821 1363 45855 1539
rect 46079 1363 46113 1539
rect 46193 1363 46227 1539
rect 46451 1363 46485 1539
rect 46565 1363 46599 1539
rect 46823 1363 46857 1539
rect 46937 1363 46971 1539
rect 47195 1363 47229 1539
rect 47309 1363 47343 1539
rect 47567 1363 47601 1539
rect 47681 1363 47715 1539
rect 47939 1363 47973 1539
rect 48053 1363 48087 1539
rect 48311 1363 48345 1539
rect 39497 945 39531 1121
rect 39755 945 39789 1121
rect 39869 945 39903 1121
rect 40127 945 40161 1121
rect 40241 945 40275 1121
rect 40499 945 40533 1121
rect 40613 945 40647 1121
rect 40871 945 40905 1121
rect 40985 945 41019 1121
rect 41243 945 41277 1121
rect 41357 945 41391 1121
rect 41615 945 41649 1121
rect 41729 945 41763 1121
rect 41987 945 42021 1121
rect 42101 945 42135 1121
rect 42359 945 42393 1121
rect 42473 945 42507 1121
rect 42731 945 42765 1121
rect 42845 945 42879 1121
rect 43103 945 43137 1121
rect 43217 945 43251 1121
rect 43475 945 43509 1121
rect 43589 945 43623 1121
rect 43847 945 43881 1121
rect 43961 945 43995 1121
rect 44219 945 44253 1121
rect 44333 945 44367 1121
rect 44591 945 44625 1121
rect 44705 945 44739 1121
rect 44963 945 44997 1121
rect 45077 945 45111 1121
rect 45335 945 45369 1121
rect 45449 945 45483 1121
rect 45707 945 45741 1121
rect 45821 945 45855 1121
rect 46079 945 46113 1121
rect 46193 945 46227 1121
rect 46451 945 46485 1121
rect 46565 945 46599 1121
rect 46823 945 46857 1121
rect 46937 945 46971 1121
rect 47195 945 47229 1121
rect 47309 945 47343 1121
rect 47567 945 47601 1121
rect 47681 945 47715 1121
rect 47939 945 47973 1121
rect 48053 945 48087 1121
rect 48311 945 48345 1121
rect 39497 527 39531 703
rect 39755 527 39789 703
rect 39869 527 39903 703
rect 40127 527 40161 703
rect 40241 527 40275 703
rect 40499 527 40533 703
rect 40613 527 40647 703
rect 40871 527 40905 703
rect 40985 527 41019 703
rect 41243 527 41277 703
rect 41357 527 41391 703
rect 41615 527 41649 703
rect 41729 527 41763 703
rect 41987 527 42021 703
rect 42101 527 42135 703
rect 42359 527 42393 703
rect 42473 527 42507 703
rect 42731 527 42765 703
rect 42845 527 42879 703
rect 43103 527 43137 703
rect 43217 527 43251 703
rect 43475 527 43509 703
rect 43589 527 43623 703
rect 43847 527 43881 703
rect 43961 527 43995 703
rect 44219 527 44253 703
rect 44333 527 44367 703
rect 44591 527 44625 703
rect 44705 527 44739 703
rect 44963 527 44997 703
rect 45077 527 45111 703
rect 45335 527 45369 703
rect 45449 527 45483 703
rect 45707 527 45741 703
rect 45821 527 45855 703
rect 46079 527 46113 703
rect 46193 527 46227 703
rect 46451 527 46485 703
rect 46565 527 46599 703
rect 46823 527 46857 703
rect 46937 527 46971 703
rect 47195 527 47229 703
rect 47309 527 47343 703
rect 47567 527 47601 703
rect 47681 527 47715 703
rect 47939 527 47973 703
rect 48053 527 48087 703
rect 48311 527 48345 703
<< pdiffc >>
rect 38009 8654 38043 9030
rect 38267 8654 38301 9030
rect 38381 8654 38415 9030
rect 38639 8654 38673 9030
rect 38753 8654 38787 9030
rect 39011 8654 39045 9030
rect 39125 8654 39159 9030
rect 39383 8654 39417 9030
rect 39497 8654 39531 9030
rect 39755 8654 39789 9030
rect 39869 8654 39903 9030
rect 40127 8654 40161 9030
rect 40241 8654 40275 9030
rect 40499 8654 40533 9030
rect 40613 8654 40647 9030
rect 40871 8654 40905 9030
rect 40985 8654 41019 9030
rect 41243 8654 41277 9030
rect 41357 8654 41391 9030
rect 41615 8654 41649 9030
rect 41729 8654 41763 9030
rect 41987 8654 42021 9030
rect 42101 8654 42135 9030
rect 42359 8654 42393 9030
rect 42473 8654 42507 9030
rect 42731 8654 42765 9030
rect 42845 8654 42879 9030
rect 43103 8654 43137 9030
rect 43217 8654 43251 9030
rect 43475 8654 43509 9030
rect 43589 8654 43623 9030
rect 43847 8654 43881 9030
rect 43961 8654 43995 9030
rect 44219 8654 44253 9030
rect 44333 8654 44367 9030
rect 44591 8654 44625 9030
rect 44705 8654 44739 9030
rect 44963 8654 44997 9030
rect 45077 8654 45111 9030
rect 45335 8654 45369 9030
rect 45449 8654 45483 9030
rect 45707 8654 45741 9030
rect 45821 8654 45855 9030
rect 46079 8654 46113 9030
rect 46193 8654 46227 9030
rect 46451 8654 46485 9030
rect 46565 8654 46599 9030
rect 46823 8654 46857 9030
rect 46937 8654 46971 9030
rect 47195 8654 47229 9030
rect 47309 8654 47343 9030
rect 47567 8654 47601 9030
rect 47681 8654 47715 9030
rect 47939 8654 47973 9030
rect 48053 8654 48087 9030
rect 48311 8654 48345 9030
rect 48425 8654 48459 9030
rect 48683 8654 48717 9030
rect 48797 8654 48831 9030
rect 49055 8654 49089 9030
rect 49169 8654 49203 9030
rect 49427 8654 49461 9030
rect 49541 8654 49575 9030
rect 49799 8654 49833 9030
rect 38009 8018 38043 8394
rect 38267 8018 38301 8394
rect 38381 8018 38415 8394
rect 38639 8018 38673 8394
rect 38753 8018 38787 8394
rect 39011 8018 39045 8394
rect 39125 8018 39159 8394
rect 39383 8018 39417 8394
rect 39497 8018 39531 8394
rect 39755 8018 39789 8394
rect 39869 8018 39903 8394
rect 40127 8018 40161 8394
rect 40241 8018 40275 8394
rect 40499 8018 40533 8394
rect 40613 8018 40647 8394
rect 40871 8018 40905 8394
rect 40985 8018 41019 8394
rect 41243 8018 41277 8394
rect 41357 8018 41391 8394
rect 41615 8018 41649 8394
rect 41729 8018 41763 8394
rect 41987 8018 42021 8394
rect 42101 8018 42135 8394
rect 42359 8018 42393 8394
rect 42473 8018 42507 8394
rect 42731 8018 42765 8394
rect 42845 8018 42879 8394
rect 43103 8018 43137 8394
rect 43217 8018 43251 8394
rect 43475 8018 43509 8394
rect 43589 8018 43623 8394
rect 43847 8018 43881 8394
rect 43961 8018 43995 8394
rect 44219 8018 44253 8394
rect 44333 8018 44367 8394
rect 44591 8018 44625 8394
rect 44705 8018 44739 8394
rect 44963 8018 44997 8394
rect 45077 8018 45111 8394
rect 45335 8018 45369 8394
rect 45449 8018 45483 8394
rect 45707 8018 45741 8394
rect 45821 8018 45855 8394
rect 46079 8018 46113 8394
rect 46193 8018 46227 8394
rect 46451 8018 46485 8394
rect 46565 8018 46599 8394
rect 46823 8018 46857 8394
rect 46937 8018 46971 8394
rect 47195 8018 47229 8394
rect 47309 8018 47343 8394
rect 47567 8018 47601 8394
rect 47681 8018 47715 8394
rect 47939 8018 47973 8394
rect 48053 8018 48087 8394
rect 48311 8018 48345 8394
rect 48425 8018 48459 8394
rect 48683 8018 48717 8394
rect 48797 8018 48831 8394
rect 49055 8018 49089 8394
rect 49169 8018 49203 8394
rect 49427 8018 49461 8394
rect 49541 8018 49575 8394
rect 49799 8018 49833 8394
rect 38009 7382 38043 7758
rect 38267 7382 38301 7758
rect 38381 7382 38415 7758
rect 38639 7382 38673 7758
rect 38753 7382 38787 7758
rect 39011 7382 39045 7758
rect 39125 7382 39159 7758
rect 39383 7382 39417 7758
rect 39497 7382 39531 7758
rect 39755 7382 39789 7758
rect 39869 7382 39903 7758
rect 40127 7382 40161 7758
rect 40241 7382 40275 7758
rect 40499 7382 40533 7758
rect 40613 7382 40647 7758
rect 40871 7382 40905 7758
rect 40985 7382 41019 7758
rect 41243 7382 41277 7758
rect 41357 7382 41391 7758
rect 41615 7382 41649 7758
rect 41729 7382 41763 7758
rect 41987 7382 42021 7758
rect 42101 7382 42135 7758
rect 42359 7382 42393 7758
rect 42473 7382 42507 7758
rect 42731 7382 42765 7758
rect 42845 7382 42879 7758
rect 43103 7382 43137 7758
rect 43217 7382 43251 7758
rect 43475 7382 43509 7758
rect 43589 7382 43623 7758
rect 43847 7382 43881 7758
rect 43961 7382 43995 7758
rect 44219 7382 44253 7758
rect 44333 7382 44367 7758
rect 44591 7382 44625 7758
rect 44705 7382 44739 7758
rect 44963 7382 44997 7758
rect 45077 7382 45111 7758
rect 45335 7382 45369 7758
rect 45449 7382 45483 7758
rect 45707 7382 45741 7758
rect 45821 7382 45855 7758
rect 46079 7382 46113 7758
rect 46193 7382 46227 7758
rect 46451 7382 46485 7758
rect 46565 7382 46599 7758
rect 46823 7382 46857 7758
rect 46937 7382 46971 7758
rect 47195 7382 47229 7758
rect 47309 7382 47343 7758
rect 47567 7382 47601 7758
rect 47681 7382 47715 7758
rect 47939 7382 47973 7758
rect 48053 7382 48087 7758
rect 48311 7382 48345 7758
rect 48425 7382 48459 7758
rect 48683 7382 48717 7758
rect 48797 7382 48831 7758
rect 49055 7382 49089 7758
rect 49169 7382 49203 7758
rect 49427 7382 49461 7758
rect 49541 7382 49575 7758
rect 49799 7382 49833 7758
rect 39497 5866 39531 6642
rect 39755 5866 39789 6642
rect 39869 5866 39903 6642
rect 40127 5866 40161 6642
rect 40241 5866 40275 6642
rect 40499 5866 40533 6642
rect 40613 5866 40647 6642
rect 40871 5866 40905 6642
rect 40985 5866 41019 6642
rect 41243 5866 41277 6642
rect 41357 5866 41391 6642
rect 41615 5866 41649 6642
rect 41729 5866 41763 6642
rect 41987 5866 42021 6642
rect 42101 5866 42135 6642
rect 42359 5866 42393 6642
rect 39497 4830 39531 5606
rect 39755 4830 39789 5606
rect 39869 4830 39903 5606
rect 40127 4830 40161 5606
rect 40241 4830 40275 5606
rect 40499 4830 40533 5606
rect 40613 4830 40647 5606
rect 40871 4830 40905 5606
rect 40985 4830 41019 5606
rect 41243 4830 41277 5606
rect 41357 4830 41391 5606
rect 41615 4830 41649 5606
rect 41729 4830 41763 5606
rect 41987 4830 42021 5606
rect 42101 4830 42135 5606
rect 42359 4830 42393 5606
rect 39497 3794 39531 4570
rect 39755 3794 39789 4570
rect 39869 3794 39903 4570
rect 40127 3794 40161 4570
rect 40241 3794 40275 4570
rect 40499 3794 40533 4570
rect 40613 3794 40647 4570
rect 40871 3794 40905 4570
rect 40985 3794 41019 4570
rect 41243 3794 41277 4570
rect 41357 3794 41391 4570
rect 41615 3794 41649 4570
rect 41729 3794 41763 4570
rect 41987 3794 42021 4570
rect 42101 3794 42135 4570
rect 42359 3794 42393 4570
rect 39497 2758 39531 3534
rect 39755 2758 39789 3534
rect 39869 2758 39903 3534
rect 40127 2758 40161 3534
rect 40241 2758 40275 3534
rect 40499 2758 40533 3534
rect 40613 2758 40647 3534
rect 40871 2758 40905 3534
rect 40985 2758 41019 3534
rect 41243 2758 41277 3534
rect 41357 2758 41391 3534
rect 41615 2758 41649 3534
rect 41729 2758 41763 3534
rect 41987 2758 42021 3534
rect 42101 2758 42135 3534
rect 42359 2758 42393 3534
<< psubdiff >>
rect 43009 4889 43105 4923
rect 43243 4889 43339 4923
rect 43009 4827 43043 4889
rect 43305 4827 43339 4889
rect 43009 3273 43043 3335
rect 43305 3273 43339 3335
rect 43009 3239 43105 3273
rect 43243 3239 43339 3273
rect 39383 2109 39479 2143
rect 48363 2109 48459 2143
rect 39383 2047 39417 2109
rect 48425 2047 48459 2109
rect 39383 375 39417 437
rect 48425 375 48459 437
rect 39383 341 39479 375
rect 48363 341 48459 375
<< nsubdiff >>
rect 37895 9191 37991 9225
rect 49851 9191 49947 9225
rect 37895 9129 37929 9191
rect 49913 9129 49947 9191
rect 37895 7221 37929 7283
rect 49913 7221 49947 7283
rect 37895 7187 37991 7221
rect 49851 7187 49947 7221
rect 39383 6803 39479 6837
rect 42411 6803 42507 6837
rect 39383 6741 39417 6803
rect 42473 6741 42507 6803
rect 39383 2597 39417 2659
rect 42473 2597 42507 2659
rect 39383 2563 39479 2597
rect 42411 2563 42507 2597
<< psubdiffcont >>
rect 43105 4889 43243 4923
rect 43009 3335 43043 4827
rect 43305 3335 43339 4827
rect 43105 3239 43243 3273
rect 39479 2109 48363 2143
rect 39383 437 39417 2047
rect 48425 437 48459 2047
rect 39479 341 48363 375
<< nsubdiffcont >>
rect 37991 9191 49851 9225
rect 37895 7283 37929 9129
rect 49913 7283 49947 9129
rect 37991 7187 49851 7221
rect 39479 6803 42411 6837
rect 39383 2659 39417 6741
rect 42473 2659 42507 6741
rect 39479 2563 42411 2597
<< poly >>
rect 38055 9123 38255 9139
rect 38055 9089 38071 9123
rect 38239 9089 38255 9123
rect 38055 9042 38255 9089
rect 38427 9123 38627 9139
rect 38427 9089 38443 9123
rect 38611 9089 38627 9123
rect 38427 9042 38627 9089
rect 38799 9123 38999 9139
rect 38799 9089 38815 9123
rect 38983 9089 38999 9123
rect 38799 9042 38999 9089
rect 39171 9123 39371 9139
rect 39171 9089 39187 9123
rect 39355 9089 39371 9123
rect 39171 9042 39371 9089
rect 39543 9123 39743 9139
rect 39543 9089 39559 9123
rect 39727 9089 39743 9123
rect 39543 9042 39743 9089
rect 39915 9123 40115 9139
rect 39915 9089 39931 9123
rect 40099 9089 40115 9123
rect 39915 9042 40115 9089
rect 40287 9123 40487 9139
rect 40287 9089 40303 9123
rect 40471 9089 40487 9123
rect 40287 9042 40487 9089
rect 40659 9123 40859 9139
rect 40659 9089 40675 9123
rect 40843 9089 40859 9123
rect 40659 9042 40859 9089
rect 41031 9123 41231 9139
rect 41031 9089 41047 9123
rect 41215 9089 41231 9123
rect 41031 9042 41231 9089
rect 41403 9123 41603 9139
rect 41403 9089 41419 9123
rect 41587 9089 41603 9123
rect 41403 9042 41603 9089
rect 41775 9123 41975 9139
rect 41775 9089 41791 9123
rect 41959 9089 41975 9123
rect 41775 9042 41975 9089
rect 42147 9123 42347 9139
rect 42147 9089 42163 9123
rect 42331 9089 42347 9123
rect 42147 9042 42347 9089
rect 42519 9123 42719 9139
rect 42519 9089 42535 9123
rect 42703 9089 42719 9123
rect 42519 9042 42719 9089
rect 42891 9123 43091 9139
rect 42891 9089 42907 9123
rect 43075 9089 43091 9123
rect 42891 9042 43091 9089
rect 43263 9123 43463 9139
rect 43263 9089 43279 9123
rect 43447 9089 43463 9123
rect 43263 9042 43463 9089
rect 43635 9123 43835 9139
rect 43635 9089 43651 9123
rect 43819 9089 43835 9123
rect 43635 9042 43835 9089
rect 44007 9123 44207 9139
rect 44007 9089 44023 9123
rect 44191 9089 44207 9123
rect 44007 9042 44207 9089
rect 44379 9123 44579 9139
rect 44379 9089 44395 9123
rect 44563 9089 44579 9123
rect 44379 9042 44579 9089
rect 44751 9123 44951 9139
rect 44751 9089 44767 9123
rect 44935 9089 44951 9123
rect 44751 9042 44951 9089
rect 45123 9123 45323 9139
rect 45123 9089 45139 9123
rect 45307 9089 45323 9123
rect 45123 9042 45323 9089
rect 45495 9123 45695 9139
rect 45495 9089 45511 9123
rect 45679 9089 45695 9123
rect 45495 9042 45695 9089
rect 45867 9123 46067 9139
rect 45867 9089 45883 9123
rect 46051 9089 46067 9123
rect 45867 9042 46067 9089
rect 46239 9123 46439 9139
rect 46239 9089 46255 9123
rect 46423 9089 46439 9123
rect 46239 9042 46439 9089
rect 46611 9123 46811 9139
rect 46611 9089 46627 9123
rect 46795 9089 46811 9123
rect 46611 9042 46811 9089
rect 46983 9123 47183 9139
rect 46983 9089 46999 9123
rect 47167 9089 47183 9123
rect 46983 9042 47183 9089
rect 47355 9123 47555 9139
rect 47355 9089 47371 9123
rect 47539 9089 47555 9123
rect 47355 9042 47555 9089
rect 47727 9123 47927 9139
rect 47727 9089 47743 9123
rect 47911 9089 47927 9123
rect 47727 9042 47927 9089
rect 48099 9123 48299 9139
rect 48099 9089 48115 9123
rect 48283 9089 48299 9123
rect 48099 9042 48299 9089
rect 48471 9123 48671 9139
rect 48471 9089 48487 9123
rect 48655 9089 48671 9123
rect 48471 9042 48671 9089
rect 48843 9123 49043 9139
rect 48843 9089 48859 9123
rect 49027 9089 49043 9123
rect 48843 9042 49043 9089
rect 49215 9123 49415 9139
rect 49215 9089 49231 9123
rect 49399 9089 49415 9123
rect 49215 9042 49415 9089
rect 49587 9123 49787 9139
rect 49587 9089 49603 9123
rect 49771 9089 49787 9123
rect 49587 9042 49787 9089
rect 38055 8595 38255 8642
rect 38055 8561 38071 8595
rect 38239 8561 38255 8595
rect 38055 8545 38255 8561
rect 38427 8595 38627 8642
rect 38427 8561 38443 8595
rect 38611 8561 38627 8595
rect 38427 8545 38627 8561
rect 38799 8595 38999 8642
rect 38799 8561 38815 8595
rect 38983 8561 38999 8595
rect 38799 8545 38999 8561
rect 39171 8595 39371 8642
rect 39171 8561 39187 8595
rect 39355 8561 39371 8595
rect 39171 8545 39371 8561
rect 39543 8595 39743 8642
rect 39543 8561 39559 8595
rect 39727 8561 39743 8595
rect 39543 8545 39743 8561
rect 39915 8595 40115 8642
rect 39915 8561 39931 8595
rect 40099 8561 40115 8595
rect 39915 8545 40115 8561
rect 40287 8595 40487 8642
rect 40287 8561 40303 8595
rect 40471 8561 40487 8595
rect 40287 8545 40487 8561
rect 40659 8595 40859 8642
rect 40659 8561 40675 8595
rect 40843 8561 40859 8595
rect 40659 8545 40859 8561
rect 41031 8595 41231 8642
rect 41031 8561 41047 8595
rect 41215 8561 41231 8595
rect 41031 8545 41231 8561
rect 41403 8595 41603 8642
rect 41403 8561 41419 8595
rect 41587 8561 41603 8595
rect 41403 8545 41603 8561
rect 41775 8595 41975 8642
rect 41775 8561 41791 8595
rect 41959 8561 41975 8595
rect 41775 8545 41975 8561
rect 42147 8595 42347 8642
rect 42147 8561 42163 8595
rect 42331 8561 42347 8595
rect 42147 8545 42347 8561
rect 42519 8595 42719 8642
rect 42519 8561 42535 8595
rect 42703 8561 42719 8595
rect 42519 8545 42719 8561
rect 42891 8595 43091 8642
rect 42891 8561 42907 8595
rect 43075 8561 43091 8595
rect 42891 8545 43091 8561
rect 43263 8595 43463 8642
rect 43263 8561 43279 8595
rect 43447 8561 43463 8595
rect 43263 8545 43463 8561
rect 43635 8595 43835 8642
rect 43635 8561 43651 8595
rect 43819 8561 43835 8595
rect 43635 8545 43835 8561
rect 44007 8595 44207 8642
rect 44007 8561 44023 8595
rect 44191 8561 44207 8595
rect 44007 8545 44207 8561
rect 44379 8595 44579 8642
rect 44379 8561 44395 8595
rect 44563 8561 44579 8595
rect 44379 8545 44579 8561
rect 44751 8595 44951 8642
rect 44751 8561 44767 8595
rect 44935 8561 44951 8595
rect 44751 8545 44951 8561
rect 45123 8595 45323 8642
rect 45123 8561 45139 8595
rect 45307 8561 45323 8595
rect 45123 8545 45323 8561
rect 45495 8595 45695 8642
rect 45495 8561 45511 8595
rect 45679 8561 45695 8595
rect 45495 8545 45695 8561
rect 45867 8595 46067 8642
rect 45867 8561 45883 8595
rect 46051 8561 46067 8595
rect 45867 8545 46067 8561
rect 46239 8595 46439 8642
rect 46239 8561 46255 8595
rect 46423 8561 46439 8595
rect 46239 8545 46439 8561
rect 46611 8595 46811 8642
rect 46611 8561 46627 8595
rect 46795 8561 46811 8595
rect 46611 8545 46811 8561
rect 46983 8595 47183 8642
rect 46983 8561 46999 8595
rect 47167 8561 47183 8595
rect 46983 8545 47183 8561
rect 47355 8595 47555 8642
rect 47355 8561 47371 8595
rect 47539 8561 47555 8595
rect 47355 8545 47555 8561
rect 47727 8595 47927 8642
rect 47727 8561 47743 8595
rect 47911 8561 47927 8595
rect 47727 8545 47927 8561
rect 48099 8595 48299 8642
rect 48099 8561 48115 8595
rect 48283 8561 48299 8595
rect 48099 8545 48299 8561
rect 48471 8595 48671 8642
rect 48471 8561 48487 8595
rect 48655 8561 48671 8595
rect 48471 8545 48671 8561
rect 48843 8595 49043 8642
rect 48843 8561 48859 8595
rect 49027 8561 49043 8595
rect 48843 8545 49043 8561
rect 49215 8595 49415 8642
rect 49215 8561 49231 8595
rect 49399 8561 49415 8595
rect 49215 8545 49415 8561
rect 49587 8595 49787 8642
rect 49587 8561 49603 8595
rect 49771 8561 49787 8595
rect 49587 8545 49787 8561
rect 38055 8487 38255 8503
rect 38055 8453 38071 8487
rect 38239 8453 38255 8487
rect 38055 8406 38255 8453
rect 38427 8487 38627 8503
rect 38427 8453 38443 8487
rect 38611 8453 38627 8487
rect 38427 8406 38627 8453
rect 38799 8487 38999 8503
rect 38799 8453 38815 8487
rect 38983 8453 38999 8487
rect 38799 8406 38999 8453
rect 39171 8487 39371 8503
rect 39171 8453 39187 8487
rect 39355 8453 39371 8487
rect 39171 8406 39371 8453
rect 39543 8487 39743 8503
rect 39543 8453 39559 8487
rect 39727 8453 39743 8487
rect 39543 8406 39743 8453
rect 39915 8487 40115 8503
rect 39915 8453 39931 8487
rect 40099 8453 40115 8487
rect 39915 8406 40115 8453
rect 40287 8487 40487 8503
rect 40287 8453 40303 8487
rect 40471 8453 40487 8487
rect 40287 8406 40487 8453
rect 40659 8487 40859 8503
rect 40659 8453 40675 8487
rect 40843 8453 40859 8487
rect 40659 8406 40859 8453
rect 41031 8487 41231 8503
rect 41031 8453 41047 8487
rect 41215 8453 41231 8487
rect 41031 8406 41231 8453
rect 41403 8487 41603 8503
rect 41403 8453 41419 8487
rect 41587 8453 41603 8487
rect 41403 8406 41603 8453
rect 41775 8487 41975 8503
rect 41775 8453 41791 8487
rect 41959 8453 41975 8487
rect 41775 8406 41975 8453
rect 42147 8487 42347 8503
rect 42147 8453 42163 8487
rect 42331 8453 42347 8487
rect 42147 8406 42347 8453
rect 42519 8487 42719 8503
rect 42519 8453 42535 8487
rect 42703 8453 42719 8487
rect 42519 8406 42719 8453
rect 42891 8487 43091 8503
rect 42891 8453 42907 8487
rect 43075 8453 43091 8487
rect 42891 8406 43091 8453
rect 43263 8487 43463 8503
rect 43263 8453 43279 8487
rect 43447 8453 43463 8487
rect 43263 8406 43463 8453
rect 43635 8487 43835 8503
rect 43635 8453 43651 8487
rect 43819 8453 43835 8487
rect 43635 8406 43835 8453
rect 44007 8487 44207 8503
rect 44007 8453 44023 8487
rect 44191 8453 44207 8487
rect 44007 8406 44207 8453
rect 44379 8487 44579 8503
rect 44379 8453 44395 8487
rect 44563 8453 44579 8487
rect 44379 8406 44579 8453
rect 44751 8487 44951 8503
rect 44751 8453 44767 8487
rect 44935 8453 44951 8487
rect 44751 8406 44951 8453
rect 45123 8487 45323 8503
rect 45123 8453 45139 8487
rect 45307 8453 45323 8487
rect 45123 8406 45323 8453
rect 45495 8487 45695 8503
rect 45495 8453 45511 8487
rect 45679 8453 45695 8487
rect 45495 8406 45695 8453
rect 45867 8487 46067 8503
rect 45867 8453 45883 8487
rect 46051 8453 46067 8487
rect 45867 8406 46067 8453
rect 46239 8487 46439 8503
rect 46239 8453 46255 8487
rect 46423 8453 46439 8487
rect 46239 8406 46439 8453
rect 46611 8487 46811 8503
rect 46611 8453 46627 8487
rect 46795 8453 46811 8487
rect 46611 8406 46811 8453
rect 46983 8487 47183 8503
rect 46983 8453 46999 8487
rect 47167 8453 47183 8487
rect 46983 8406 47183 8453
rect 47355 8487 47555 8503
rect 47355 8453 47371 8487
rect 47539 8453 47555 8487
rect 47355 8406 47555 8453
rect 47727 8487 47927 8503
rect 47727 8453 47743 8487
rect 47911 8453 47927 8487
rect 47727 8406 47927 8453
rect 48099 8487 48299 8503
rect 48099 8453 48115 8487
rect 48283 8453 48299 8487
rect 48099 8406 48299 8453
rect 48471 8487 48671 8503
rect 48471 8453 48487 8487
rect 48655 8453 48671 8487
rect 48471 8406 48671 8453
rect 48843 8487 49043 8503
rect 48843 8453 48859 8487
rect 49027 8453 49043 8487
rect 48843 8406 49043 8453
rect 49215 8487 49415 8503
rect 49215 8453 49231 8487
rect 49399 8453 49415 8487
rect 49215 8406 49415 8453
rect 49587 8487 49787 8503
rect 49587 8453 49603 8487
rect 49771 8453 49787 8487
rect 49587 8406 49787 8453
rect 38055 7959 38255 8006
rect 38055 7925 38071 7959
rect 38239 7925 38255 7959
rect 38055 7909 38255 7925
rect 38427 7959 38627 8006
rect 38427 7925 38443 7959
rect 38611 7925 38627 7959
rect 38427 7909 38627 7925
rect 38799 7959 38999 8006
rect 38799 7925 38815 7959
rect 38983 7925 38999 7959
rect 38799 7909 38999 7925
rect 39171 7959 39371 8006
rect 39171 7925 39187 7959
rect 39355 7925 39371 7959
rect 39171 7909 39371 7925
rect 39543 7959 39743 8006
rect 39543 7925 39559 7959
rect 39727 7925 39743 7959
rect 39543 7909 39743 7925
rect 39915 7959 40115 8006
rect 39915 7925 39931 7959
rect 40099 7925 40115 7959
rect 39915 7909 40115 7925
rect 40287 7959 40487 8006
rect 40287 7925 40303 7959
rect 40471 7925 40487 7959
rect 40287 7909 40487 7925
rect 40659 7959 40859 8006
rect 40659 7925 40675 7959
rect 40843 7925 40859 7959
rect 40659 7909 40859 7925
rect 41031 7959 41231 8006
rect 41031 7925 41047 7959
rect 41215 7925 41231 7959
rect 41031 7909 41231 7925
rect 41403 7959 41603 8006
rect 41403 7925 41419 7959
rect 41587 7925 41603 7959
rect 41403 7909 41603 7925
rect 41775 7959 41975 8006
rect 41775 7925 41791 7959
rect 41959 7925 41975 7959
rect 41775 7909 41975 7925
rect 42147 7959 42347 8006
rect 42147 7925 42163 7959
rect 42331 7925 42347 7959
rect 42147 7909 42347 7925
rect 42519 7959 42719 8006
rect 42519 7925 42535 7959
rect 42703 7925 42719 7959
rect 42519 7909 42719 7925
rect 42891 7959 43091 8006
rect 42891 7925 42907 7959
rect 43075 7925 43091 7959
rect 42891 7909 43091 7925
rect 43263 7959 43463 8006
rect 43263 7925 43279 7959
rect 43447 7925 43463 7959
rect 43263 7909 43463 7925
rect 43635 7959 43835 8006
rect 43635 7925 43651 7959
rect 43819 7925 43835 7959
rect 43635 7909 43835 7925
rect 44007 7959 44207 8006
rect 44007 7925 44023 7959
rect 44191 7925 44207 7959
rect 44007 7909 44207 7925
rect 44379 7959 44579 8006
rect 44379 7925 44395 7959
rect 44563 7925 44579 7959
rect 44379 7909 44579 7925
rect 44751 7959 44951 8006
rect 44751 7925 44767 7959
rect 44935 7925 44951 7959
rect 44751 7909 44951 7925
rect 45123 7959 45323 8006
rect 45123 7925 45139 7959
rect 45307 7925 45323 7959
rect 45123 7909 45323 7925
rect 45495 7959 45695 8006
rect 45495 7925 45511 7959
rect 45679 7925 45695 7959
rect 45495 7909 45695 7925
rect 45867 7959 46067 8006
rect 45867 7925 45883 7959
rect 46051 7925 46067 7959
rect 45867 7909 46067 7925
rect 46239 7959 46439 8006
rect 46239 7925 46255 7959
rect 46423 7925 46439 7959
rect 46239 7909 46439 7925
rect 46611 7959 46811 8006
rect 46611 7925 46627 7959
rect 46795 7925 46811 7959
rect 46611 7909 46811 7925
rect 46983 7959 47183 8006
rect 46983 7925 46999 7959
rect 47167 7925 47183 7959
rect 46983 7909 47183 7925
rect 47355 7959 47555 8006
rect 47355 7925 47371 7959
rect 47539 7925 47555 7959
rect 47355 7909 47555 7925
rect 47727 7959 47927 8006
rect 47727 7925 47743 7959
rect 47911 7925 47927 7959
rect 47727 7909 47927 7925
rect 48099 7959 48299 8006
rect 48099 7925 48115 7959
rect 48283 7925 48299 7959
rect 48099 7909 48299 7925
rect 48471 7959 48671 8006
rect 48471 7925 48487 7959
rect 48655 7925 48671 7959
rect 48471 7909 48671 7925
rect 48843 7959 49043 8006
rect 48843 7925 48859 7959
rect 49027 7925 49043 7959
rect 48843 7909 49043 7925
rect 49215 7959 49415 8006
rect 49215 7925 49231 7959
rect 49399 7925 49415 7959
rect 49215 7909 49415 7925
rect 49587 7959 49787 8006
rect 49587 7925 49603 7959
rect 49771 7925 49787 7959
rect 49587 7909 49787 7925
rect 38055 7851 38255 7867
rect 38055 7817 38071 7851
rect 38239 7817 38255 7851
rect 38055 7770 38255 7817
rect 38427 7851 38627 7867
rect 38427 7817 38443 7851
rect 38611 7817 38627 7851
rect 38427 7770 38627 7817
rect 38799 7851 38999 7867
rect 38799 7817 38815 7851
rect 38983 7817 38999 7851
rect 38799 7770 38999 7817
rect 39171 7851 39371 7867
rect 39171 7817 39187 7851
rect 39355 7817 39371 7851
rect 39171 7770 39371 7817
rect 39543 7851 39743 7867
rect 39543 7817 39559 7851
rect 39727 7817 39743 7851
rect 39543 7770 39743 7817
rect 39915 7851 40115 7867
rect 39915 7817 39931 7851
rect 40099 7817 40115 7851
rect 39915 7770 40115 7817
rect 40287 7851 40487 7867
rect 40287 7817 40303 7851
rect 40471 7817 40487 7851
rect 40287 7770 40487 7817
rect 40659 7851 40859 7867
rect 40659 7817 40675 7851
rect 40843 7817 40859 7851
rect 40659 7770 40859 7817
rect 41031 7851 41231 7867
rect 41031 7817 41047 7851
rect 41215 7817 41231 7851
rect 41031 7770 41231 7817
rect 41403 7851 41603 7867
rect 41403 7817 41419 7851
rect 41587 7817 41603 7851
rect 41403 7770 41603 7817
rect 41775 7851 41975 7867
rect 41775 7817 41791 7851
rect 41959 7817 41975 7851
rect 41775 7770 41975 7817
rect 42147 7851 42347 7867
rect 42147 7817 42163 7851
rect 42331 7817 42347 7851
rect 42147 7770 42347 7817
rect 42519 7851 42719 7867
rect 42519 7817 42535 7851
rect 42703 7817 42719 7851
rect 42519 7770 42719 7817
rect 42891 7851 43091 7867
rect 42891 7817 42907 7851
rect 43075 7817 43091 7851
rect 42891 7770 43091 7817
rect 43263 7851 43463 7867
rect 43263 7817 43279 7851
rect 43447 7817 43463 7851
rect 43263 7770 43463 7817
rect 43635 7851 43835 7867
rect 43635 7817 43651 7851
rect 43819 7817 43835 7851
rect 43635 7770 43835 7817
rect 44007 7851 44207 7867
rect 44007 7817 44023 7851
rect 44191 7817 44207 7851
rect 44007 7770 44207 7817
rect 44379 7851 44579 7867
rect 44379 7817 44395 7851
rect 44563 7817 44579 7851
rect 44379 7770 44579 7817
rect 44751 7851 44951 7867
rect 44751 7817 44767 7851
rect 44935 7817 44951 7851
rect 44751 7770 44951 7817
rect 45123 7851 45323 7867
rect 45123 7817 45139 7851
rect 45307 7817 45323 7851
rect 45123 7770 45323 7817
rect 45495 7851 45695 7867
rect 45495 7817 45511 7851
rect 45679 7817 45695 7851
rect 45495 7770 45695 7817
rect 45867 7851 46067 7867
rect 45867 7817 45883 7851
rect 46051 7817 46067 7851
rect 45867 7770 46067 7817
rect 46239 7851 46439 7867
rect 46239 7817 46255 7851
rect 46423 7817 46439 7851
rect 46239 7770 46439 7817
rect 46611 7851 46811 7867
rect 46611 7817 46627 7851
rect 46795 7817 46811 7851
rect 46611 7770 46811 7817
rect 46983 7851 47183 7867
rect 46983 7817 46999 7851
rect 47167 7817 47183 7851
rect 46983 7770 47183 7817
rect 47355 7851 47555 7867
rect 47355 7817 47371 7851
rect 47539 7817 47555 7851
rect 47355 7770 47555 7817
rect 47727 7851 47927 7867
rect 47727 7817 47743 7851
rect 47911 7817 47927 7851
rect 47727 7770 47927 7817
rect 48099 7851 48299 7867
rect 48099 7817 48115 7851
rect 48283 7817 48299 7851
rect 48099 7770 48299 7817
rect 48471 7851 48671 7867
rect 48471 7817 48487 7851
rect 48655 7817 48671 7851
rect 48471 7770 48671 7817
rect 48843 7851 49043 7867
rect 48843 7817 48859 7851
rect 49027 7817 49043 7851
rect 48843 7770 49043 7817
rect 49215 7851 49415 7867
rect 49215 7817 49231 7851
rect 49399 7817 49415 7851
rect 49215 7770 49415 7817
rect 49587 7851 49787 7867
rect 49587 7817 49603 7851
rect 49771 7817 49787 7851
rect 49587 7770 49787 7817
rect 38055 7323 38255 7370
rect 38055 7289 38071 7323
rect 38239 7289 38255 7323
rect 38055 7273 38255 7289
rect 38427 7323 38627 7370
rect 38427 7289 38443 7323
rect 38611 7289 38627 7323
rect 38427 7273 38627 7289
rect 38799 7323 38999 7370
rect 38799 7289 38815 7323
rect 38983 7289 38999 7323
rect 38799 7273 38999 7289
rect 39171 7323 39371 7370
rect 39171 7289 39187 7323
rect 39355 7289 39371 7323
rect 39171 7273 39371 7289
rect 39543 7323 39743 7370
rect 39543 7289 39559 7323
rect 39727 7289 39743 7323
rect 39543 7273 39743 7289
rect 39915 7323 40115 7370
rect 39915 7289 39931 7323
rect 40099 7289 40115 7323
rect 39915 7273 40115 7289
rect 40287 7323 40487 7370
rect 40287 7289 40303 7323
rect 40471 7289 40487 7323
rect 40287 7273 40487 7289
rect 40659 7323 40859 7370
rect 40659 7289 40675 7323
rect 40843 7289 40859 7323
rect 40659 7273 40859 7289
rect 41031 7323 41231 7370
rect 41031 7289 41047 7323
rect 41215 7289 41231 7323
rect 41031 7273 41231 7289
rect 41403 7323 41603 7370
rect 41403 7289 41419 7323
rect 41587 7289 41603 7323
rect 41403 7273 41603 7289
rect 41775 7323 41975 7370
rect 41775 7289 41791 7323
rect 41959 7289 41975 7323
rect 41775 7273 41975 7289
rect 42147 7323 42347 7370
rect 42147 7289 42163 7323
rect 42331 7289 42347 7323
rect 42147 7273 42347 7289
rect 42519 7323 42719 7370
rect 42519 7289 42535 7323
rect 42703 7289 42719 7323
rect 42519 7273 42719 7289
rect 42891 7323 43091 7370
rect 42891 7289 42907 7323
rect 43075 7289 43091 7323
rect 42891 7273 43091 7289
rect 43263 7323 43463 7370
rect 43263 7289 43279 7323
rect 43447 7289 43463 7323
rect 43263 7273 43463 7289
rect 43635 7323 43835 7370
rect 43635 7289 43651 7323
rect 43819 7289 43835 7323
rect 43635 7273 43835 7289
rect 44007 7323 44207 7370
rect 44007 7289 44023 7323
rect 44191 7289 44207 7323
rect 44007 7273 44207 7289
rect 44379 7323 44579 7370
rect 44379 7289 44395 7323
rect 44563 7289 44579 7323
rect 44379 7273 44579 7289
rect 44751 7323 44951 7370
rect 44751 7289 44767 7323
rect 44935 7289 44951 7323
rect 44751 7273 44951 7289
rect 45123 7323 45323 7370
rect 45123 7289 45139 7323
rect 45307 7289 45323 7323
rect 45123 7273 45323 7289
rect 45495 7323 45695 7370
rect 45495 7289 45511 7323
rect 45679 7289 45695 7323
rect 45495 7273 45695 7289
rect 45867 7323 46067 7370
rect 45867 7289 45883 7323
rect 46051 7289 46067 7323
rect 45867 7273 46067 7289
rect 46239 7323 46439 7370
rect 46239 7289 46255 7323
rect 46423 7289 46439 7323
rect 46239 7273 46439 7289
rect 46611 7323 46811 7370
rect 46611 7289 46627 7323
rect 46795 7289 46811 7323
rect 46611 7273 46811 7289
rect 46983 7323 47183 7370
rect 46983 7289 46999 7323
rect 47167 7289 47183 7323
rect 46983 7273 47183 7289
rect 47355 7323 47555 7370
rect 47355 7289 47371 7323
rect 47539 7289 47555 7323
rect 47355 7273 47555 7289
rect 47727 7323 47927 7370
rect 47727 7289 47743 7323
rect 47911 7289 47927 7323
rect 47727 7273 47927 7289
rect 48099 7323 48299 7370
rect 48099 7289 48115 7323
rect 48283 7289 48299 7323
rect 48099 7273 48299 7289
rect 48471 7323 48671 7370
rect 48471 7289 48487 7323
rect 48655 7289 48671 7323
rect 48471 7273 48671 7289
rect 48843 7323 49043 7370
rect 48843 7289 48859 7323
rect 49027 7289 49043 7323
rect 48843 7273 49043 7289
rect 49215 7323 49415 7370
rect 49215 7289 49231 7323
rect 49399 7289 49415 7323
rect 49215 7273 49415 7289
rect 49587 7323 49787 7370
rect 49587 7289 49603 7323
rect 49771 7289 49787 7323
rect 49587 7273 49787 7289
rect 39543 6735 39743 6751
rect 39543 6701 39559 6735
rect 39727 6701 39743 6735
rect 39543 6654 39743 6701
rect 39915 6735 40115 6751
rect 39915 6701 39931 6735
rect 40099 6701 40115 6735
rect 39915 6654 40115 6701
rect 40287 6735 40487 6751
rect 40287 6701 40303 6735
rect 40471 6701 40487 6735
rect 40287 6654 40487 6701
rect 40659 6735 40859 6751
rect 40659 6701 40675 6735
rect 40843 6701 40859 6735
rect 40659 6654 40859 6701
rect 41031 6735 41231 6751
rect 41031 6701 41047 6735
rect 41215 6701 41231 6735
rect 41031 6654 41231 6701
rect 41403 6735 41603 6751
rect 41403 6701 41419 6735
rect 41587 6701 41603 6735
rect 41403 6654 41603 6701
rect 41775 6735 41975 6751
rect 41775 6701 41791 6735
rect 41959 6701 41975 6735
rect 41775 6654 41975 6701
rect 42147 6735 42347 6751
rect 42147 6701 42163 6735
rect 42331 6701 42347 6735
rect 42147 6654 42347 6701
rect 39543 5807 39743 5854
rect 39543 5773 39559 5807
rect 39727 5773 39743 5807
rect 39543 5757 39743 5773
rect 39915 5807 40115 5854
rect 39915 5773 39931 5807
rect 40099 5773 40115 5807
rect 39915 5757 40115 5773
rect 40287 5807 40487 5854
rect 40287 5773 40303 5807
rect 40471 5773 40487 5807
rect 40287 5757 40487 5773
rect 40659 5807 40859 5854
rect 40659 5773 40675 5807
rect 40843 5773 40859 5807
rect 40659 5757 40859 5773
rect 41031 5807 41231 5854
rect 41031 5773 41047 5807
rect 41215 5773 41231 5807
rect 41031 5757 41231 5773
rect 41403 5807 41603 5854
rect 41403 5773 41419 5807
rect 41587 5773 41603 5807
rect 41403 5757 41603 5773
rect 41775 5807 41975 5854
rect 41775 5773 41791 5807
rect 41959 5773 41975 5807
rect 41775 5757 41975 5773
rect 42147 5807 42347 5854
rect 42147 5773 42163 5807
rect 42331 5773 42347 5807
rect 42147 5757 42347 5773
rect 39543 5699 39743 5715
rect 39543 5665 39559 5699
rect 39727 5665 39743 5699
rect 39543 5618 39743 5665
rect 39915 5699 40115 5715
rect 39915 5665 39931 5699
rect 40099 5665 40115 5699
rect 39915 5618 40115 5665
rect 40287 5699 40487 5715
rect 40287 5665 40303 5699
rect 40471 5665 40487 5699
rect 40287 5618 40487 5665
rect 40659 5699 40859 5715
rect 40659 5665 40675 5699
rect 40843 5665 40859 5699
rect 40659 5618 40859 5665
rect 41031 5699 41231 5715
rect 41031 5665 41047 5699
rect 41215 5665 41231 5699
rect 41031 5618 41231 5665
rect 41403 5699 41603 5715
rect 41403 5665 41419 5699
rect 41587 5665 41603 5699
rect 41403 5618 41603 5665
rect 41775 5699 41975 5715
rect 41775 5665 41791 5699
rect 41959 5665 41975 5699
rect 41775 5618 41975 5665
rect 42147 5699 42347 5715
rect 42147 5665 42163 5699
rect 42331 5665 42347 5699
rect 42147 5618 42347 5665
rect 39543 4771 39743 4818
rect 39543 4737 39559 4771
rect 39727 4737 39743 4771
rect 39543 4721 39743 4737
rect 39915 4771 40115 4818
rect 39915 4737 39931 4771
rect 40099 4737 40115 4771
rect 39915 4721 40115 4737
rect 40287 4771 40487 4818
rect 40287 4737 40303 4771
rect 40471 4737 40487 4771
rect 40287 4721 40487 4737
rect 40659 4771 40859 4818
rect 40659 4737 40675 4771
rect 40843 4737 40859 4771
rect 40659 4721 40859 4737
rect 41031 4771 41231 4818
rect 41031 4737 41047 4771
rect 41215 4737 41231 4771
rect 41031 4721 41231 4737
rect 41403 4771 41603 4818
rect 41403 4737 41419 4771
rect 41587 4737 41603 4771
rect 41403 4721 41603 4737
rect 41775 4771 41975 4818
rect 41775 4737 41791 4771
rect 41959 4737 41975 4771
rect 41775 4721 41975 4737
rect 42147 4771 42347 4818
rect 42147 4737 42163 4771
rect 42331 4737 42347 4771
rect 42147 4721 42347 4737
rect 39543 4663 39743 4679
rect 39543 4629 39559 4663
rect 39727 4629 39743 4663
rect 39543 4582 39743 4629
rect 39915 4663 40115 4679
rect 39915 4629 39931 4663
rect 40099 4629 40115 4663
rect 39915 4582 40115 4629
rect 40287 4663 40487 4679
rect 40287 4629 40303 4663
rect 40471 4629 40487 4663
rect 40287 4582 40487 4629
rect 40659 4663 40859 4679
rect 40659 4629 40675 4663
rect 40843 4629 40859 4663
rect 40659 4582 40859 4629
rect 41031 4663 41231 4679
rect 41031 4629 41047 4663
rect 41215 4629 41231 4663
rect 41031 4582 41231 4629
rect 41403 4663 41603 4679
rect 41403 4629 41419 4663
rect 41587 4629 41603 4663
rect 41403 4582 41603 4629
rect 41775 4663 41975 4679
rect 41775 4629 41791 4663
rect 41959 4629 41975 4663
rect 41775 4582 41975 4629
rect 42147 4663 42347 4679
rect 42147 4629 42163 4663
rect 42331 4629 42347 4663
rect 42147 4582 42347 4629
rect 39543 3735 39743 3782
rect 39543 3701 39559 3735
rect 39727 3701 39743 3735
rect 39543 3685 39743 3701
rect 39915 3735 40115 3782
rect 39915 3701 39931 3735
rect 40099 3701 40115 3735
rect 39915 3685 40115 3701
rect 40287 3735 40487 3782
rect 40287 3701 40303 3735
rect 40471 3701 40487 3735
rect 40287 3685 40487 3701
rect 40659 3735 40859 3782
rect 40659 3701 40675 3735
rect 40843 3701 40859 3735
rect 40659 3685 40859 3701
rect 41031 3735 41231 3782
rect 41031 3701 41047 3735
rect 41215 3701 41231 3735
rect 41031 3685 41231 3701
rect 41403 3735 41603 3782
rect 41403 3701 41419 3735
rect 41587 3701 41603 3735
rect 41403 3685 41603 3701
rect 41775 3735 41975 3782
rect 41775 3701 41791 3735
rect 41959 3701 41975 3735
rect 41775 3685 41975 3701
rect 42147 3735 42347 3782
rect 42147 3701 42163 3735
rect 42331 3701 42347 3735
rect 42147 3685 42347 3701
rect 39543 3627 39743 3643
rect 39543 3593 39559 3627
rect 39727 3593 39743 3627
rect 39543 3546 39743 3593
rect 39915 3627 40115 3643
rect 39915 3593 39931 3627
rect 40099 3593 40115 3627
rect 39915 3546 40115 3593
rect 40287 3627 40487 3643
rect 40287 3593 40303 3627
rect 40471 3593 40487 3627
rect 40287 3546 40487 3593
rect 40659 3627 40859 3643
rect 40659 3593 40675 3627
rect 40843 3593 40859 3627
rect 40659 3546 40859 3593
rect 41031 3627 41231 3643
rect 41031 3593 41047 3627
rect 41215 3593 41231 3627
rect 41031 3546 41231 3593
rect 41403 3627 41603 3643
rect 41403 3593 41419 3627
rect 41587 3593 41603 3627
rect 41403 3546 41603 3593
rect 41775 3627 41975 3643
rect 41775 3593 41791 3627
rect 41959 3593 41975 3627
rect 41775 3546 41975 3593
rect 42147 3627 42347 3643
rect 42147 3593 42163 3627
rect 42331 3593 42347 3627
rect 42147 3546 42347 3593
rect 39543 2699 39743 2746
rect 39543 2665 39559 2699
rect 39727 2665 39743 2699
rect 39543 2649 39743 2665
rect 39915 2699 40115 2746
rect 39915 2665 39931 2699
rect 40099 2665 40115 2699
rect 39915 2649 40115 2665
rect 40287 2699 40487 2746
rect 40287 2665 40303 2699
rect 40471 2665 40487 2699
rect 40287 2649 40487 2665
rect 40659 2699 40859 2746
rect 40659 2665 40675 2699
rect 40843 2665 40859 2699
rect 40659 2649 40859 2665
rect 41031 2699 41231 2746
rect 41031 2665 41047 2699
rect 41215 2665 41231 2699
rect 41031 2649 41231 2665
rect 41403 2699 41603 2746
rect 41403 2665 41419 2699
rect 41587 2665 41603 2699
rect 41403 2649 41603 2665
rect 41775 2699 41975 2746
rect 41775 2665 41791 2699
rect 41959 2665 41975 2699
rect 41775 2649 41975 2665
rect 42147 2699 42347 2746
rect 42147 2665 42163 2699
rect 42331 2665 42347 2699
rect 42147 2649 42347 2665
rect 39543 2041 39743 2057
rect 39543 2007 39559 2041
rect 39727 2007 39743 2041
rect 39543 1969 39743 2007
rect 39915 2041 40115 2057
rect 39915 2007 39931 2041
rect 40099 2007 40115 2041
rect 39915 1969 40115 2007
rect 40287 2041 40487 2057
rect 40287 2007 40303 2041
rect 40471 2007 40487 2041
rect 40287 1969 40487 2007
rect 40659 2041 40859 2057
rect 40659 2007 40675 2041
rect 40843 2007 40859 2041
rect 40659 1969 40859 2007
rect 41031 2041 41231 2057
rect 41031 2007 41047 2041
rect 41215 2007 41231 2041
rect 41031 1969 41231 2007
rect 41403 2041 41603 2057
rect 41403 2007 41419 2041
rect 41587 2007 41603 2041
rect 41403 1969 41603 2007
rect 41775 2041 41975 2057
rect 41775 2007 41791 2041
rect 41959 2007 41975 2041
rect 41775 1969 41975 2007
rect 42147 2041 42347 2057
rect 42147 2007 42163 2041
rect 42331 2007 42347 2041
rect 42147 1969 42347 2007
rect 42519 2041 42719 2057
rect 42519 2007 42535 2041
rect 42703 2007 42719 2041
rect 42519 1969 42719 2007
rect 42891 2041 43091 2057
rect 42891 2007 42907 2041
rect 43075 2007 43091 2041
rect 42891 1969 43091 2007
rect 43263 2041 43463 2057
rect 43263 2007 43279 2041
rect 43447 2007 43463 2041
rect 43263 1969 43463 2007
rect 43635 2041 43835 2057
rect 43635 2007 43651 2041
rect 43819 2007 43835 2041
rect 43635 1969 43835 2007
rect 44007 2041 44207 2057
rect 44007 2007 44023 2041
rect 44191 2007 44207 2041
rect 44007 1969 44207 2007
rect 44379 2041 44579 2057
rect 44379 2007 44395 2041
rect 44563 2007 44579 2041
rect 44379 1969 44579 2007
rect 44751 2041 44951 2057
rect 44751 2007 44767 2041
rect 44935 2007 44951 2041
rect 44751 1969 44951 2007
rect 45123 2041 45323 2057
rect 45123 2007 45139 2041
rect 45307 2007 45323 2041
rect 45123 1969 45323 2007
rect 45495 2041 45695 2057
rect 45495 2007 45511 2041
rect 45679 2007 45695 2041
rect 45495 1969 45695 2007
rect 45867 2041 46067 2057
rect 45867 2007 45883 2041
rect 46051 2007 46067 2041
rect 45867 1969 46067 2007
rect 46239 2041 46439 2057
rect 46239 2007 46255 2041
rect 46423 2007 46439 2041
rect 46239 1969 46439 2007
rect 46611 2041 46811 2057
rect 46611 2007 46627 2041
rect 46795 2007 46811 2041
rect 46611 1969 46811 2007
rect 46983 2041 47183 2057
rect 46983 2007 46999 2041
rect 47167 2007 47183 2041
rect 46983 1969 47183 2007
rect 47355 2041 47555 2057
rect 47355 2007 47371 2041
rect 47539 2007 47555 2041
rect 47355 1969 47555 2007
rect 47727 2041 47927 2057
rect 47727 2007 47743 2041
rect 47911 2007 47927 2041
rect 47727 1969 47927 2007
rect 48099 2041 48299 2057
rect 48099 2007 48115 2041
rect 48283 2007 48299 2041
rect 48099 1969 48299 2007
rect 39543 1731 39743 1769
rect 39543 1697 39559 1731
rect 39727 1697 39743 1731
rect 39543 1681 39743 1697
rect 39915 1731 40115 1769
rect 39915 1697 39931 1731
rect 40099 1697 40115 1731
rect 39915 1681 40115 1697
rect 40287 1731 40487 1769
rect 40287 1697 40303 1731
rect 40471 1697 40487 1731
rect 40287 1681 40487 1697
rect 40659 1731 40859 1769
rect 40659 1697 40675 1731
rect 40843 1697 40859 1731
rect 40659 1681 40859 1697
rect 41031 1731 41231 1769
rect 41031 1697 41047 1731
rect 41215 1697 41231 1731
rect 41031 1681 41231 1697
rect 41403 1731 41603 1769
rect 41403 1697 41419 1731
rect 41587 1697 41603 1731
rect 41403 1681 41603 1697
rect 41775 1731 41975 1769
rect 41775 1697 41791 1731
rect 41959 1697 41975 1731
rect 41775 1681 41975 1697
rect 42147 1731 42347 1769
rect 42147 1697 42163 1731
rect 42331 1697 42347 1731
rect 42147 1681 42347 1697
rect 42519 1731 42719 1769
rect 42519 1697 42535 1731
rect 42703 1697 42719 1731
rect 42519 1681 42719 1697
rect 42891 1731 43091 1769
rect 42891 1697 42907 1731
rect 43075 1697 43091 1731
rect 42891 1681 43091 1697
rect 43263 1731 43463 1769
rect 43263 1697 43279 1731
rect 43447 1697 43463 1731
rect 43263 1681 43463 1697
rect 43635 1731 43835 1769
rect 43635 1697 43651 1731
rect 43819 1697 43835 1731
rect 43635 1681 43835 1697
rect 44007 1731 44207 1769
rect 44007 1697 44023 1731
rect 44191 1697 44207 1731
rect 44007 1681 44207 1697
rect 44379 1731 44579 1769
rect 44379 1697 44395 1731
rect 44563 1697 44579 1731
rect 44379 1681 44579 1697
rect 44751 1731 44951 1769
rect 44751 1697 44767 1731
rect 44935 1697 44951 1731
rect 44751 1681 44951 1697
rect 45123 1731 45323 1769
rect 45123 1697 45139 1731
rect 45307 1697 45323 1731
rect 45123 1681 45323 1697
rect 45495 1731 45695 1769
rect 45495 1697 45511 1731
rect 45679 1697 45695 1731
rect 45495 1681 45695 1697
rect 45867 1731 46067 1769
rect 45867 1697 45883 1731
rect 46051 1697 46067 1731
rect 45867 1681 46067 1697
rect 46239 1731 46439 1769
rect 46239 1697 46255 1731
rect 46423 1697 46439 1731
rect 46239 1681 46439 1697
rect 46611 1731 46811 1769
rect 46611 1697 46627 1731
rect 46795 1697 46811 1731
rect 46611 1681 46811 1697
rect 46983 1731 47183 1769
rect 46983 1697 46999 1731
rect 47167 1697 47183 1731
rect 46983 1681 47183 1697
rect 47355 1731 47555 1769
rect 47355 1697 47371 1731
rect 47539 1697 47555 1731
rect 47355 1681 47555 1697
rect 47727 1731 47927 1769
rect 47727 1697 47743 1731
rect 47911 1697 47927 1731
rect 47727 1681 47927 1697
rect 48099 1731 48299 1769
rect 48099 1697 48115 1731
rect 48283 1697 48299 1731
rect 48099 1681 48299 1697
rect 39543 1623 39743 1639
rect 39543 1589 39559 1623
rect 39727 1589 39743 1623
rect 39543 1551 39743 1589
rect 39915 1623 40115 1639
rect 39915 1589 39931 1623
rect 40099 1589 40115 1623
rect 39915 1551 40115 1589
rect 40287 1623 40487 1639
rect 40287 1589 40303 1623
rect 40471 1589 40487 1623
rect 40287 1551 40487 1589
rect 40659 1623 40859 1639
rect 40659 1589 40675 1623
rect 40843 1589 40859 1623
rect 40659 1551 40859 1589
rect 41031 1623 41231 1639
rect 41031 1589 41047 1623
rect 41215 1589 41231 1623
rect 41031 1551 41231 1589
rect 41403 1623 41603 1639
rect 41403 1589 41419 1623
rect 41587 1589 41603 1623
rect 41403 1551 41603 1589
rect 41775 1623 41975 1639
rect 41775 1589 41791 1623
rect 41959 1589 41975 1623
rect 41775 1551 41975 1589
rect 42147 1623 42347 1639
rect 42147 1589 42163 1623
rect 42331 1589 42347 1623
rect 42147 1551 42347 1589
rect 42519 1623 42719 1639
rect 42519 1589 42535 1623
rect 42703 1589 42719 1623
rect 42519 1551 42719 1589
rect 42891 1623 43091 1639
rect 42891 1589 42907 1623
rect 43075 1589 43091 1623
rect 42891 1551 43091 1589
rect 43263 1623 43463 1639
rect 43263 1589 43279 1623
rect 43447 1589 43463 1623
rect 43263 1551 43463 1589
rect 43635 1623 43835 1639
rect 43635 1589 43651 1623
rect 43819 1589 43835 1623
rect 43635 1551 43835 1589
rect 44007 1623 44207 1639
rect 44007 1589 44023 1623
rect 44191 1589 44207 1623
rect 44007 1551 44207 1589
rect 44379 1623 44579 1639
rect 44379 1589 44395 1623
rect 44563 1589 44579 1623
rect 44379 1551 44579 1589
rect 44751 1623 44951 1639
rect 44751 1589 44767 1623
rect 44935 1589 44951 1623
rect 44751 1551 44951 1589
rect 45123 1623 45323 1639
rect 45123 1589 45139 1623
rect 45307 1589 45323 1623
rect 45123 1551 45323 1589
rect 45495 1623 45695 1639
rect 45495 1589 45511 1623
rect 45679 1589 45695 1623
rect 45495 1551 45695 1589
rect 45867 1623 46067 1639
rect 45867 1589 45883 1623
rect 46051 1589 46067 1623
rect 45867 1551 46067 1589
rect 46239 1623 46439 1639
rect 46239 1589 46255 1623
rect 46423 1589 46439 1623
rect 46239 1551 46439 1589
rect 46611 1623 46811 1639
rect 46611 1589 46627 1623
rect 46795 1589 46811 1623
rect 46611 1551 46811 1589
rect 46983 1623 47183 1639
rect 46983 1589 46999 1623
rect 47167 1589 47183 1623
rect 46983 1551 47183 1589
rect 47355 1623 47555 1639
rect 47355 1589 47371 1623
rect 47539 1589 47555 1623
rect 47355 1551 47555 1589
rect 47727 1623 47927 1639
rect 47727 1589 47743 1623
rect 47911 1589 47927 1623
rect 47727 1551 47927 1589
rect 48099 1623 48299 1639
rect 48099 1589 48115 1623
rect 48283 1589 48299 1623
rect 48099 1551 48299 1589
rect 39543 1313 39743 1351
rect 39543 1279 39559 1313
rect 39727 1279 39743 1313
rect 39543 1263 39743 1279
rect 39915 1313 40115 1351
rect 39915 1279 39931 1313
rect 40099 1279 40115 1313
rect 39915 1263 40115 1279
rect 40287 1313 40487 1351
rect 40287 1279 40303 1313
rect 40471 1279 40487 1313
rect 40287 1263 40487 1279
rect 40659 1313 40859 1351
rect 40659 1279 40675 1313
rect 40843 1279 40859 1313
rect 40659 1263 40859 1279
rect 41031 1313 41231 1351
rect 41031 1279 41047 1313
rect 41215 1279 41231 1313
rect 41031 1263 41231 1279
rect 41403 1313 41603 1351
rect 41403 1279 41419 1313
rect 41587 1279 41603 1313
rect 41403 1263 41603 1279
rect 41775 1313 41975 1351
rect 41775 1279 41791 1313
rect 41959 1279 41975 1313
rect 41775 1263 41975 1279
rect 42147 1313 42347 1351
rect 42147 1279 42163 1313
rect 42331 1279 42347 1313
rect 42147 1263 42347 1279
rect 42519 1313 42719 1351
rect 42519 1279 42535 1313
rect 42703 1279 42719 1313
rect 42519 1263 42719 1279
rect 42891 1313 43091 1351
rect 42891 1279 42907 1313
rect 43075 1279 43091 1313
rect 42891 1263 43091 1279
rect 43263 1313 43463 1351
rect 43263 1279 43279 1313
rect 43447 1279 43463 1313
rect 43263 1263 43463 1279
rect 43635 1313 43835 1351
rect 43635 1279 43651 1313
rect 43819 1279 43835 1313
rect 43635 1263 43835 1279
rect 44007 1313 44207 1351
rect 44007 1279 44023 1313
rect 44191 1279 44207 1313
rect 44007 1263 44207 1279
rect 44379 1313 44579 1351
rect 44379 1279 44395 1313
rect 44563 1279 44579 1313
rect 44379 1263 44579 1279
rect 44751 1313 44951 1351
rect 44751 1279 44767 1313
rect 44935 1279 44951 1313
rect 44751 1263 44951 1279
rect 45123 1313 45323 1351
rect 45123 1279 45139 1313
rect 45307 1279 45323 1313
rect 45123 1263 45323 1279
rect 45495 1313 45695 1351
rect 45495 1279 45511 1313
rect 45679 1279 45695 1313
rect 45495 1263 45695 1279
rect 45867 1313 46067 1351
rect 45867 1279 45883 1313
rect 46051 1279 46067 1313
rect 45867 1263 46067 1279
rect 46239 1313 46439 1351
rect 46239 1279 46255 1313
rect 46423 1279 46439 1313
rect 46239 1263 46439 1279
rect 46611 1313 46811 1351
rect 46611 1279 46627 1313
rect 46795 1279 46811 1313
rect 46611 1263 46811 1279
rect 46983 1313 47183 1351
rect 46983 1279 46999 1313
rect 47167 1279 47183 1313
rect 46983 1263 47183 1279
rect 47355 1313 47555 1351
rect 47355 1279 47371 1313
rect 47539 1279 47555 1313
rect 47355 1263 47555 1279
rect 47727 1313 47927 1351
rect 47727 1279 47743 1313
rect 47911 1279 47927 1313
rect 47727 1263 47927 1279
rect 48099 1313 48299 1351
rect 48099 1279 48115 1313
rect 48283 1279 48299 1313
rect 48099 1263 48299 1279
rect 39543 1205 39743 1221
rect 39543 1171 39559 1205
rect 39727 1171 39743 1205
rect 39543 1133 39743 1171
rect 39915 1205 40115 1221
rect 39915 1171 39931 1205
rect 40099 1171 40115 1205
rect 39915 1133 40115 1171
rect 40287 1205 40487 1221
rect 40287 1171 40303 1205
rect 40471 1171 40487 1205
rect 40287 1133 40487 1171
rect 40659 1205 40859 1221
rect 40659 1171 40675 1205
rect 40843 1171 40859 1205
rect 40659 1133 40859 1171
rect 41031 1205 41231 1221
rect 41031 1171 41047 1205
rect 41215 1171 41231 1205
rect 41031 1133 41231 1171
rect 41403 1205 41603 1221
rect 41403 1171 41419 1205
rect 41587 1171 41603 1205
rect 41403 1133 41603 1171
rect 41775 1205 41975 1221
rect 41775 1171 41791 1205
rect 41959 1171 41975 1205
rect 41775 1133 41975 1171
rect 42147 1205 42347 1221
rect 42147 1171 42163 1205
rect 42331 1171 42347 1205
rect 42147 1133 42347 1171
rect 42519 1205 42719 1221
rect 42519 1171 42535 1205
rect 42703 1171 42719 1205
rect 42519 1133 42719 1171
rect 42891 1205 43091 1221
rect 42891 1171 42907 1205
rect 43075 1171 43091 1205
rect 42891 1133 43091 1171
rect 43263 1205 43463 1221
rect 43263 1171 43279 1205
rect 43447 1171 43463 1205
rect 43263 1133 43463 1171
rect 43635 1205 43835 1221
rect 43635 1171 43651 1205
rect 43819 1171 43835 1205
rect 43635 1133 43835 1171
rect 44007 1205 44207 1221
rect 44007 1171 44023 1205
rect 44191 1171 44207 1205
rect 44007 1133 44207 1171
rect 44379 1205 44579 1221
rect 44379 1171 44395 1205
rect 44563 1171 44579 1205
rect 44379 1133 44579 1171
rect 44751 1205 44951 1221
rect 44751 1171 44767 1205
rect 44935 1171 44951 1205
rect 44751 1133 44951 1171
rect 45123 1205 45323 1221
rect 45123 1171 45139 1205
rect 45307 1171 45323 1205
rect 45123 1133 45323 1171
rect 45495 1205 45695 1221
rect 45495 1171 45511 1205
rect 45679 1171 45695 1205
rect 45495 1133 45695 1171
rect 45867 1205 46067 1221
rect 45867 1171 45883 1205
rect 46051 1171 46067 1205
rect 45867 1133 46067 1171
rect 46239 1205 46439 1221
rect 46239 1171 46255 1205
rect 46423 1171 46439 1205
rect 46239 1133 46439 1171
rect 46611 1205 46811 1221
rect 46611 1171 46627 1205
rect 46795 1171 46811 1205
rect 46611 1133 46811 1171
rect 46983 1205 47183 1221
rect 46983 1171 46999 1205
rect 47167 1171 47183 1205
rect 46983 1133 47183 1171
rect 47355 1205 47555 1221
rect 47355 1171 47371 1205
rect 47539 1171 47555 1205
rect 47355 1133 47555 1171
rect 47727 1205 47927 1221
rect 47727 1171 47743 1205
rect 47911 1171 47927 1205
rect 47727 1133 47927 1171
rect 48099 1205 48299 1221
rect 48099 1171 48115 1205
rect 48283 1171 48299 1205
rect 48099 1133 48299 1171
rect 39543 895 39743 933
rect 39543 861 39559 895
rect 39727 861 39743 895
rect 39543 845 39743 861
rect 39915 895 40115 933
rect 39915 861 39931 895
rect 40099 861 40115 895
rect 39915 845 40115 861
rect 40287 895 40487 933
rect 40287 861 40303 895
rect 40471 861 40487 895
rect 40287 845 40487 861
rect 40659 895 40859 933
rect 40659 861 40675 895
rect 40843 861 40859 895
rect 40659 845 40859 861
rect 41031 895 41231 933
rect 41031 861 41047 895
rect 41215 861 41231 895
rect 41031 845 41231 861
rect 41403 895 41603 933
rect 41403 861 41419 895
rect 41587 861 41603 895
rect 41403 845 41603 861
rect 41775 895 41975 933
rect 41775 861 41791 895
rect 41959 861 41975 895
rect 41775 845 41975 861
rect 42147 895 42347 933
rect 42147 861 42163 895
rect 42331 861 42347 895
rect 42147 845 42347 861
rect 42519 895 42719 933
rect 42519 861 42535 895
rect 42703 861 42719 895
rect 42519 845 42719 861
rect 42891 895 43091 933
rect 42891 861 42907 895
rect 43075 861 43091 895
rect 42891 845 43091 861
rect 43263 895 43463 933
rect 43263 861 43279 895
rect 43447 861 43463 895
rect 43263 845 43463 861
rect 43635 895 43835 933
rect 43635 861 43651 895
rect 43819 861 43835 895
rect 43635 845 43835 861
rect 44007 895 44207 933
rect 44007 861 44023 895
rect 44191 861 44207 895
rect 44007 845 44207 861
rect 44379 895 44579 933
rect 44379 861 44395 895
rect 44563 861 44579 895
rect 44379 845 44579 861
rect 44751 895 44951 933
rect 44751 861 44767 895
rect 44935 861 44951 895
rect 44751 845 44951 861
rect 45123 895 45323 933
rect 45123 861 45139 895
rect 45307 861 45323 895
rect 45123 845 45323 861
rect 45495 895 45695 933
rect 45495 861 45511 895
rect 45679 861 45695 895
rect 45495 845 45695 861
rect 45867 895 46067 933
rect 45867 861 45883 895
rect 46051 861 46067 895
rect 45867 845 46067 861
rect 46239 895 46439 933
rect 46239 861 46255 895
rect 46423 861 46439 895
rect 46239 845 46439 861
rect 46611 895 46811 933
rect 46611 861 46627 895
rect 46795 861 46811 895
rect 46611 845 46811 861
rect 46983 895 47183 933
rect 46983 861 46999 895
rect 47167 861 47183 895
rect 46983 845 47183 861
rect 47355 895 47555 933
rect 47355 861 47371 895
rect 47539 861 47555 895
rect 47355 845 47555 861
rect 47727 895 47927 933
rect 47727 861 47743 895
rect 47911 861 47927 895
rect 47727 845 47927 861
rect 48099 895 48299 933
rect 48099 861 48115 895
rect 48283 861 48299 895
rect 48099 845 48299 861
rect 39543 787 39743 803
rect 39543 753 39559 787
rect 39727 753 39743 787
rect 39543 715 39743 753
rect 39915 787 40115 803
rect 39915 753 39931 787
rect 40099 753 40115 787
rect 39915 715 40115 753
rect 40287 787 40487 803
rect 40287 753 40303 787
rect 40471 753 40487 787
rect 40287 715 40487 753
rect 40659 787 40859 803
rect 40659 753 40675 787
rect 40843 753 40859 787
rect 40659 715 40859 753
rect 41031 787 41231 803
rect 41031 753 41047 787
rect 41215 753 41231 787
rect 41031 715 41231 753
rect 41403 787 41603 803
rect 41403 753 41419 787
rect 41587 753 41603 787
rect 41403 715 41603 753
rect 41775 787 41975 803
rect 41775 753 41791 787
rect 41959 753 41975 787
rect 41775 715 41975 753
rect 42147 787 42347 803
rect 42147 753 42163 787
rect 42331 753 42347 787
rect 42147 715 42347 753
rect 42519 787 42719 803
rect 42519 753 42535 787
rect 42703 753 42719 787
rect 42519 715 42719 753
rect 42891 787 43091 803
rect 42891 753 42907 787
rect 43075 753 43091 787
rect 42891 715 43091 753
rect 43263 787 43463 803
rect 43263 753 43279 787
rect 43447 753 43463 787
rect 43263 715 43463 753
rect 43635 787 43835 803
rect 43635 753 43651 787
rect 43819 753 43835 787
rect 43635 715 43835 753
rect 44007 787 44207 803
rect 44007 753 44023 787
rect 44191 753 44207 787
rect 44007 715 44207 753
rect 44379 787 44579 803
rect 44379 753 44395 787
rect 44563 753 44579 787
rect 44379 715 44579 753
rect 44751 787 44951 803
rect 44751 753 44767 787
rect 44935 753 44951 787
rect 44751 715 44951 753
rect 45123 787 45323 803
rect 45123 753 45139 787
rect 45307 753 45323 787
rect 45123 715 45323 753
rect 45495 787 45695 803
rect 45495 753 45511 787
rect 45679 753 45695 787
rect 45495 715 45695 753
rect 45867 787 46067 803
rect 45867 753 45883 787
rect 46051 753 46067 787
rect 45867 715 46067 753
rect 46239 787 46439 803
rect 46239 753 46255 787
rect 46423 753 46439 787
rect 46239 715 46439 753
rect 46611 787 46811 803
rect 46611 753 46627 787
rect 46795 753 46811 787
rect 46611 715 46811 753
rect 46983 787 47183 803
rect 46983 753 46999 787
rect 47167 753 47183 787
rect 46983 715 47183 753
rect 47355 787 47555 803
rect 47355 753 47371 787
rect 47539 753 47555 787
rect 47355 715 47555 753
rect 47727 787 47927 803
rect 47727 753 47743 787
rect 47911 753 47927 787
rect 47727 715 47927 753
rect 48099 787 48299 803
rect 48099 753 48115 787
rect 48283 753 48299 787
rect 48099 715 48299 753
rect 39543 477 39743 515
rect 39543 443 39559 477
rect 39727 443 39743 477
rect 39543 427 39743 443
rect 39915 477 40115 515
rect 39915 443 39931 477
rect 40099 443 40115 477
rect 39915 427 40115 443
rect 40287 477 40487 515
rect 40287 443 40303 477
rect 40471 443 40487 477
rect 40287 427 40487 443
rect 40659 477 40859 515
rect 40659 443 40675 477
rect 40843 443 40859 477
rect 40659 427 40859 443
rect 41031 477 41231 515
rect 41031 443 41047 477
rect 41215 443 41231 477
rect 41031 427 41231 443
rect 41403 477 41603 515
rect 41403 443 41419 477
rect 41587 443 41603 477
rect 41403 427 41603 443
rect 41775 477 41975 515
rect 41775 443 41791 477
rect 41959 443 41975 477
rect 41775 427 41975 443
rect 42147 477 42347 515
rect 42147 443 42163 477
rect 42331 443 42347 477
rect 42147 427 42347 443
rect 42519 477 42719 515
rect 42519 443 42535 477
rect 42703 443 42719 477
rect 42519 427 42719 443
rect 42891 477 43091 515
rect 42891 443 42907 477
rect 43075 443 43091 477
rect 42891 427 43091 443
rect 43263 477 43463 515
rect 43263 443 43279 477
rect 43447 443 43463 477
rect 43263 427 43463 443
rect 43635 477 43835 515
rect 43635 443 43651 477
rect 43819 443 43835 477
rect 43635 427 43835 443
rect 44007 477 44207 515
rect 44007 443 44023 477
rect 44191 443 44207 477
rect 44007 427 44207 443
rect 44379 477 44579 515
rect 44379 443 44395 477
rect 44563 443 44579 477
rect 44379 427 44579 443
rect 44751 477 44951 515
rect 44751 443 44767 477
rect 44935 443 44951 477
rect 44751 427 44951 443
rect 45123 477 45323 515
rect 45123 443 45139 477
rect 45307 443 45323 477
rect 45123 427 45323 443
rect 45495 477 45695 515
rect 45495 443 45511 477
rect 45679 443 45695 477
rect 45495 427 45695 443
rect 45867 477 46067 515
rect 45867 443 45883 477
rect 46051 443 46067 477
rect 45867 427 46067 443
rect 46239 477 46439 515
rect 46239 443 46255 477
rect 46423 443 46439 477
rect 46239 427 46439 443
rect 46611 477 46811 515
rect 46611 443 46627 477
rect 46795 443 46811 477
rect 46611 427 46811 443
rect 46983 477 47183 515
rect 46983 443 46999 477
rect 47167 443 47183 477
rect 46983 427 47183 443
rect 47355 477 47555 515
rect 47355 443 47371 477
rect 47539 443 47555 477
rect 47355 427 47555 443
rect 47727 477 47927 515
rect 47727 443 47743 477
rect 47911 443 47927 477
rect 47727 427 47927 443
rect 48099 477 48299 515
rect 48099 443 48115 477
rect 48283 443 48299 477
rect 48099 427 48299 443
<< polycont >>
rect 38071 9089 38239 9123
rect 38443 9089 38611 9123
rect 38815 9089 38983 9123
rect 39187 9089 39355 9123
rect 39559 9089 39727 9123
rect 39931 9089 40099 9123
rect 40303 9089 40471 9123
rect 40675 9089 40843 9123
rect 41047 9089 41215 9123
rect 41419 9089 41587 9123
rect 41791 9089 41959 9123
rect 42163 9089 42331 9123
rect 42535 9089 42703 9123
rect 42907 9089 43075 9123
rect 43279 9089 43447 9123
rect 43651 9089 43819 9123
rect 44023 9089 44191 9123
rect 44395 9089 44563 9123
rect 44767 9089 44935 9123
rect 45139 9089 45307 9123
rect 45511 9089 45679 9123
rect 45883 9089 46051 9123
rect 46255 9089 46423 9123
rect 46627 9089 46795 9123
rect 46999 9089 47167 9123
rect 47371 9089 47539 9123
rect 47743 9089 47911 9123
rect 48115 9089 48283 9123
rect 48487 9089 48655 9123
rect 48859 9089 49027 9123
rect 49231 9089 49399 9123
rect 49603 9089 49771 9123
rect 38071 8561 38239 8595
rect 38443 8561 38611 8595
rect 38815 8561 38983 8595
rect 39187 8561 39355 8595
rect 39559 8561 39727 8595
rect 39931 8561 40099 8595
rect 40303 8561 40471 8595
rect 40675 8561 40843 8595
rect 41047 8561 41215 8595
rect 41419 8561 41587 8595
rect 41791 8561 41959 8595
rect 42163 8561 42331 8595
rect 42535 8561 42703 8595
rect 42907 8561 43075 8595
rect 43279 8561 43447 8595
rect 43651 8561 43819 8595
rect 44023 8561 44191 8595
rect 44395 8561 44563 8595
rect 44767 8561 44935 8595
rect 45139 8561 45307 8595
rect 45511 8561 45679 8595
rect 45883 8561 46051 8595
rect 46255 8561 46423 8595
rect 46627 8561 46795 8595
rect 46999 8561 47167 8595
rect 47371 8561 47539 8595
rect 47743 8561 47911 8595
rect 48115 8561 48283 8595
rect 48487 8561 48655 8595
rect 48859 8561 49027 8595
rect 49231 8561 49399 8595
rect 49603 8561 49771 8595
rect 38071 8453 38239 8487
rect 38443 8453 38611 8487
rect 38815 8453 38983 8487
rect 39187 8453 39355 8487
rect 39559 8453 39727 8487
rect 39931 8453 40099 8487
rect 40303 8453 40471 8487
rect 40675 8453 40843 8487
rect 41047 8453 41215 8487
rect 41419 8453 41587 8487
rect 41791 8453 41959 8487
rect 42163 8453 42331 8487
rect 42535 8453 42703 8487
rect 42907 8453 43075 8487
rect 43279 8453 43447 8487
rect 43651 8453 43819 8487
rect 44023 8453 44191 8487
rect 44395 8453 44563 8487
rect 44767 8453 44935 8487
rect 45139 8453 45307 8487
rect 45511 8453 45679 8487
rect 45883 8453 46051 8487
rect 46255 8453 46423 8487
rect 46627 8453 46795 8487
rect 46999 8453 47167 8487
rect 47371 8453 47539 8487
rect 47743 8453 47911 8487
rect 48115 8453 48283 8487
rect 48487 8453 48655 8487
rect 48859 8453 49027 8487
rect 49231 8453 49399 8487
rect 49603 8453 49771 8487
rect 38071 7925 38239 7959
rect 38443 7925 38611 7959
rect 38815 7925 38983 7959
rect 39187 7925 39355 7959
rect 39559 7925 39727 7959
rect 39931 7925 40099 7959
rect 40303 7925 40471 7959
rect 40675 7925 40843 7959
rect 41047 7925 41215 7959
rect 41419 7925 41587 7959
rect 41791 7925 41959 7959
rect 42163 7925 42331 7959
rect 42535 7925 42703 7959
rect 42907 7925 43075 7959
rect 43279 7925 43447 7959
rect 43651 7925 43819 7959
rect 44023 7925 44191 7959
rect 44395 7925 44563 7959
rect 44767 7925 44935 7959
rect 45139 7925 45307 7959
rect 45511 7925 45679 7959
rect 45883 7925 46051 7959
rect 46255 7925 46423 7959
rect 46627 7925 46795 7959
rect 46999 7925 47167 7959
rect 47371 7925 47539 7959
rect 47743 7925 47911 7959
rect 48115 7925 48283 7959
rect 48487 7925 48655 7959
rect 48859 7925 49027 7959
rect 49231 7925 49399 7959
rect 49603 7925 49771 7959
rect 38071 7817 38239 7851
rect 38443 7817 38611 7851
rect 38815 7817 38983 7851
rect 39187 7817 39355 7851
rect 39559 7817 39727 7851
rect 39931 7817 40099 7851
rect 40303 7817 40471 7851
rect 40675 7817 40843 7851
rect 41047 7817 41215 7851
rect 41419 7817 41587 7851
rect 41791 7817 41959 7851
rect 42163 7817 42331 7851
rect 42535 7817 42703 7851
rect 42907 7817 43075 7851
rect 43279 7817 43447 7851
rect 43651 7817 43819 7851
rect 44023 7817 44191 7851
rect 44395 7817 44563 7851
rect 44767 7817 44935 7851
rect 45139 7817 45307 7851
rect 45511 7817 45679 7851
rect 45883 7817 46051 7851
rect 46255 7817 46423 7851
rect 46627 7817 46795 7851
rect 46999 7817 47167 7851
rect 47371 7817 47539 7851
rect 47743 7817 47911 7851
rect 48115 7817 48283 7851
rect 48487 7817 48655 7851
rect 48859 7817 49027 7851
rect 49231 7817 49399 7851
rect 49603 7817 49771 7851
rect 38071 7289 38239 7323
rect 38443 7289 38611 7323
rect 38815 7289 38983 7323
rect 39187 7289 39355 7323
rect 39559 7289 39727 7323
rect 39931 7289 40099 7323
rect 40303 7289 40471 7323
rect 40675 7289 40843 7323
rect 41047 7289 41215 7323
rect 41419 7289 41587 7323
rect 41791 7289 41959 7323
rect 42163 7289 42331 7323
rect 42535 7289 42703 7323
rect 42907 7289 43075 7323
rect 43279 7289 43447 7323
rect 43651 7289 43819 7323
rect 44023 7289 44191 7323
rect 44395 7289 44563 7323
rect 44767 7289 44935 7323
rect 45139 7289 45307 7323
rect 45511 7289 45679 7323
rect 45883 7289 46051 7323
rect 46255 7289 46423 7323
rect 46627 7289 46795 7323
rect 46999 7289 47167 7323
rect 47371 7289 47539 7323
rect 47743 7289 47911 7323
rect 48115 7289 48283 7323
rect 48487 7289 48655 7323
rect 48859 7289 49027 7323
rect 49231 7289 49399 7323
rect 49603 7289 49771 7323
rect 39559 6701 39727 6735
rect 39931 6701 40099 6735
rect 40303 6701 40471 6735
rect 40675 6701 40843 6735
rect 41047 6701 41215 6735
rect 41419 6701 41587 6735
rect 41791 6701 41959 6735
rect 42163 6701 42331 6735
rect 39559 5773 39727 5807
rect 39931 5773 40099 5807
rect 40303 5773 40471 5807
rect 40675 5773 40843 5807
rect 41047 5773 41215 5807
rect 41419 5773 41587 5807
rect 41791 5773 41959 5807
rect 42163 5773 42331 5807
rect 39559 5665 39727 5699
rect 39931 5665 40099 5699
rect 40303 5665 40471 5699
rect 40675 5665 40843 5699
rect 41047 5665 41215 5699
rect 41419 5665 41587 5699
rect 41791 5665 41959 5699
rect 42163 5665 42331 5699
rect 39559 4737 39727 4771
rect 39931 4737 40099 4771
rect 40303 4737 40471 4771
rect 40675 4737 40843 4771
rect 41047 4737 41215 4771
rect 41419 4737 41587 4771
rect 41791 4737 41959 4771
rect 42163 4737 42331 4771
rect 39559 4629 39727 4663
rect 39931 4629 40099 4663
rect 40303 4629 40471 4663
rect 40675 4629 40843 4663
rect 41047 4629 41215 4663
rect 41419 4629 41587 4663
rect 41791 4629 41959 4663
rect 42163 4629 42331 4663
rect 39559 3701 39727 3735
rect 39931 3701 40099 3735
rect 40303 3701 40471 3735
rect 40675 3701 40843 3735
rect 41047 3701 41215 3735
rect 41419 3701 41587 3735
rect 41791 3701 41959 3735
rect 42163 3701 42331 3735
rect 39559 3593 39727 3627
rect 39931 3593 40099 3627
rect 40303 3593 40471 3627
rect 40675 3593 40843 3627
rect 41047 3593 41215 3627
rect 41419 3593 41587 3627
rect 41791 3593 41959 3627
rect 42163 3593 42331 3627
rect 39559 2665 39727 2699
rect 39931 2665 40099 2699
rect 40303 2665 40471 2699
rect 40675 2665 40843 2699
rect 41047 2665 41215 2699
rect 41419 2665 41587 2699
rect 41791 2665 41959 2699
rect 42163 2665 42331 2699
rect 39559 2007 39727 2041
rect 39931 2007 40099 2041
rect 40303 2007 40471 2041
rect 40675 2007 40843 2041
rect 41047 2007 41215 2041
rect 41419 2007 41587 2041
rect 41791 2007 41959 2041
rect 42163 2007 42331 2041
rect 42535 2007 42703 2041
rect 42907 2007 43075 2041
rect 43279 2007 43447 2041
rect 43651 2007 43819 2041
rect 44023 2007 44191 2041
rect 44395 2007 44563 2041
rect 44767 2007 44935 2041
rect 45139 2007 45307 2041
rect 45511 2007 45679 2041
rect 45883 2007 46051 2041
rect 46255 2007 46423 2041
rect 46627 2007 46795 2041
rect 46999 2007 47167 2041
rect 47371 2007 47539 2041
rect 47743 2007 47911 2041
rect 48115 2007 48283 2041
rect 39559 1697 39727 1731
rect 39931 1697 40099 1731
rect 40303 1697 40471 1731
rect 40675 1697 40843 1731
rect 41047 1697 41215 1731
rect 41419 1697 41587 1731
rect 41791 1697 41959 1731
rect 42163 1697 42331 1731
rect 42535 1697 42703 1731
rect 42907 1697 43075 1731
rect 43279 1697 43447 1731
rect 43651 1697 43819 1731
rect 44023 1697 44191 1731
rect 44395 1697 44563 1731
rect 44767 1697 44935 1731
rect 45139 1697 45307 1731
rect 45511 1697 45679 1731
rect 45883 1697 46051 1731
rect 46255 1697 46423 1731
rect 46627 1697 46795 1731
rect 46999 1697 47167 1731
rect 47371 1697 47539 1731
rect 47743 1697 47911 1731
rect 48115 1697 48283 1731
rect 39559 1589 39727 1623
rect 39931 1589 40099 1623
rect 40303 1589 40471 1623
rect 40675 1589 40843 1623
rect 41047 1589 41215 1623
rect 41419 1589 41587 1623
rect 41791 1589 41959 1623
rect 42163 1589 42331 1623
rect 42535 1589 42703 1623
rect 42907 1589 43075 1623
rect 43279 1589 43447 1623
rect 43651 1589 43819 1623
rect 44023 1589 44191 1623
rect 44395 1589 44563 1623
rect 44767 1589 44935 1623
rect 45139 1589 45307 1623
rect 45511 1589 45679 1623
rect 45883 1589 46051 1623
rect 46255 1589 46423 1623
rect 46627 1589 46795 1623
rect 46999 1589 47167 1623
rect 47371 1589 47539 1623
rect 47743 1589 47911 1623
rect 48115 1589 48283 1623
rect 39559 1279 39727 1313
rect 39931 1279 40099 1313
rect 40303 1279 40471 1313
rect 40675 1279 40843 1313
rect 41047 1279 41215 1313
rect 41419 1279 41587 1313
rect 41791 1279 41959 1313
rect 42163 1279 42331 1313
rect 42535 1279 42703 1313
rect 42907 1279 43075 1313
rect 43279 1279 43447 1313
rect 43651 1279 43819 1313
rect 44023 1279 44191 1313
rect 44395 1279 44563 1313
rect 44767 1279 44935 1313
rect 45139 1279 45307 1313
rect 45511 1279 45679 1313
rect 45883 1279 46051 1313
rect 46255 1279 46423 1313
rect 46627 1279 46795 1313
rect 46999 1279 47167 1313
rect 47371 1279 47539 1313
rect 47743 1279 47911 1313
rect 48115 1279 48283 1313
rect 39559 1171 39727 1205
rect 39931 1171 40099 1205
rect 40303 1171 40471 1205
rect 40675 1171 40843 1205
rect 41047 1171 41215 1205
rect 41419 1171 41587 1205
rect 41791 1171 41959 1205
rect 42163 1171 42331 1205
rect 42535 1171 42703 1205
rect 42907 1171 43075 1205
rect 43279 1171 43447 1205
rect 43651 1171 43819 1205
rect 44023 1171 44191 1205
rect 44395 1171 44563 1205
rect 44767 1171 44935 1205
rect 45139 1171 45307 1205
rect 45511 1171 45679 1205
rect 45883 1171 46051 1205
rect 46255 1171 46423 1205
rect 46627 1171 46795 1205
rect 46999 1171 47167 1205
rect 47371 1171 47539 1205
rect 47743 1171 47911 1205
rect 48115 1171 48283 1205
rect 39559 861 39727 895
rect 39931 861 40099 895
rect 40303 861 40471 895
rect 40675 861 40843 895
rect 41047 861 41215 895
rect 41419 861 41587 895
rect 41791 861 41959 895
rect 42163 861 42331 895
rect 42535 861 42703 895
rect 42907 861 43075 895
rect 43279 861 43447 895
rect 43651 861 43819 895
rect 44023 861 44191 895
rect 44395 861 44563 895
rect 44767 861 44935 895
rect 45139 861 45307 895
rect 45511 861 45679 895
rect 45883 861 46051 895
rect 46255 861 46423 895
rect 46627 861 46795 895
rect 46999 861 47167 895
rect 47371 861 47539 895
rect 47743 861 47911 895
rect 48115 861 48283 895
rect 39559 753 39727 787
rect 39931 753 40099 787
rect 40303 753 40471 787
rect 40675 753 40843 787
rect 41047 753 41215 787
rect 41419 753 41587 787
rect 41791 753 41959 787
rect 42163 753 42331 787
rect 42535 753 42703 787
rect 42907 753 43075 787
rect 43279 753 43447 787
rect 43651 753 43819 787
rect 44023 753 44191 787
rect 44395 753 44563 787
rect 44767 753 44935 787
rect 45139 753 45307 787
rect 45511 753 45679 787
rect 45883 753 46051 787
rect 46255 753 46423 787
rect 46627 753 46795 787
rect 46999 753 47167 787
rect 47371 753 47539 787
rect 47743 753 47911 787
rect 48115 753 48283 787
rect 39559 443 39727 477
rect 39931 443 40099 477
rect 40303 443 40471 477
rect 40675 443 40843 477
rect 41047 443 41215 477
rect 41419 443 41587 477
rect 41791 443 41959 477
rect 42163 443 42331 477
rect 42535 443 42703 477
rect 42907 443 43075 477
rect 43279 443 43447 477
rect 43651 443 43819 477
rect 44023 443 44191 477
rect 44395 443 44563 477
rect 44767 443 44935 477
rect 45139 443 45307 477
rect 45511 443 45679 477
rect 45883 443 46051 477
rect 46255 443 46423 477
rect 46627 443 46795 477
rect 46999 443 47167 477
rect 47371 443 47539 477
rect 47743 443 47911 477
rect 48115 443 48283 477
<< xpolycontact >>
rect 43139 4361 43209 4793
rect 43139 3369 43209 3801
<< xpolyres >>
rect 43139 3801 43209 4361
<< locali >>
rect 37895 9191 37991 9225
rect 49854 9191 49947 9225
rect 37895 9129 37929 9191
rect 49913 9129 49947 9191
rect 38055 9089 38071 9123
rect 38239 9089 38255 9123
rect 38427 9089 38443 9123
rect 38611 9089 38627 9123
rect 38799 9089 38815 9123
rect 38983 9089 38999 9123
rect 39171 9089 39187 9123
rect 39355 9089 39371 9123
rect 39543 9089 39559 9123
rect 39727 9089 39743 9123
rect 39915 9089 39931 9123
rect 40099 9089 40115 9123
rect 40287 9089 40303 9123
rect 40471 9089 40487 9123
rect 40659 9089 40675 9123
rect 40843 9089 40859 9123
rect 41031 9089 41047 9123
rect 41215 9089 41231 9123
rect 41403 9089 41419 9123
rect 41587 9089 41603 9123
rect 41775 9089 41791 9123
rect 41959 9089 41975 9123
rect 42147 9089 42163 9123
rect 42331 9089 42347 9123
rect 42519 9089 42535 9123
rect 42703 9089 42719 9123
rect 42891 9089 42907 9123
rect 43075 9089 43091 9123
rect 43263 9089 43279 9123
rect 43447 9089 43463 9123
rect 43635 9089 43651 9123
rect 43819 9089 43835 9123
rect 44007 9089 44023 9123
rect 44191 9089 44207 9123
rect 44379 9089 44395 9123
rect 44563 9089 44579 9123
rect 44751 9089 44767 9123
rect 44935 9089 44951 9123
rect 45123 9089 45139 9123
rect 45307 9089 45323 9123
rect 45495 9089 45511 9123
rect 45679 9089 45695 9123
rect 45867 9089 45883 9123
rect 46051 9089 46067 9123
rect 46239 9089 46255 9123
rect 46423 9089 46439 9123
rect 46611 9089 46627 9123
rect 46795 9089 46811 9123
rect 46983 9089 46999 9123
rect 47167 9089 47183 9123
rect 47355 9089 47371 9123
rect 47539 9089 47555 9123
rect 47727 9089 47743 9123
rect 47911 9089 47927 9123
rect 48099 9089 48115 9123
rect 48283 9089 48299 9123
rect 48471 9089 48487 9123
rect 48655 9089 48671 9123
rect 48843 9089 48859 9123
rect 49027 9089 49043 9123
rect 49215 9089 49231 9123
rect 49399 9089 49415 9123
rect 49587 9089 49603 9123
rect 49771 9089 49787 9123
rect 38009 9030 38043 9046
rect 38009 8638 38043 8654
rect 38267 9030 38301 9046
rect 38267 8638 38301 8654
rect 38381 9030 38415 9046
rect 38381 8638 38415 8654
rect 38639 9030 38673 9046
rect 38639 8638 38673 8654
rect 38753 9030 38787 9046
rect 38753 8638 38787 8654
rect 39011 9030 39045 9046
rect 39011 8638 39045 8654
rect 39125 9030 39159 9046
rect 39125 8638 39159 8654
rect 39383 9030 39417 9046
rect 39383 8638 39417 8654
rect 39497 9030 39531 9046
rect 39497 8638 39531 8654
rect 39755 9030 39789 9046
rect 39755 8638 39789 8654
rect 39869 9030 39903 9046
rect 39869 8638 39903 8654
rect 40127 9030 40161 9046
rect 40127 8638 40161 8654
rect 40241 9030 40275 9046
rect 40241 8638 40275 8654
rect 40499 9030 40533 9046
rect 40499 8638 40533 8654
rect 40613 9030 40647 9046
rect 40613 8638 40647 8654
rect 40871 9030 40905 9046
rect 40871 8638 40905 8654
rect 40985 9030 41019 9046
rect 40985 8638 41019 8654
rect 41243 9030 41277 9046
rect 41243 8638 41277 8654
rect 41357 9030 41391 9046
rect 41357 8638 41391 8654
rect 41615 9030 41649 9046
rect 41615 8638 41649 8654
rect 41729 9030 41763 9046
rect 41729 8638 41763 8654
rect 41987 9030 42021 9046
rect 41987 8638 42021 8654
rect 42101 9030 42135 9046
rect 42101 8638 42135 8654
rect 42359 9030 42393 9046
rect 42359 8638 42393 8654
rect 42473 9030 42507 9046
rect 42473 8638 42507 8654
rect 42731 9030 42765 9046
rect 42731 8638 42765 8654
rect 42845 9030 42879 9046
rect 42845 8638 42879 8654
rect 43103 9030 43137 9046
rect 43103 8638 43137 8654
rect 43217 9030 43251 9046
rect 43217 8638 43251 8654
rect 43475 9030 43509 9046
rect 43475 8638 43509 8654
rect 43589 9030 43623 9046
rect 43589 8638 43623 8654
rect 43847 9030 43881 9046
rect 43847 8638 43881 8654
rect 43961 9030 43995 9046
rect 43961 8638 43995 8654
rect 44219 9030 44253 9046
rect 44219 8638 44253 8654
rect 44333 9030 44367 9046
rect 44333 8638 44367 8654
rect 44591 9030 44625 9046
rect 44591 8638 44625 8654
rect 44705 9030 44739 9046
rect 44705 8638 44739 8654
rect 44963 9030 44997 9046
rect 44963 8638 44997 8654
rect 45077 9030 45111 9046
rect 45077 8638 45111 8654
rect 45335 9030 45369 9046
rect 45335 8638 45369 8654
rect 45449 9030 45483 9046
rect 45449 8638 45483 8654
rect 45707 9030 45741 9046
rect 45707 8638 45741 8654
rect 45821 9030 45855 9046
rect 45821 8638 45855 8654
rect 46079 9030 46113 9046
rect 46079 8638 46113 8654
rect 46193 9030 46227 9046
rect 46193 8638 46227 8654
rect 46451 9030 46485 9046
rect 46451 8638 46485 8654
rect 46565 9030 46599 9046
rect 46565 8638 46599 8654
rect 46823 9030 46857 9046
rect 46823 8638 46857 8654
rect 46937 9030 46971 9046
rect 46937 8638 46971 8654
rect 47195 9030 47229 9046
rect 47195 8638 47229 8654
rect 47309 9030 47343 9046
rect 47309 8638 47343 8654
rect 47567 9030 47601 9046
rect 47567 8638 47601 8654
rect 47681 9030 47715 9046
rect 47681 8638 47715 8654
rect 47939 9030 47973 9046
rect 47939 8638 47973 8654
rect 48053 9030 48087 9046
rect 48053 8638 48087 8654
rect 48311 9030 48345 9046
rect 48311 8638 48345 8654
rect 48425 9030 48459 9046
rect 48425 8638 48459 8654
rect 48683 9030 48717 9046
rect 48683 8638 48717 8654
rect 48797 9030 48831 9046
rect 48797 8638 48831 8654
rect 49055 9030 49089 9046
rect 49055 8638 49089 8654
rect 49169 9030 49203 9046
rect 49169 8638 49203 8654
rect 49427 9030 49461 9046
rect 49427 8638 49461 8654
rect 49541 9030 49575 9046
rect 49541 8638 49575 8654
rect 49799 9030 49833 9046
rect 49799 8638 49833 8654
rect 38055 8561 38071 8595
rect 38239 8561 38255 8595
rect 38427 8561 38443 8595
rect 38611 8561 38627 8595
rect 38799 8561 38815 8595
rect 38983 8561 38999 8595
rect 39171 8561 39187 8595
rect 39355 8561 39371 8595
rect 39543 8561 39559 8595
rect 39727 8561 39743 8595
rect 39915 8561 39931 8595
rect 40099 8561 40115 8595
rect 40287 8561 40303 8595
rect 40471 8561 40487 8595
rect 40659 8561 40675 8595
rect 40843 8561 40859 8595
rect 41031 8561 41047 8595
rect 41215 8561 41231 8595
rect 41403 8561 41419 8595
rect 41587 8561 41603 8595
rect 41775 8561 41791 8595
rect 41959 8561 41975 8595
rect 42147 8561 42163 8595
rect 42331 8561 42347 8595
rect 42519 8561 42535 8595
rect 42703 8561 42719 8595
rect 42891 8561 42907 8595
rect 43075 8561 43091 8595
rect 43263 8561 43279 8595
rect 43447 8561 43463 8595
rect 43635 8561 43651 8595
rect 43819 8561 43835 8595
rect 44007 8561 44023 8595
rect 44191 8561 44207 8595
rect 44379 8561 44395 8595
rect 44563 8561 44579 8595
rect 44751 8561 44767 8595
rect 44935 8561 44951 8595
rect 45123 8561 45139 8595
rect 45307 8561 45323 8595
rect 45495 8561 45511 8595
rect 45679 8561 45695 8595
rect 45867 8561 45883 8595
rect 46051 8561 46067 8595
rect 46239 8561 46255 8595
rect 46423 8561 46439 8595
rect 46611 8561 46627 8595
rect 46795 8561 46811 8595
rect 46983 8561 46999 8595
rect 47167 8561 47183 8595
rect 47355 8561 47371 8595
rect 47539 8561 47555 8595
rect 47727 8561 47743 8595
rect 47911 8561 47927 8595
rect 48099 8561 48115 8595
rect 48283 8561 48299 8595
rect 48471 8561 48487 8595
rect 48655 8561 48671 8595
rect 48843 8561 48859 8595
rect 49027 8561 49043 8595
rect 49215 8561 49231 8595
rect 49399 8561 49415 8595
rect 49587 8561 49603 8595
rect 49771 8561 49787 8595
rect 38055 8453 38071 8487
rect 38239 8453 38255 8487
rect 38427 8453 38443 8487
rect 38611 8453 38627 8487
rect 38799 8453 38815 8487
rect 38983 8453 38999 8487
rect 39171 8453 39187 8487
rect 39355 8453 39371 8487
rect 39543 8453 39559 8487
rect 39727 8453 39743 8487
rect 39915 8453 39931 8487
rect 40099 8453 40115 8487
rect 40287 8453 40303 8487
rect 40471 8453 40487 8487
rect 40659 8453 40675 8487
rect 40843 8453 40859 8487
rect 41031 8453 41047 8487
rect 41215 8453 41231 8487
rect 41403 8453 41419 8487
rect 41587 8453 41603 8487
rect 41775 8453 41791 8487
rect 41959 8453 41975 8487
rect 42147 8453 42163 8487
rect 42331 8453 42347 8487
rect 42519 8453 42535 8487
rect 42703 8453 42719 8487
rect 42891 8453 42907 8487
rect 43075 8453 43091 8487
rect 43263 8453 43279 8487
rect 43447 8453 43463 8487
rect 43635 8453 43651 8487
rect 43819 8453 43835 8487
rect 44007 8453 44023 8487
rect 44191 8453 44207 8487
rect 44379 8453 44395 8487
rect 44563 8453 44579 8487
rect 44751 8453 44767 8487
rect 44935 8453 44951 8487
rect 45123 8453 45139 8487
rect 45307 8453 45323 8487
rect 45495 8453 45511 8487
rect 45679 8453 45695 8487
rect 45867 8453 45883 8487
rect 46051 8453 46067 8487
rect 46239 8453 46255 8487
rect 46423 8453 46439 8487
rect 46611 8453 46627 8487
rect 46795 8453 46811 8487
rect 46983 8453 46999 8487
rect 47167 8453 47183 8487
rect 47355 8453 47371 8487
rect 47539 8453 47555 8487
rect 47727 8453 47743 8487
rect 47911 8453 47927 8487
rect 48099 8453 48115 8487
rect 48283 8453 48299 8487
rect 48471 8453 48487 8487
rect 48655 8453 48671 8487
rect 48843 8453 48859 8487
rect 49027 8453 49043 8487
rect 49215 8453 49231 8487
rect 49399 8453 49415 8487
rect 49587 8453 49603 8487
rect 49771 8453 49787 8487
rect 38009 8394 38043 8410
rect 38009 8002 38043 8018
rect 38267 8394 38301 8410
rect 38267 8002 38301 8018
rect 38381 8394 38415 8410
rect 38381 8002 38415 8018
rect 38639 8394 38673 8410
rect 38639 8002 38673 8018
rect 38753 8394 38787 8410
rect 38753 8002 38787 8018
rect 39011 8394 39045 8410
rect 39011 8002 39045 8018
rect 39125 8394 39159 8410
rect 39125 8002 39159 8018
rect 39383 8394 39417 8410
rect 39383 8002 39417 8018
rect 39497 8394 39531 8410
rect 39497 8002 39531 8018
rect 39755 8394 39789 8410
rect 39755 8002 39789 8018
rect 39869 8394 39903 8410
rect 39869 8002 39903 8018
rect 40127 8394 40161 8410
rect 40127 8002 40161 8018
rect 40241 8394 40275 8410
rect 40241 8002 40275 8018
rect 40499 8394 40533 8410
rect 40499 8002 40533 8018
rect 40613 8394 40647 8410
rect 40613 8002 40647 8018
rect 40871 8394 40905 8410
rect 40871 8002 40905 8018
rect 40985 8394 41019 8410
rect 40985 8002 41019 8018
rect 41243 8394 41277 8410
rect 41243 8002 41277 8018
rect 41357 8394 41391 8410
rect 41357 8002 41391 8018
rect 41615 8394 41649 8410
rect 41615 8002 41649 8018
rect 41729 8394 41763 8410
rect 41729 8002 41763 8018
rect 41987 8394 42021 8410
rect 41987 8002 42021 8018
rect 42101 8394 42135 8410
rect 42101 8002 42135 8018
rect 42359 8394 42393 8410
rect 42359 8002 42393 8018
rect 42473 8394 42507 8410
rect 42473 8002 42507 8018
rect 42731 8394 42765 8410
rect 42731 8002 42765 8018
rect 42845 8394 42879 8410
rect 42845 8002 42879 8018
rect 43103 8394 43137 8410
rect 43103 8002 43137 8018
rect 43217 8394 43251 8410
rect 43217 8002 43251 8018
rect 43475 8394 43509 8410
rect 43475 8002 43509 8018
rect 43589 8394 43623 8410
rect 43589 8002 43623 8018
rect 43847 8394 43881 8410
rect 43847 8002 43881 8018
rect 43961 8394 43995 8410
rect 43961 8002 43995 8018
rect 44219 8394 44253 8410
rect 44219 8002 44253 8018
rect 44333 8394 44367 8410
rect 44333 8002 44367 8018
rect 44591 8394 44625 8410
rect 44591 8002 44625 8018
rect 44705 8394 44739 8410
rect 44705 8002 44739 8018
rect 44963 8394 44997 8410
rect 44963 8002 44997 8018
rect 45077 8394 45111 8410
rect 45077 8002 45111 8018
rect 45335 8394 45369 8410
rect 45335 8002 45369 8018
rect 45449 8394 45483 8410
rect 45449 8002 45483 8018
rect 45707 8394 45741 8410
rect 45707 8002 45741 8018
rect 45821 8394 45855 8410
rect 45821 8002 45855 8018
rect 46079 8394 46113 8410
rect 46079 8002 46113 8018
rect 46193 8394 46227 8410
rect 46193 8002 46227 8018
rect 46451 8394 46485 8410
rect 46451 8002 46485 8018
rect 46565 8394 46599 8410
rect 46565 8002 46599 8018
rect 46823 8394 46857 8410
rect 46823 8002 46857 8018
rect 46937 8394 46971 8410
rect 46937 8002 46971 8018
rect 47195 8394 47229 8410
rect 47195 8002 47229 8018
rect 47309 8394 47343 8410
rect 47309 8002 47343 8018
rect 47567 8394 47601 8410
rect 47567 8002 47601 8018
rect 47681 8394 47715 8410
rect 47681 8002 47715 8018
rect 47939 8394 47973 8410
rect 47939 8002 47973 8018
rect 48053 8394 48087 8410
rect 48053 8002 48087 8018
rect 48311 8394 48345 8410
rect 48311 8002 48345 8018
rect 48425 8394 48459 8410
rect 48425 8002 48459 8018
rect 48683 8394 48717 8410
rect 48683 8002 48717 8018
rect 48797 8394 48831 8410
rect 48797 8002 48831 8018
rect 49055 8394 49089 8410
rect 49055 8002 49089 8018
rect 49169 8394 49203 8410
rect 49169 8002 49203 8018
rect 49427 8394 49461 8410
rect 49427 8002 49461 8018
rect 49541 8394 49575 8410
rect 49541 8002 49575 8018
rect 49799 8394 49833 8410
rect 49799 8002 49833 8018
rect 38055 7925 38071 7959
rect 38239 7925 38255 7959
rect 38427 7925 38443 7959
rect 38611 7925 38627 7959
rect 38799 7925 38815 7959
rect 38983 7925 38999 7959
rect 39171 7925 39187 7959
rect 39355 7925 39371 7959
rect 39543 7925 39559 7959
rect 39727 7925 39743 7959
rect 39915 7925 39931 7959
rect 40099 7925 40115 7959
rect 40287 7925 40303 7959
rect 40471 7925 40487 7959
rect 40659 7925 40675 7959
rect 40843 7925 40859 7959
rect 41031 7925 41047 7959
rect 41215 7925 41231 7959
rect 41403 7925 41419 7959
rect 41587 7925 41603 7959
rect 41775 7925 41791 7959
rect 41959 7925 41975 7959
rect 42147 7925 42163 7959
rect 42331 7925 42347 7959
rect 42519 7925 42535 7959
rect 42703 7925 42719 7959
rect 42891 7925 42907 7959
rect 43075 7925 43091 7959
rect 43263 7925 43279 7959
rect 43447 7925 43463 7959
rect 43635 7925 43651 7959
rect 43819 7925 43835 7959
rect 44007 7925 44023 7959
rect 44191 7925 44207 7959
rect 44379 7925 44395 7959
rect 44563 7925 44579 7959
rect 44751 7925 44767 7959
rect 44935 7925 44951 7959
rect 45123 7925 45139 7959
rect 45307 7925 45323 7959
rect 45495 7925 45511 7959
rect 45679 7925 45695 7959
rect 45867 7925 45883 7959
rect 46051 7925 46067 7959
rect 46239 7925 46255 7959
rect 46423 7925 46439 7959
rect 46611 7925 46627 7959
rect 46795 7925 46811 7959
rect 46983 7925 46999 7959
rect 47167 7925 47183 7959
rect 47355 7925 47371 7959
rect 47539 7925 47555 7959
rect 47727 7925 47743 7959
rect 47911 7925 47927 7959
rect 48099 7925 48115 7959
rect 48283 7925 48299 7959
rect 48471 7925 48487 7959
rect 48655 7925 48671 7959
rect 48843 7925 48859 7959
rect 49027 7925 49043 7959
rect 49215 7925 49231 7959
rect 49399 7925 49415 7959
rect 49587 7925 49603 7959
rect 49771 7925 49787 7959
rect 38055 7817 38071 7851
rect 38239 7817 38255 7851
rect 38427 7817 38443 7851
rect 38611 7817 38627 7851
rect 38799 7817 38815 7851
rect 38983 7817 38999 7851
rect 39171 7817 39187 7851
rect 39355 7817 39371 7851
rect 39543 7817 39559 7851
rect 39727 7817 39743 7851
rect 39915 7817 39931 7851
rect 40099 7817 40115 7851
rect 40287 7817 40303 7851
rect 40471 7817 40487 7851
rect 40659 7817 40675 7851
rect 40843 7817 40859 7851
rect 41031 7817 41047 7851
rect 41215 7817 41231 7851
rect 41403 7817 41419 7851
rect 41587 7817 41603 7851
rect 41775 7817 41791 7851
rect 41959 7817 41975 7851
rect 42147 7817 42163 7851
rect 42331 7817 42347 7851
rect 42519 7817 42535 7851
rect 42703 7817 42719 7851
rect 42891 7817 42907 7851
rect 43075 7817 43091 7851
rect 43263 7817 43279 7851
rect 43447 7817 43463 7851
rect 43635 7817 43651 7851
rect 43819 7817 43835 7851
rect 44007 7817 44023 7851
rect 44191 7817 44207 7851
rect 44379 7817 44395 7851
rect 44563 7817 44579 7851
rect 44751 7817 44767 7851
rect 44935 7817 44951 7851
rect 45123 7817 45139 7851
rect 45307 7817 45323 7851
rect 45495 7817 45511 7851
rect 45679 7817 45695 7851
rect 45867 7817 45883 7851
rect 46051 7817 46067 7851
rect 46239 7817 46255 7851
rect 46423 7817 46439 7851
rect 46611 7817 46627 7851
rect 46795 7817 46811 7851
rect 46983 7817 46999 7851
rect 47167 7817 47183 7851
rect 47355 7817 47371 7851
rect 47539 7817 47555 7851
rect 47727 7817 47743 7851
rect 47911 7817 47927 7851
rect 48099 7817 48115 7851
rect 48283 7817 48299 7851
rect 48471 7817 48487 7851
rect 48655 7817 48671 7851
rect 48843 7817 48859 7851
rect 49027 7817 49043 7851
rect 49215 7817 49231 7851
rect 49399 7817 49415 7851
rect 49587 7817 49603 7851
rect 49771 7817 49787 7851
rect 38009 7758 38043 7774
rect 38009 7366 38043 7382
rect 38267 7758 38301 7774
rect 38267 7366 38301 7382
rect 38381 7758 38415 7774
rect 38381 7366 38415 7382
rect 38639 7758 38673 7774
rect 38639 7366 38673 7382
rect 38753 7758 38787 7774
rect 38753 7366 38787 7382
rect 39011 7758 39045 7774
rect 39011 7366 39045 7382
rect 39125 7758 39159 7774
rect 39125 7366 39159 7382
rect 39383 7758 39417 7774
rect 39383 7366 39417 7382
rect 39497 7758 39531 7774
rect 39497 7366 39531 7382
rect 39755 7758 39789 7774
rect 39755 7366 39789 7382
rect 39869 7758 39903 7774
rect 39869 7366 39903 7382
rect 40127 7758 40161 7774
rect 40127 7366 40161 7382
rect 40241 7758 40275 7774
rect 40241 7366 40275 7382
rect 40499 7758 40533 7774
rect 40499 7366 40533 7382
rect 40613 7758 40647 7774
rect 40613 7366 40647 7382
rect 40871 7758 40905 7774
rect 40871 7366 40905 7382
rect 40985 7758 41019 7774
rect 40985 7366 41019 7382
rect 41243 7758 41277 7774
rect 41243 7366 41277 7382
rect 41357 7758 41391 7774
rect 41357 7366 41391 7382
rect 41615 7758 41649 7774
rect 41615 7366 41649 7382
rect 41729 7758 41763 7774
rect 41729 7366 41763 7382
rect 41987 7758 42021 7774
rect 41987 7366 42021 7382
rect 42101 7758 42135 7774
rect 42101 7366 42135 7382
rect 42359 7758 42393 7774
rect 42359 7366 42393 7382
rect 42473 7758 42507 7774
rect 42473 7366 42507 7382
rect 42731 7758 42765 7774
rect 42731 7366 42765 7382
rect 42845 7758 42879 7774
rect 42845 7366 42879 7382
rect 43103 7758 43137 7774
rect 43103 7366 43137 7382
rect 43217 7758 43251 7774
rect 43217 7366 43251 7382
rect 43475 7758 43509 7774
rect 43475 7366 43509 7382
rect 43589 7758 43623 7774
rect 43589 7366 43623 7382
rect 43847 7758 43881 7774
rect 43847 7366 43881 7382
rect 43961 7758 43995 7774
rect 43961 7366 43995 7382
rect 44219 7758 44253 7774
rect 44219 7366 44253 7382
rect 44333 7758 44367 7774
rect 44333 7366 44367 7382
rect 44591 7758 44625 7774
rect 44591 7366 44625 7382
rect 44705 7758 44739 7774
rect 44705 7366 44739 7382
rect 44963 7758 44997 7774
rect 44963 7366 44997 7382
rect 45077 7758 45111 7774
rect 45077 7366 45111 7382
rect 45335 7758 45369 7774
rect 45335 7366 45369 7382
rect 45449 7758 45483 7774
rect 45449 7366 45483 7382
rect 45707 7758 45741 7774
rect 45707 7366 45741 7382
rect 45821 7758 45855 7774
rect 45821 7366 45855 7382
rect 46079 7758 46113 7774
rect 46079 7366 46113 7382
rect 46193 7758 46227 7774
rect 46193 7366 46227 7382
rect 46451 7758 46485 7774
rect 46451 7366 46485 7382
rect 46565 7758 46599 7774
rect 46565 7366 46599 7382
rect 46823 7758 46857 7774
rect 46823 7366 46857 7382
rect 46937 7758 46971 7774
rect 46937 7366 46971 7382
rect 47195 7758 47229 7774
rect 47195 7366 47229 7382
rect 47309 7758 47343 7774
rect 47309 7366 47343 7382
rect 47567 7758 47601 7774
rect 47567 7366 47601 7382
rect 47681 7758 47715 7774
rect 47681 7366 47715 7382
rect 47939 7758 47973 7774
rect 47939 7366 47973 7382
rect 48053 7758 48087 7774
rect 48053 7366 48087 7382
rect 48311 7758 48345 7774
rect 48311 7366 48345 7382
rect 48425 7758 48459 7774
rect 48425 7366 48459 7382
rect 48683 7758 48717 7774
rect 48683 7366 48717 7382
rect 48797 7758 48831 7774
rect 48797 7366 48831 7382
rect 49055 7758 49089 7774
rect 49055 7366 49089 7382
rect 49169 7758 49203 7774
rect 49169 7366 49203 7382
rect 49427 7758 49461 7774
rect 49427 7366 49461 7382
rect 49541 7758 49575 7774
rect 49541 7366 49575 7382
rect 49799 7758 49833 7774
rect 49799 7366 49833 7382
rect 38055 7289 38071 7323
rect 38239 7289 38255 7323
rect 38427 7289 38443 7323
rect 38611 7289 38627 7323
rect 38799 7289 38815 7323
rect 38983 7289 38999 7323
rect 39171 7289 39187 7323
rect 39355 7289 39371 7323
rect 39543 7289 39559 7323
rect 39727 7289 39743 7323
rect 39915 7289 39931 7323
rect 40099 7289 40115 7323
rect 40287 7289 40303 7323
rect 40471 7289 40487 7323
rect 40659 7289 40675 7323
rect 40843 7289 40859 7323
rect 41031 7289 41047 7323
rect 41215 7289 41231 7323
rect 41403 7289 41419 7323
rect 41587 7289 41603 7323
rect 41775 7289 41791 7323
rect 41959 7289 41975 7323
rect 42147 7289 42163 7323
rect 42331 7289 42347 7323
rect 42519 7289 42535 7323
rect 42703 7289 42719 7323
rect 42891 7289 42907 7323
rect 43075 7289 43091 7323
rect 43263 7289 43279 7323
rect 43447 7289 43463 7323
rect 43635 7289 43651 7323
rect 43819 7289 43835 7323
rect 44007 7289 44023 7323
rect 44191 7289 44207 7323
rect 44379 7289 44395 7323
rect 44563 7289 44579 7323
rect 44751 7289 44767 7323
rect 44935 7289 44951 7323
rect 45123 7289 45139 7323
rect 45307 7289 45323 7323
rect 45495 7289 45511 7323
rect 45679 7289 45695 7323
rect 45867 7289 45883 7323
rect 46051 7289 46067 7323
rect 46239 7289 46255 7323
rect 46423 7289 46439 7323
rect 46611 7289 46627 7323
rect 46795 7289 46811 7323
rect 46983 7289 46999 7323
rect 47167 7289 47183 7323
rect 47355 7289 47371 7323
rect 47539 7289 47555 7323
rect 47727 7289 47743 7323
rect 47911 7289 47927 7323
rect 48099 7289 48115 7323
rect 48283 7289 48299 7323
rect 48471 7289 48487 7323
rect 48655 7289 48671 7323
rect 48843 7289 48859 7323
rect 49027 7289 49043 7323
rect 49215 7289 49231 7323
rect 49399 7289 49415 7323
rect 49587 7289 49603 7323
rect 49771 7289 49787 7323
rect 37895 7221 37929 7283
rect 49913 7221 49947 7283
rect 37895 7187 37991 7221
rect 49851 7187 49947 7221
rect 39383 6803 39468 6837
rect 42411 6803 42507 6837
rect 39383 6741 39417 6803
rect 42473 6741 42507 6803
rect 39543 6701 39559 6735
rect 39727 6701 39743 6735
rect 39915 6701 39931 6735
rect 40099 6701 40115 6735
rect 40287 6701 40303 6735
rect 40471 6701 40487 6735
rect 40659 6701 40675 6735
rect 40843 6701 40859 6735
rect 41031 6701 41047 6735
rect 41215 6701 41231 6735
rect 41403 6701 41419 6735
rect 41587 6701 41603 6735
rect 41775 6701 41791 6735
rect 41959 6701 41975 6735
rect 42147 6701 42163 6735
rect 42331 6701 42347 6735
rect 39497 6642 39531 6658
rect 39497 5850 39531 5866
rect 39755 6642 39789 6658
rect 39755 5850 39789 5866
rect 39869 6642 39903 6658
rect 39869 5850 39903 5866
rect 40127 6642 40161 6658
rect 40127 5850 40161 5866
rect 40241 6642 40275 6658
rect 40241 5850 40275 5866
rect 40499 6642 40533 6658
rect 40499 5850 40533 5866
rect 40613 6642 40647 6658
rect 40613 5850 40647 5866
rect 40871 6642 40905 6658
rect 40871 5850 40905 5866
rect 40985 6642 41019 6658
rect 40985 5850 41019 5866
rect 41243 6642 41277 6658
rect 41243 5850 41277 5866
rect 41357 6642 41391 6658
rect 41357 5850 41391 5866
rect 41615 6642 41649 6658
rect 41615 5850 41649 5866
rect 41729 6642 41763 6658
rect 41729 5850 41763 5866
rect 41987 6642 42021 6658
rect 41987 5850 42021 5866
rect 42101 6642 42135 6658
rect 42101 5850 42135 5866
rect 42359 6642 42393 6658
rect 42359 5850 42393 5866
rect 39543 5773 39559 5807
rect 39727 5773 39743 5807
rect 39915 5773 39931 5807
rect 40099 5773 40115 5807
rect 40287 5773 40303 5807
rect 40471 5773 40487 5807
rect 40659 5773 40675 5807
rect 40843 5773 40859 5807
rect 41031 5773 41047 5807
rect 41215 5773 41231 5807
rect 41403 5773 41419 5807
rect 41587 5773 41603 5807
rect 41775 5773 41791 5807
rect 41959 5773 41975 5807
rect 42147 5773 42163 5807
rect 42331 5773 42347 5807
rect 39543 5665 39559 5699
rect 39727 5665 39743 5699
rect 39915 5665 39931 5699
rect 40099 5665 40115 5699
rect 40287 5665 40303 5699
rect 40471 5665 40487 5699
rect 40659 5665 40675 5699
rect 40843 5665 40859 5699
rect 41031 5665 41047 5699
rect 41215 5665 41231 5699
rect 41403 5665 41419 5699
rect 41587 5665 41603 5699
rect 41775 5665 41791 5699
rect 41959 5665 41975 5699
rect 42147 5665 42163 5699
rect 42331 5665 42347 5699
rect 39497 5606 39531 5622
rect 39497 4814 39531 4830
rect 39755 5606 39789 5622
rect 39755 4814 39789 4830
rect 39869 5606 39903 5622
rect 39869 4814 39903 4830
rect 40127 5606 40161 5622
rect 40127 4814 40161 4830
rect 40241 5606 40275 5622
rect 40241 4814 40275 4830
rect 40499 5606 40533 5622
rect 40499 4814 40533 4830
rect 40613 5606 40647 5622
rect 40613 4814 40647 4830
rect 40871 5606 40905 5622
rect 40871 4814 40905 4830
rect 40985 5606 41019 5622
rect 40985 4814 41019 4830
rect 41243 5606 41277 5622
rect 41243 4814 41277 4830
rect 41357 5606 41391 5622
rect 41357 4814 41391 4830
rect 41615 5606 41649 5622
rect 41615 4814 41649 4830
rect 41729 5606 41763 5622
rect 41729 4814 41763 4830
rect 41987 5606 42021 5622
rect 41987 4814 42021 4830
rect 42101 5606 42135 5622
rect 42101 4814 42135 4830
rect 42359 5606 42393 5622
rect 42359 4814 42393 4830
rect 39543 4737 39559 4771
rect 39727 4737 39743 4771
rect 39915 4737 39931 4771
rect 40099 4737 40115 4771
rect 40287 4737 40303 4771
rect 40471 4737 40487 4771
rect 40659 4737 40675 4771
rect 40843 4737 40859 4771
rect 41031 4737 41047 4771
rect 41215 4737 41231 4771
rect 41403 4737 41419 4771
rect 41587 4737 41603 4771
rect 41775 4737 41791 4771
rect 41959 4737 41975 4771
rect 42147 4737 42163 4771
rect 42331 4737 42347 4771
rect 39543 4629 39559 4663
rect 39727 4629 39743 4663
rect 39915 4629 39931 4663
rect 40099 4629 40115 4663
rect 40287 4629 40303 4663
rect 40471 4629 40487 4663
rect 40659 4629 40675 4663
rect 40843 4629 40859 4663
rect 41031 4629 41047 4663
rect 41215 4629 41231 4663
rect 41403 4629 41419 4663
rect 41587 4629 41603 4663
rect 41775 4629 41791 4663
rect 41959 4629 41975 4663
rect 42147 4629 42163 4663
rect 42331 4629 42347 4663
rect 39497 4570 39531 4586
rect 39497 3778 39531 3794
rect 39755 4570 39789 4586
rect 39755 3778 39789 3794
rect 39869 4570 39903 4586
rect 39869 3778 39903 3794
rect 40127 4570 40161 4586
rect 40127 3778 40161 3794
rect 40241 4570 40275 4586
rect 40241 3778 40275 3794
rect 40499 4570 40533 4586
rect 40499 3778 40533 3794
rect 40613 4570 40647 4586
rect 40613 3778 40647 3794
rect 40871 4570 40905 4586
rect 40871 3778 40905 3794
rect 40985 4570 41019 4586
rect 40985 3778 41019 3794
rect 41243 4570 41277 4586
rect 41243 3778 41277 3794
rect 41357 4570 41391 4586
rect 41357 3778 41391 3794
rect 41615 4570 41649 4586
rect 41615 3778 41649 3794
rect 41729 4570 41763 4586
rect 41729 3778 41763 3794
rect 41987 4570 42021 4586
rect 41987 3778 42021 3794
rect 42101 4570 42135 4586
rect 42101 3778 42135 3794
rect 42359 4570 42393 4586
rect 42359 3778 42393 3794
rect 39543 3701 39559 3735
rect 39727 3701 39743 3735
rect 39915 3701 39931 3735
rect 40099 3701 40115 3735
rect 40287 3701 40303 3735
rect 40471 3701 40487 3735
rect 40659 3701 40675 3735
rect 40843 3701 40859 3735
rect 41031 3701 41047 3735
rect 41215 3701 41231 3735
rect 41403 3701 41419 3735
rect 41587 3701 41603 3735
rect 41775 3701 41791 3735
rect 41959 3701 41975 3735
rect 42147 3701 42163 3735
rect 42331 3701 42347 3735
rect 39543 3593 39559 3627
rect 39727 3593 39743 3627
rect 39915 3593 39931 3627
rect 40099 3593 40115 3627
rect 40287 3593 40303 3627
rect 40471 3593 40487 3627
rect 40659 3593 40675 3627
rect 40843 3593 40859 3627
rect 41031 3593 41047 3627
rect 41215 3593 41231 3627
rect 41403 3593 41419 3627
rect 41587 3593 41603 3627
rect 41775 3593 41791 3627
rect 41959 3593 41975 3627
rect 42147 3593 42163 3627
rect 42331 3593 42347 3627
rect 39497 3534 39531 3550
rect 39497 2742 39531 2758
rect 39755 3534 39789 3550
rect 39755 2742 39789 2758
rect 39869 3534 39903 3550
rect 39869 2742 39903 2758
rect 40127 3534 40161 3550
rect 40127 2742 40161 2758
rect 40241 3534 40275 3550
rect 40241 2742 40275 2758
rect 40499 3534 40533 3550
rect 40499 2742 40533 2758
rect 40613 3534 40647 3550
rect 40613 2742 40647 2758
rect 40871 3534 40905 3550
rect 40871 2742 40905 2758
rect 40985 3534 41019 3550
rect 40985 2742 41019 2758
rect 41243 3534 41277 3550
rect 41243 2742 41277 2758
rect 41357 3534 41391 3550
rect 41357 2742 41391 2758
rect 41615 3534 41649 3550
rect 41615 2742 41649 2758
rect 41729 3534 41763 3550
rect 41729 2742 41763 2758
rect 41987 3534 42021 3550
rect 41987 2742 42021 2758
rect 42101 3534 42135 3550
rect 42101 2742 42135 2758
rect 42359 3534 42393 3550
rect 42359 2742 42393 2758
rect 39543 2665 39559 2699
rect 39727 2665 39743 2699
rect 39915 2665 39931 2699
rect 40099 2665 40115 2699
rect 40287 2665 40303 2699
rect 40471 2665 40487 2699
rect 40659 2665 40675 2699
rect 40843 2665 40859 2699
rect 41031 2665 41047 2699
rect 41215 2665 41231 2699
rect 41403 2665 41419 2699
rect 41587 2665 41603 2699
rect 41775 2665 41791 2699
rect 41959 2665 41975 2699
rect 42147 2665 42163 2699
rect 42331 2665 42347 2699
rect 39383 2597 39417 2659
rect 43009 4889 43105 4923
rect 43243 4889 43339 4923
rect 43009 4827 43043 4889
rect 43305 4827 43339 4889
rect 43009 3273 43043 3335
rect 43305 3273 43339 3335
rect 43009 3239 43105 3273
rect 43243 3239 43339 3273
rect 42473 2597 42507 2659
rect 39383 2563 39479 2597
rect 42411 2563 42507 2597
rect 39383 2109 39479 2143
rect 48363 2109 48459 2143
rect 39383 2047 39417 2109
rect 48425 2047 48459 2109
rect 39543 2007 39559 2041
rect 39727 2007 39743 2041
rect 39915 2007 39931 2041
rect 40099 2007 40115 2041
rect 40287 2007 40303 2041
rect 40471 2007 40487 2041
rect 40659 2007 40675 2041
rect 40843 2007 40859 2041
rect 41031 2007 41047 2041
rect 41215 2007 41231 2041
rect 41403 2007 41419 2041
rect 41587 2007 41603 2041
rect 41775 2007 41791 2041
rect 41959 2007 41975 2041
rect 42147 2007 42163 2041
rect 42331 2007 42347 2041
rect 42519 2007 42535 2041
rect 42703 2007 42719 2041
rect 42891 2007 42907 2041
rect 43075 2007 43091 2041
rect 43263 2007 43279 2041
rect 43447 2007 43463 2041
rect 43635 2007 43651 2041
rect 43819 2007 43835 2041
rect 44007 2007 44023 2041
rect 44191 2007 44207 2041
rect 44379 2007 44395 2041
rect 44563 2007 44579 2041
rect 44751 2007 44767 2041
rect 44935 2007 44951 2041
rect 45123 2007 45139 2041
rect 45307 2007 45323 2041
rect 45495 2007 45511 2041
rect 45679 2007 45695 2041
rect 45867 2007 45883 2041
rect 46051 2007 46067 2041
rect 46239 2007 46255 2041
rect 46423 2007 46439 2041
rect 46611 2007 46627 2041
rect 46795 2007 46811 2041
rect 46983 2007 46999 2041
rect 47167 2007 47183 2041
rect 47355 2007 47371 2041
rect 47539 2007 47555 2041
rect 47727 2007 47743 2041
rect 47911 2007 47927 2041
rect 48099 2007 48115 2041
rect 48283 2007 48299 2041
rect 39497 1957 39531 1973
rect 39497 1765 39531 1781
rect 39755 1957 39789 1973
rect 39755 1765 39789 1781
rect 39869 1957 39903 1973
rect 39869 1765 39903 1781
rect 40127 1957 40161 1973
rect 40127 1765 40161 1781
rect 40241 1957 40275 1973
rect 40241 1765 40275 1781
rect 40499 1957 40533 1973
rect 40499 1765 40533 1781
rect 40613 1957 40647 1973
rect 40613 1765 40647 1781
rect 40871 1957 40905 1973
rect 40871 1765 40905 1781
rect 40985 1957 41019 1973
rect 40985 1765 41019 1781
rect 41243 1957 41277 1973
rect 41243 1765 41277 1781
rect 41357 1957 41391 1973
rect 41357 1765 41391 1781
rect 41615 1957 41649 1973
rect 41615 1765 41649 1781
rect 41729 1957 41763 1973
rect 41729 1765 41763 1781
rect 41987 1957 42021 1973
rect 41987 1765 42021 1781
rect 42101 1957 42135 1973
rect 42101 1765 42135 1781
rect 42359 1957 42393 1973
rect 42359 1765 42393 1781
rect 42473 1957 42507 1973
rect 42473 1765 42507 1781
rect 42731 1957 42765 1973
rect 42731 1765 42765 1781
rect 42845 1957 42879 1973
rect 42845 1765 42879 1781
rect 43103 1957 43137 1973
rect 43103 1765 43137 1781
rect 43217 1957 43251 1973
rect 43217 1765 43251 1781
rect 43475 1957 43509 1973
rect 43475 1765 43509 1781
rect 43589 1957 43623 1973
rect 43589 1765 43623 1781
rect 43847 1957 43881 1973
rect 43847 1765 43881 1781
rect 43961 1957 43995 1973
rect 43961 1765 43995 1781
rect 44219 1957 44253 1973
rect 44219 1765 44253 1781
rect 44333 1957 44367 1973
rect 44333 1765 44367 1781
rect 44591 1957 44625 1973
rect 44591 1765 44625 1781
rect 44705 1957 44739 1973
rect 44705 1765 44739 1781
rect 44963 1957 44997 1973
rect 44963 1765 44997 1781
rect 45077 1957 45111 1973
rect 45077 1765 45111 1781
rect 45335 1957 45369 1973
rect 45335 1765 45369 1781
rect 45449 1957 45483 1973
rect 45449 1765 45483 1781
rect 45707 1957 45741 1973
rect 45707 1765 45741 1781
rect 45821 1957 45855 1973
rect 45821 1765 45855 1781
rect 46079 1957 46113 1973
rect 46079 1765 46113 1781
rect 46193 1957 46227 1973
rect 46193 1765 46227 1781
rect 46451 1957 46485 1973
rect 46451 1765 46485 1781
rect 46565 1957 46599 1973
rect 46565 1765 46599 1781
rect 46823 1957 46857 1973
rect 46823 1765 46857 1781
rect 46937 1957 46971 1973
rect 46937 1765 46971 1781
rect 47195 1957 47229 1973
rect 47195 1765 47229 1781
rect 47309 1957 47343 1973
rect 47309 1765 47343 1781
rect 47567 1957 47601 1973
rect 47567 1765 47601 1781
rect 47681 1957 47715 1973
rect 47681 1765 47715 1781
rect 47939 1957 47973 1973
rect 47939 1765 47973 1781
rect 48053 1957 48087 1973
rect 48053 1765 48087 1781
rect 48311 1957 48345 1973
rect 48311 1765 48345 1781
rect 39543 1697 39559 1731
rect 39727 1697 39743 1731
rect 39915 1697 39931 1731
rect 40099 1697 40115 1731
rect 40287 1697 40303 1731
rect 40471 1697 40487 1731
rect 40659 1697 40675 1731
rect 40843 1697 40859 1731
rect 41031 1697 41047 1731
rect 41215 1697 41231 1731
rect 41403 1697 41419 1731
rect 41587 1697 41603 1731
rect 41775 1697 41791 1731
rect 41959 1697 41975 1731
rect 42147 1697 42163 1731
rect 42331 1697 42347 1731
rect 42519 1697 42535 1731
rect 42703 1697 42719 1731
rect 42891 1697 42907 1731
rect 43075 1697 43091 1731
rect 43263 1697 43279 1731
rect 43447 1697 43463 1731
rect 43635 1697 43651 1731
rect 43819 1697 43835 1731
rect 44007 1697 44023 1731
rect 44191 1697 44207 1731
rect 44379 1697 44395 1731
rect 44563 1697 44579 1731
rect 44751 1697 44767 1731
rect 44935 1697 44951 1731
rect 45123 1697 45139 1731
rect 45307 1697 45323 1731
rect 45495 1697 45511 1731
rect 45679 1697 45695 1731
rect 45867 1697 45883 1731
rect 46051 1697 46067 1731
rect 46239 1697 46255 1731
rect 46423 1697 46439 1731
rect 46611 1697 46627 1731
rect 46795 1697 46811 1731
rect 46983 1697 46999 1731
rect 47167 1697 47183 1731
rect 47355 1697 47371 1731
rect 47539 1697 47555 1731
rect 47727 1697 47743 1731
rect 47911 1697 47927 1731
rect 48099 1697 48115 1731
rect 48283 1697 48299 1731
rect 39543 1589 39559 1623
rect 39727 1589 39743 1623
rect 39915 1589 39931 1623
rect 40099 1589 40115 1623
rect 40287 1589 40303 1623
rect 40471 1589 40487 1623
rect 40659 1589 40675 1623
rect 40843 1589 40859 1623
rect 41031 1589 41047 1623
rect 41215 1589 41231 1623
rect 41403 1589 41419 1623
rect 41587 1589 41603 1623
rect 41775 1589 41791 1623
rect 41959 1589 41975 1623
rect 42147 1589 42163 1623
rect 42331 1589 42347 1623
rect 42519 1589 42535 1623
rect 42703 1589 42719 1623
rect 42891 1589 42907 1623
rect 43075 1589 43091 1623
rect 43263 1589 43279 1623
rect 43447 1589 43463 1623
rect 43635 1589 43651 1623
rect 43819 1589 43835 1623
rect 44007 1589 44023 1623
rect 44191 1589 44207 1623
rect 44379 1589 44395 1623
rect 44563 1589 44579 1623
rect 44751 1589 44767 1623
rect 44935 1589 44951 1623
rect 45123 1589 45139 1623
rect 45307 1589 45323 1623
rect 45495 1589 45511 1623
rect 45679 1589 45695 1623
rect 45867 1589 45883 1623
rect 46051 1589 46067 1623
rect 46239 1589 46255 1623
rect 46423 1589 46439 1623
rect 46611 1589 46627 1623
rect 46795 1589 46811 1623
rect 46983 1589 46999 1623
rect 47167 1589 47183 1623
rect 47355 1589 47371 1623
rect 47539 1589 47555 1623
rect 47727 1589 47743 1623
rect 47911 1589 47927 1623
rect 48099 1589 48115 1623
rect 48283 1589 48299 1623
rect 39497 1539 39531 1555
rect 39497 1347 39531 1363
rect 39755 1539 39789 1555
rect 39755 1347 39789 1363
rect 39869 1539 39903 1555
rect 39869 1347 39903 1363
rect 40127 1539 40161 1555
rect 40127 1347 40161 1363
rect 40241 1539 40275 1555
rect 40241 1347 40275 1363
rect 40499 1539 40533 1555
rect 40499 1347 40533 1363
rect 40613 1539 40647 1555
rect 40613 1347 40647 1363
rect 40871 1539 40905 1555
rect 40871 1347 40905 1363
rect 40985 1539 41019 1555
rect 40985 1347 41019 1363
rect 41243 1539 41277 1555
rect 41243 1347 41277 1363
rect 41357 1539 41391 1555
rect 41357 1347 41391 1363
rect 41615 1539 41649 1555
rect 41615 1347 41649 1363
rect 41729 1539 41763 1555
rect 41729 1347 41763 1363
rect 41987 1539 42021 1555
rect 41987 1347 42021 1363
rect 42101 1539 42135 1555
rect 42101 1347 42135 1363
rect 42359 1539 42393 1555
rect 42359 1347 42393 1363
rect 42473 1539 42507 1555
rect 42473 1347 42507 1363
rect 42731 1539 42765 1555
rect 42731 1347 42765 1363
rect 42845 1539 42879 1555
rect 42845 1347 42879 1363
rect 43103 1539 43137 1555
rect 43103 1347 43137 1363
rect 43217 1539 43251 1555
rect 43217 1347 43251 1363
rect 43475 1539 43509 1555
rect 43475 1347 43509 1363
rect 43589 1539 43623 1555
rect 43589 1347 43623 1363
rect 43847 1539 43881 1555
rect 43847 1347 43881 1363
rect 43961 1539 43995 1555
rect 43961 1347 43995 1363
rect 44219 1539 44253 1555
rect 44219 1347 44253 1363
rect 44333 1539 44367 1555
rect 44333 1347 44367 1363
rect 44591 1539 44625 1555
rect 44591 1347 44625 1363
rect 44705 1539 44739 1555
rect 44705 1347 44739 1363
rect 44963 1539 44997 1555
rect 44963 1347 44997 1363
rect 45077 1539 45111 1555
rect 45077 1347 45111 1363
rect 45335 1539 45369 1555
rect 45335 1347 45369 1363
rect 45449 1539 45483 1555
rect 45449 1347 45483 1363
rect 45707 1539 45741 1555
rect 45707 1347 45741 1363
rect 45821 1539 45855 1555
rect 45821 1347 45855 1363
rect 46079 1539 46113 1555
rect 46079 1347 46113 1363
rect 46193 1539 46227 1555
rect 46193 1347 46227 1363
rect 46451 1539 46485 1555
rect 46451 1347 46485 1363
rect 46565 1539 46599 1555
rect 46565 1347 46599 1363
rect 46823 1539 46857 1555
rect 46823 1347 46857 1363
rect 46937 1539 46971 1555
rect 46937 1347 46971 1363
rect 47195 1539 47229 1555
rect 47195 1347 47229 1363
rect 47309 1539 47343 1555
rect 47309 1347 47343 1363
rect 47567 1539 47601 1555
rect 47567 1347 47601 1363
rect 47681 1539 47715 1555
rect 47681 1347 47715 1363
rect 47939 1539 47973 1555
rect 47939 1347 47973 1363
rect 48053 1539 48087 1555
rect 48053 1347 48087 1363
rect 48311 1539 48345 1555
rect 48311 1347 48345 1363
rect 39543 1279 39559 1313
rect 39727 1279 39743 1313
rect 39915 1279 39931 1313
rect 40099 1279 40115 1313
rect 40287 1279 40303 1313
rect 40471 1279 40487 1313
rect 40659 1279 40675 1313
rect 40843 1279 40859 1313
rect 41031 1279 41047 1313
rect 41215 1279 41231 1313
rect 41403 1279 41419 1313
rect 41587 1279 41603 1313
rect 41775 1279 41791 1313
rect 41959 1279 41975 1313
rect 42147 1279 42163 1313
rect 42331 1279 42347 1313
rect 42519 1279 42535 1313
rect 42703 1279 42719 1313
rect 42891 1279 42907 1313
rect 43075 1279 43091 1313
rect 43263 1279 43279 1313
rect 43447 1279 43463 1313
rect 43635 1279 43651 1313
rect 43819 1279 43835 1313
rect 44007 1279 44023 1313
rect 44191 1279 44207 1313
rect 44379 1279 44395 1313
rect 44563 1279 44579 1313
rect 44751 1279 44767 1313
rect 44935 1279 44951 1313
rect 45123 1279 45139 1313
rect 45307 1279 45323 1313
rect 45495 1279 45511 1313
rect 45679 1279 45695 1313
rect 45867 1279 45883 1313
rect 46051 1279 46067 1313
rect 46239 1279 46255 1313
rect 46423 1279 46439 1313
rect 46611 1279 46627 1313
rect 46795 1279 46811 1313
rect 46983 1279 46999 1313
rect 47167 1279 47183 1313
rect 47355 1279 47371 1313
rect 47539 1279 47555 1313
rect 47727 1279 47743 1313
rect 47911 1279 47927 1313
rect 48099 1279 48115 1313
rect 48283 1279 48299 1313
rect 39543 1171 39559 1205
rect 39727 1171 39743 1205
rect 39915 1171 39931 1205
rect 40099 1171 40115 1205
rect 40287 1171 40303 1205
rect 40471 1171 40487 1205
rect 40659 1171 40675 1205
rect 40843 1171 40859 1205
rect 41031 1171 41047 1205
rect 41215 1171 41231 1205
rect 41403 1171 41419 1205
rect 41587 1171 41603 1205
rect 41775 1171 41791 1205
rect 41959 1171 41975 1205
rect 42147 1171 42163 1205
rect 42331 1171 42347 1205
rect 42519 1171 42535 1205
rect 42703 1171 42719 1205
rect 42891 1171 42907 1205
rect 43075 1171 43091 1205
rect 43263 1171 43279 1205
rect 43447 1171 43463 1205
rect 43635 1171 43651 1205
rect 43819 1171 43835 1205
rect 44007 1171 44023 1205
rect 44191 1171 44207 1205
rect 44379 1171 44395 1205
rect 44563 1171 44579 1205
rect 44751 1171 44767 1205
rect 44935 1171 44951 1205
rect 45123 1171 45139 1205
rect 45307 1171 45323 1205
rect 45495 1171 45511 1205
rect 45679 1171 45695 1205
rect 45867 1171 45883 1205
rect 46051 1171 46067 1205
rect 46239 1171 46255 1205
rect 46423 1171 46439 1205
rect 46611 1171 46627 1205
rect 46795 1171 46811 1205
rect 46983 1171 46999 1205
rect 47167 1171 47183 1205
rect 47355 1171 47371 1205
rect 47539 1171 47555 1205
rect 47727 1171 47743 1205
rect 47911 1171 47927 1205
rect 48099 1171 48115 1205
rect 48283 1171 48299 1205
rect 39497 1121 39531 1137
rect 39497 929 39531 945
rect 39755 1121 39789 1137
rect 39755 929 39789 945
rect 39869 1121 39903 1137
rect 39869 929 39903 945
rect 40127 1121 40161 1137
rect 40127 929 40161 945
rect 40241 1121 40275 1137
rect 40241 929 40275 945
rect 40499 1121 40533 1137
rect 40499 929 40533 945
rect 40613 1121 40647 1137
rect 40613 929 40647 945
rect 40871 1121 40905 1137
rect 40871 929 40905 945
rect 40985 1121 41019 1137
rect 40985 929 41019 945
rect 41243 1121 41277 1137
rect 41243 929 41277 945
rect 41357 1121 41391 1137
rect 41357 929 41391 945
rect 41615 1121 41649 1137
rect 41615 929 41649 945
rect 41729 1121 41763 1137
rect 41729 929 41763 945
rect 41987 1121 42021 1137
rect 41987 929 42021 945
rect 42101 1121 42135 1137
rect 42101 929 42135 945
rect 42359 1121 42393 1137
rect 42359 929 42393 945
rect 42473 1121 42507 1137
rect 42473 929 42507 945
rect 42731 1121 42765 1137
rect 42731 929 42765 945
rect 42845 1121 42879 1137
rect 42845 929 42879 945
rect 43103 1121 43137 1137
rect 43103 929 43137 945
rect 43217 1121 43251 1137
rect 43217 929 43251 945
rect 43475 1121 43509 1137
rect 43475 929 43509 945
rect 43589 1121 43623 1137
rect 43589 929 43623 945
rect 43847 1121 43881 1137
rect 43847 929 43881 945
rect 43961 1121 43995 1137
rect 43961 929 43995 945
rect 44219 1121 44253 1137
rect 44219 929 44253 945
rect 44333 1121 44367 1137
rect 44333 929 44367 945
rect 44591 1121 44625 1137
rect 44591 929 44625 945
rect 44705 1121 44739 1137
rect 44705 929 44739 945
rect 44963 1121 44997 1137
rect 44963 929 44997 945
rect 45077 1121 45111 1137
rect 45077 929 45111 945
rect 45335 1121 45369 1137
rect 45335 929 45369 945
rect 45449 1121 45483 1137
rect 45449 929 45483 945
rect 45707 1121 45741 1137
rect 45707 929 45741 945
rect 45821 1121 45855 1137
rect 45821 929 45855 945
rect 46079 1121 46113 1137
rect 46079 929 46113 945
rect 46193 1121 46227 1137
rect 46193 929 46227 945
rect 46451 1121 46485 1137
rect 46451 929 46485 945
rect 46565 1121 46599 1137
rect 46565 929 46599 945
rect 46823 1121 46857 1137
rect 46823 929 46857 945
rect 46937 1121 46971 1137
rect 46937 929 46971 945
rect 47195 1121 47229 1137
rect 47195 929 47229 945
rect 47309 1121 47343 1137
rect 47309 929 47343 945
rect 47567 1121 47601 1137
rect 47567 929 47601 945
rect 47681 1121 47715 1137
rect 47681 929 47715 945
rect 47939 1121 47973 1137
rect 47939 929 47973 945
rect 48053 1121 48087 1137
rect 48053 929 48087 945
rect 48311 1121 48345 1137
rect 48311 929 48345 945
rect 39543 861 39559 895
rect 39727 861 39743 895
rect 39915 861 39931 895
rect 40099 861 40115 895
rect 40287 861 40303 895
rect 40471 861 40487 895
rect 40659 861 40675 895
rect 40843 861 40859 895
rect 41031 861 41047 895
rect 41215 861 41231 895
rect 41403 861 41419 895
rect 41587 861 41603 895
rect 41775 861 41791 895
rect 41959 861 41975 895
rect 42147 861 42163 895
rect 42331 861 42347 895
rect 42519 861 42535 895
rect 42703 861 42719 895
rect 42891 861 42907 895
rect 43075 861 43091 895
rect 43263 861 43279 895
rect 43447 861 43463 895
rect 43635 861 43651 895
rect 43819 861 43835 895
rect 44007 861 44023 895
rect 44191 861 44207 895
rect 44379 861 44395 895
rect 44563 861 44579 895
rect 44751 861 44767 895
rect 44935 861 44951 895
rect 45123 861 45139 895
rect 45307 861 45323 895
rect 45495 861 45511 895
rect 45679 861 45695 895
rect 45867 861 45883 895
rect 46051 861 46067 895
rect 46239 861 46255 895
rect 46423 861 46439 895
rect 46611 861 46627 895
rect 46795 861 46811 895
rect 46983 861 46999 895
rect 47167 861 47183 895
rect 47355 861 47371 895
rect 47539 861 47555 895
rect 47727 861 47743 895
rect 47911 861 47927 895
rect 48099 861 48115 895
rect 48283 861 48299 895
rect 39543 753 39559 787
rect 39727 753 39743 787
rect 39915 753 39931 787
rect 40099 753 40115 787
rect 40287 753 40303 787
rect 40471 753 40487 787
rect 40659 753 40675 787
rect 40843 753 40859 787
rect 41031 753 41047 787
rect 41215 753 41231 787
rect 41403 753 41419 787
rect 41587 753 41603 787
rect 41775 753 41791 787
rect 41959 753 41975 787
rect 42147 753 42163 787
rect 42331 753 42347 787
rect 42519 753 42535 787
rect 42703 753 42719 787
rect 42891 753 42907 787
rect 43075 753 43091 787
rect 43263 753 43279 787
rect 43447 753 43463 787
rect 43635 753 43651 787
rect 43819 753 43835 787
rect 44007 753 44023 787
rect 44191 753 44207 787
rect 44379 753 44395 787
rect 44563 753 44579 787
rect 44751 753 44767 787
rect 44935 753 44951 787
rect 45123 753 45139 787
rect 45307 753 45323 787
rect 45495 753 45511 787
rect 45679 753 45695 787
rect 45867 753 45883 787
rect 46051 753 46067 787
rect 46239 753 46255 787
rect 46423 753 46439 787
rect 46611 753 46627 787
rect 46795 753 46811 787
rect 46983 753 46999 787
rect 47167 753 47183 787
rect 47355 753 47371 787
rect 47539 753 47555 787
rect 47727 753 47743 787
rect 47911 753 47927 787
rect 48099 753 48115 787
rect 48283 753 48299 787
rect 39497 703 39531 719
rect 39497 511 39531 527
rect 39755 703 39789 719
rect 39755 511 39789 527
rect 39869 703 39903 719
rect 39869 511 39903 527
rect 40127 703 40161 719
rect 40127 511 40161 527
rect 40241 703 40275 719
rect 40241 511 40275 527
rect 40499 703 40533 719
rect 40499 511 40533 527
rect 40613 703 40647 719
rect 40613 511 40647 527
rect 40871 703 40905 719
rect 40871 511 40905 527
rect 40985 703 41019 719
rect 40985 511 41019 527
rect 41243 703 41277 719
rect 41243 511 41277 527
rect 41357 703 41391 719
rect 41357 511 41391 527
rect 41615 703 41649 719
rect 41615 511 41649 527
rect 41729 703 41763 719
rect 41729 511 41763 527
rect 41987 703 42021 719
rect 41987 511 42021 527
rect 42101 703 42135 719
rect 42101 511 42135 527
rect 42359 703 42393 719
rect 42359 511 42393 527
rect 42473 703 42507 719
rect 42473 511 42507 527
rect 42731 703 42765 719
rect 42731 511 42765 527
rect 42845 703 42879 719
rect 42845 511 42879 527
rect 43103 703 43137 719
rect 43103 511 43137 527
rect 43217 703 43251 719
rect 43217 511 43251 527
rect 43475 703 43509 719
rect 43475 511 43509 527
rect 43589 703 43623 719
rect 43589 511 43623 527
rect 43847 703 43881 719
rect 43847 511 43881 527
rect 43961 703 43995 719
rect 43961 511 43995 527
rect 44219 703 44253 719
rect 44219 511 44253 527
rect 44333 703 44367 719
rect 44333 511 44367 527
rect 44591 703 44625 719
rect 44591 511 44625 527
rect 44705 703 44739 719
rect 44705 511 44739 527
rect 44963 703 44997 719
rect 44963 511 44997 527
rect 45077 703 45111 719
rect 45077 511 45111 527
rect 45335 703 45369 719
rect 45335 511 45369 527
rect 45449 703 45483 719
rect 45449 511 45483 527
rect 45707 703 45741 719
rect 45707 511 45741 527
rect 45821 703 45855 719
rect 45821 511 45855 527
rect 46079 703 46113 719
rect 46079 511 46113 527
rect 46193 703 46227 719
rect 46193 511 46227 527
rect 46451 703 46485 719
rect 46451 511 46485 527
rect 46565 703 46599 719
rect 46565 511 46599 527
rect 46823 703 46857 719
rect 46823 511 46857 527
rect 46937 703 46971 719
rect 46937 511 46971 527
rect 47195 703 47229 719
rect 47195 511 47229 527
rect 47309 703 47343 719
rect 47309 511 47343 527
rect 47567 703 47601 719
rect 47567 511 47601 527
rect 47681 703 47715 719
rect 47681 511 47715 527
rect 47939 703 47973 719
rect 47939 511 47973 527
rect 48053 703 48087 719
rect 48053 511 48087 527
rect 48311 703 48345 719
rect 48311 511 48345 527
rect 39543 443 39559 477
rect 39727 443 39743 477
rect 39915 443 39931 477
rect 40099 443 40115 477
rect 40287 443 40303 477
rect 40471 443 40487 477
rect 40659 443 40675 477
rect 40843 443 40859 477
rect 41031 443 41047 477
rect 41215 443 41231 477
rect 41403 443 41419 477
rect 41587 443 41603 477
rect 41775 443 41791 477
rect 41959 443 41975 477
rect 42147 443 42163 477
rect 42331 443 42347 477
rect 42519 443 42535 477
rect 42703 443 42719 477
rect 42891 443 42907 477
rect 43075 443 43091 477
rect 43263 443 43279 477
rect 43447 443 43463 477
rect 43635 443 43651 477
rect 43819 443 43835 477
rect 44007 443 44023 477
rect 44191 443 44207 477
rect 44379 443 44395 477
rect 44563 443 44579 477
rect 44751 443 44767 477
rect 44935 443 44951 477
rect 45123 443 45139 477
rect 45307 443 45323 477
rect 45495 443 45511 477
rect 45679 443 45695 477
rect 45867 443 45883 477
rect 46051 443 46067 477
rect 46239 443 46255 477
rect 46423 443 46439 477
rect 46611 443 46627 477
rect 46795 443 46811 477
rect 46983 443 46999 477
rect 47167 443 47183 477
rect 47355 443 47371 477
rect 47539 443 47555 477
rect 47727 443 47743 477
rect 47911 443 47927 477
rect 48099 443 48115 477
rect 48283 443 48299 477
rect 39383 375 39417 437
rect 48425 375 48459 437
rect 39383 341 39479 375
rect 48363 341 48459 375
<< viali >>
rect 38306 9225 38376 9242
rect 39050 9225 39120 9242
rect 39794 9225 39864 9242
rect 40538 9225 40608 9242
rect 41282 9225 41352 9242
rect 42026 9225 42096 9242
rect 42770 9225 42840 9242
rect 43514 9225 43584 9242
rect 43886 9225 43956 9242
rect 44630 9225 44700 9242
rect 45374 9225 45444 9242
rect 46118 9225 46188 9242
rect 46862 9225 46932 9242
rect 47606 9225 47676 9242
rect 48350 9225 48420 9242
rect 49094 9225 49164 9242
rect 49784 9225 49854 9242
rect 38306 9191 38376 9225
rect 39050 9191 39120 9225
rect 39794 9191 39864 9225
rect 40538 9191 40608 9225
rect 41282 9191 41352 9225
rect 42026 9191 42096 9225
rect 42770 9191 42840 9225
rect 43514 9191 43584 9225
rect 43886 9191 43956 9225
rect 44630 9191 44700 9225
rect 45374 9191 45444 9225
rect 46118 9191 46188 9225
rect 46862 9191 46932 9225
rect 47606 9191 47676 9225
rect 48350 9191 48420 9225
rect 49094 9191 49164 9225
rect 49784 9191 49851 9225
rect 49851 9191 49854 9225
rect 38306 9172 38376 9191
rect 39050 9172 39120 9191
rect 39794 9172 39864 9191
rect 40538 9172 40608 9191
rect 41282 9172 41352 9191
rect 42026 9172 42096 9191
rect 42770 9172 42840 9191
rect 43514 9172 43584 9191
rect 43886 9172 43956 9191
rect 44630 9172 44700 9191
rect 45374 9172 45444 9191
rect 46118 9172 46188 9191
rect 46862 9172 46932 9191
rect 47606 9172 47676 9191
rect 48350 9172 48420 9191
rect 49094 9172 49164 9191
rect 49784 9172 49854 9191
rect 38071 9089 38239 9123
rect 38443 9089 38611 9123
rect 38815 9089 38983 9123
rect 39187 9089 39355 9123
rect 39559 9089 39727 9123
rect 39931 9089 40099 9123
rect 40303 9089 40471 9123
rect 40675 9089 40843 9123
rect 41047 9089 41215 9123
rect 41419 9089 41587 9123
rect 41791 9089 41959 9123
rect 42163 9089 42331 9123
rect 42535 9089 42703 9123
rect 42907 9089 43075 9123
rect 43279 9089 43447 9123
rect 43651 9089 43819 9123
rect 44023 9089 44191 9123
rect 44395 9089 44563 9123
rect 44767 9089 44935 9123
rect 45139 9089 45307 9123
rect 45511 9089 45679 9123
rect 45883 9089 46051 9123
rect 46255 9089 46423 9123
rect 46627 9089 46795 9123
rect 46999 9089 47167 9123
rect 47371 9089 47539 9123
rect 47743 9089 47911 9123
rect 48115 9089 48283 9123
rect 48487 9089 48655 9123
rect 48859 9089 49027 9123
rect 49231 9089 49399 9123
rect 49603 9089 49771 9123
rect 38009 8654 38043 9030
rect 38267 8654 38301 9030
rect 38381 8654 38415 9030
rect 38639 8654 38673 9030
rect 38753 8654 38787 9030
rect 39011 8654 39045 9030
rect 39125 8654 39159 9030
rect 39383 8654 39417 9030
rect 39497 8654 39531 9030
rect 39755 8654 39789 9030
rect 39869 8654 39903 9030
rect 40127 8654 40161 9030
rect 40241 8654 40275 9030
rect 40499 8654 40533 9030
rect 40613 8654 40647 9030
rect 40871 8654 40905 9030
rect 40985 8654 41019 9030
rect 41243 8654 41277 9030
rect 41357 8654 41391 9030
rect 41615 8654 41649 9030
rect 41729 8654 41763 9030
rect 41987 8654 42021 9030
rect 42101 8654 42135 9030
rect 42359 8654 42393 9030
rect 42473 8654 42507 9030
rect 42731 8654 42765 9030
rect 42845 8654 42879 9030
rect 43103 8654 43137 9030
rect 43217 8654 43251 9030
rect 43475 8654 43509 9030
rect 43589 8654 43623 9030
rect 43847 8654 43881 9030
rect 43961 8654 43995 9030
rect 44219 8654 44253 9030
rect 44333 8654 44367 9030
rect 44591 8654 44625 9030
rect 44705 8654 44739 9030
rect 44963 8654 44997 9030
rect 45077 8654 45111 9030
rect 45335 8654 45369 9030
rect 45449 8654 45483 9030
rect 45707 8654 45741 9030
rect 45821 8654 45855 9030
rect 46079 8654 46113 9030
rect 46193 8654 46227 9030
rect 46451 8654 46485 9030
rect 46565 8654 46599 9030
rect 46823 8654 46857 9030
rect 46937 8654 46971 9030
rect 47195 8654 47229 9030
rect 47309 8654 47343 9030
rect 47567 8654 47601 9030
rect 47681 8654 47715 9030
rect 47939 8654 47973 9030
rect 48053 8654 48087 9030
rect 48311 8654 48345 9030
rect 48425 8654 48459 9030
rect 48683 8654 48717 9030
rect 48797 8654 48831 9030
rect 49055 8654 49089 9030
rect 49169 8654 49203 9030
rect 49427 8654 49461 9030
rect 49541 8654 49575 9030
rect 49799 8654 49833 9030
rect 38071 8561 38239 8595
rect 38443 8561 38611 8595
rect 38815 8561 38983 8595
rect 39187 8561 39355 8595
rect 39559 8561 39727 8595
rect 39931 8561 40099 8595
rect 40303 8561 40471 8595
rect 40675 8561 40843 8595
rect 41047 8561 41215 8595
rect 41419 8561 41587 8595
rect 41791 8561 41959 8595
rect 42163 8561 42331 8595
rect 42535 8561 42703 8595
rect 42907 8561 43075 8595
rect 43279 8561 43447 8595
rect 43651 8561 43819 8595
rect 44023 8561 44191 8595
rect 44395 8561 44563 8595
rect 44767 8561 44935 8595
rect 45139 8561 45307 8595
rect 45511 8561 45679 8595
rect 45883 8561 46051 8595
rect 46255 8561 46423 8595
rect 46627 8561 46795 8595
rect 46999 8561 47167 8595
rect 47371 8561 47539 8595
rect 47743 8561 47911 8595
rect 48115 8561 48283 8595
rect 48487 8561 48655 8595
rect 48859 8561 49027 8595
rect 49231 8561 49399 8595
rect 49603 8561 49771 8595
rect 38071 8453 38239 8487
rect 38443 8453 38611 8487
rect 38815 8453 38983 8487
rect 39187 8453 39355 8487
rect 39559 8453 39727 8487
rect 39931 8453 40099 8487
rect 40303 8453 40471 8487
rect 40675 8453 40843 8487
rect 41047 8453 41215 8487
rect 41419 8453 41587 8487
rect 41791 8453 41959 8487
rect 42163 8453 42331 8487
rect 42535 8453 42703 8487
rect 42907 8453 43075 8487
rect 43279 8453 43447 8487
rect 43651 8453 43819 8487
rect 44023 8453 44191 8487
rect 44395 8453 44563 8487
rect 44767 8453 44935 8487
rect 45139 8453 45307 8487
rect 45511 8453 45679 8487
rect 45883 8453 46051 8487
rect 46255 8453 46423 8487
rect 46627 8453 46795 8487
rect 46999 8453 47167 8487
rect 47371 8453 47539 8487
rect 47743 8453 47911 8487
rect 48115 8453 48283 8487
rect 48487 8453 48655 8487
rect 48859 8453 49027 8487
rect 49231 8453 49399 8487
rect 49603 8453 49771 8487
rect 38009 8018 38043 8394
rect 38267 8018 38301 8394
rect 38381 8018 38415 8394
rect 38639 8018 38673 8394
rect 38753 8018 38787 8394
rect 39011 8018 39045 8394
rect 39125 8018 39159 8394
rect 39383 8018 39417 8394
rect 39497 8018 39531 8394
rect 39755 8018 39789 8394
rect 39869 8018 39903 8394
rect 40127 8018 40161 8394
rect 40241 8018 40275 8394
rect 40499 8018 40533 8394
rect 40613 8018 40647 8394
rect 40871 8018 40905 8394
rect 40985 8018 41019 8394
rect 41243 8018 41277 8394
rect 41357 8018 41391 8394
rect 41615 8018 41649 8394
rect 41729 8018 41763 8394
rect 41987 8018 42021 8394
rect 42101 8018 42135 8394
rect 42359 8018 42393 8394
rect 42473 8018 42507 8394
rect 42731 8018 42765 8394
rect 42845 8018 42879 8394
rect 43103 8018 43137 8394
rect 43217 8018 43251 8394
rect 43475 8018 43509 8394
rect 43589 8018 43623 8394
rect 43847 8018 43881 8394
rect 43961 8018 43995 8394
rect 44219 8018 44253 8394
rect 44333 8018 44367 8394
rect 44591 8018 44625 8394
rect 44705 8018 44739 8394
rect 44963 8018 44997 8394
rect 45077 8018 45111 8394
rect 45335 8018 45369 8394
rect 45449 8018 45483 8394
rect 45707 8018 45741 8394
rect 45821 8018 45855 8394
rect 46079 8018 46113 8394
rect 46193 8018 46227 8394
rect 46451 8018 46485 8394
rect 46565 8018 46599 8394
rect 46823 8018 46857 8394
rect 46937 8018 46971 8394
rect 47195 8018 47229 8394
rect 47309 8018 47343 8394
rect 47567 8018 47601 8394
rect 47681 8018 47715 8394
rect 47939 8018 47973 8394
rect 48053 8018 48087 8394
rect 48311 8018 48345 8394
rect 48425 8018 48459 8394
rect 48683 8018 48717 8394
rect 48797 8018 48831 8394
rect 49055 8018 49089 8394
rect 49169 8018 49203 8394
rect 49427 8018 49461 8394
rect 49541 8018 49575 8394
rect 49799 8018 49833 8394
rect 38071 7925 38239 7959
rect 38443 7925 38611 7959
rect 38815 7925 38983 7959
rect 39187 7925 39355 7959
rect 39559 7925 39727 7959
rect 39931 7925 40099 7959
rect 40303 7925 40471 7959
rect 40675 7925 40843 7959
rect 41047 7925 41215 7959
rect 41419 7925 41587 7959
rect 41791 7925 41959 7959
rect 42163 7925 42331 7959
rect 42535 7925 42703 7959
rect 42907 7925 43075 7959
rect 43279 7925 43447 7959
rect 43651 7925 43819 7959
rect 44023 7925 44191 7959
rect 44395 7925 44563 7959
rect 44767 7925 44935 7959
rect 45139 7925 45307 7959
rect 45511 7925 45679 7959
rect 45883 7925 46051 7959
rect 46255 7925 46423 7959
rect 46627 7925 46795 7959
rect 46999 7925 47167 7959
rect 47371 7925 47539 7959
rect 47743 7925 47911 7959
rect 48115 7925 48283 7959
rect 48487 7925 48655 7959
rect 48859 7925 49027 7959
rect 49231 7925 49399 7959
rect 49603 7925 49771 7959
rect 38071 7817 38239 7851
rect 38443 7817 38611 7851
rect 38815 7817 38983 7851
rect 39187 7817 39355 7851
rect 39559 7817 39727 7851
rect 39931 7817 40099 7851
rect 40303 7817 40471 7851
rect 40675 7817 40843 7851
rect 41047 7817 41215 7851
rect 41419 7817 41587 7851
rect 41791 7817 41959 7851
rect 42163 7817 42331 7851
rect 42535 7817 42703 7851
rect 42907 7817 43075 7851
rect 43279 7817 43447 7851
rect 43651 7817 43819 7851
rect 44023 7817 44191 7851
rect 44395 7817 44563 7851
rect 44767 7817 44935 7851
rect 45139 7817 45307 7851
rect 45511 7817 45679 7851
rect 45883 7817 46051 7851
rect 46255 7817 46423 7851
rect 46627 7817 46795 7851
rect 46999 7817 47167 7851
rect 47371 7817 47539 7851
rect 47743 7817 47911 7851
rect 48115 7817 48283 7851
rect 48487 7817 48655 7851
rect 48859 7817 49027 7851
rect 49231 7817 49399 7851
rect 49603 7817 49771 7851
rect 38009 7382 38043 7758
rect 38267 7382 38301 7758
rect 38381 7382 38415 7758
rect 38639 7382 38673 7758
rect 38753 7382 38787 7758
rect 39011 7382 39045 7758
rect 39125 7382 39159 7758
rect 39383 7382 39417 7758
rect 39497 7382 39531 7758
rect 39755 7382 39789 7758
rect 39869 7382 39903 7758
rect 40127 7382 40161 7758
rect 40241 7382 40275 7758
rect 40499 7382 40533 7758
rect 40613 7382 40647 7758
rect 40871 7382 40905 7758
rect 40985 7382 41019 7758
rect 41243 7382 41277 7758
rect 41357 7382 41391 7758
rect 41615 7382 41649 7758
rect 41729 7382 41763 7758
rect 41987 7382 42021 7758
rect 42101 7382 42135 7758
rect 42359 7382 42393 7758
rect 42473 7382 42507 7758
rect 42731 7382 42765 7758
rect 42845 7382 42879 7758
rect 43103 7382 43137 7758
rect 43217 7382 43251 7758
rect 43475 7382 43509 7758
rect 43589 7382 43623 7758
rect 43847 7382 43881 7758
rect 43961 7382 43995 7758
rect 44219 7382 44253 7758
rect 44333 7382 44367 7758
rect 44591 7382 44625 7758
rect 44705 7382 44739 7758
rect 44963 7382 44997 7758
rect 45077 7382 45111 7758
rect 45335 7382 45369 7758
rect 45449 7382 45483 7758
rect 45707 7382 45741 7758
rect 45821 7382 45855 7758
rect 46079 7382 46113 7758
rect 46193 7382 46227 7758
rect 46451 7382 46485 7758
rect 46565 7382 46599 7758
rect 46823 7382 46857 7758
rect 46937 7382 46971 7758
rect 47195 7382 47229 7758
rect 47309 7382 47343 7758
rect 47567 7382 47601 7758
rect 47681 7382 47715 7758
rect 47939 7382 47973 7758
rect 48053 7382 48087 7758
rect 48311 7382 48345 7758
rect 48425 7382 48459 7758
rect 48683 7382 48717 7758
rect 48797 7382 48831 7758
rect 49055 7382 49089 7758
rect 49169 7382 49203 7758
rect 49427 7382 49461 7758
rect 49541 7382 49575 7758
rect 49799 7382 49833 7758
rect 38071 7289 38239 7323
rect 38443 7289 38611 7323
rect 38815 7289 38983 7323
rect 39187 7289 39355 7323
rect 39559 7289 39727 7323
rect 39931 7289 40099 7323
rect 40303 7289 40471 7323
rect 40675 7289 40843 7323
rect 41047 7289 41215 7323
rect 41419 7289 41587 7323
rect 41791 7289 41959 7323
rect 42163 7289 42331 7323
rect 42535 7289 42703 7323
rect 42907 7289 43075 7323
rect 43279 7289 43447 7323
rect 43651 7289 43819 7323
rect 44023 7289 44191 7323
rect 44395 7289 44563 7323
rect 44767 7289 44935 7323
rect 45139 7289 45307 7323
rect 45511 7289 45679 7323
rect 45883 7289 46051 7323
rect 46255 7289 46423 7323
rect 46627 7289 46795 7323
rect 46999 7289 47167 7323
rect 47371 7289 47539 7323
rect 47743 7289 47911 7323
rect 48115 7289 48283 7323
rect 48487 7289 48655 7323
rect 48859 7289 49027 7323
rect 49231 7289 49399 7323
rect 49603 7289 49771 7323
rect 39468 6837 39538 6854
rect 39840 6837 39910 6854
rect 40212 6837 40282 6854
rect 40584 6837 40654 6854
rect 40956 6837 41026 6854
rect 41328 6837 41398 6854
rect 41700 6837 41770 6854
rect 42072 6837 42142 6854
rect 42334 6837 42404 6854
rect 39468 6803 39479 6837
rect 39479 6803 39538 6837
rect 39840 6803 39910 6837
rect 40212 6803 40282 6837
rect 40584 6803 40654 6837
rect 40956 6803 41026 6837
rect 41328 6803 41398 6837
rect 41700 6803 41770 6837
rect 42072 6803 42142 6837
rect 42334 6803 42404 6837
rect 39468 6784 39538 6803
rect 39840 6784 39910 6803
rect 40212 6784 40282 6803
rect 40584 6784 40654 6803
rect 40956 6784 41026 6803
rect 41328 6784 41398 6803
rect 41700 6784 41770 6803
rect 42072 6784 42142 6803
rect 42334 6784 42404 6803
rect 39559 6701 39727 6735
rect 39931 6701 40099 6735
rect 40303 6701 40471 6735
rect 40675 6701 40843 6735
rect 41047 6701 41215 6735
rect 41419 6701 41587 6735
rect 41791 6701 41959 6735
rect 42163 6701 42331 6735
rect 39497 5866 39531 6642
rect 39755 5866 39789 6642
rect 39869 5866 39903 6642
rect 40127 5866 40161 6642
rect 40241 5866 40275 6642
rect 40499 5866 40533 6642
rect 40613 5866 40647 6642
rect 40871 5866 40905 6642
rect 40985 5866 41019 6642
rect 41243 5866 41277 6642
rect 41357 5866 41391 6642
rect 41615 5866 41649 6642
rect 41729 5866 41763 6642
rect 41987 5866 42021 6642
rect 42101 5866 42135 6642
rect 42359 5866 42393 6642
rect 39559 5773 39727 5807
rect 39931 5773 40099 5807
rect 40303 5773 40471 5807
rect 40675 5773 40843 5807
rect 41047 5773 41215 5807
rect 41419 5773 41587 5807
rect 41791 5773 41959 5807
rect 42163 5773 42331 5807
rect 39559 5665 39727 5699
rect 39931 5665 40099 5699
rect 40303 5665 40471 5699
rect 40675 5665 40843 5699
rect 41047 5665 41215 5699
rect 41419 5665 41587 5699
rect 41791 5665 41959 5699
rect 42163 5665 42331 5699
rect 39497 4830 39531 5606
rect 39755 4830 39789 5606
rect 39869 4830 39903 5606
rect 40127 4830 40161 5606
rect 40241 4830 40275 5606
rect 40499 4830 40533 5606
rect 40613 4830 40647 5606
rect 40871 4830 40905 5606
rect 40985 4830 41019 5606
rect 41243 4830 41277 5606
rect 41357 4830 41391 5606
rect 41615 4830 41649 5606
rect 41729 4830 41763 5606
rect 41987 4830 42021 5606
rect 42101 4830 42135 5606
rect 42359 4830 42393 5606
rect 39559 4737 39727 4771
rect 39931 4737 40099 4771
rect 40303 4737 40471 4771
rect 40675 4737 40843 4771
rect 41047 4737 41215 4771
rect 41419 4737 41587 4771
rect 41791 4737 41959 4771
rect 42163 4737 42331 4771
rect 39559 4629 39727 4663
rect 39931 4629 40099 4663
rect 40303 4629 40471 4663
rect 40675 4629 40843 4663
rect 41047 4629 41215 4663
rect 41419 4629 41587 4663
rect 41791 4629 41959 4663
rect 42163 4629 42331 4663
rect 39497 3794 39531 4570
rect 39755 3794 39789 4570
rect 39869 3794 39903 4570
rect 40127 3794 40161 4570
rect 40241 3794 40275 4570
rect 40499 3794 40533 4570
rect 40613 3794 40647 4570
rect 40871 3794 40905 4570
rect 40985 3794 41019 4570
rect 41243 3794 41277 4570
rect 41357 3794 41391 4570
rect 41615 3794 41649 4570
rect 41729 3794 41763 4570
rect 41987 3794 42021 4570
rect 42101 3794 42135 4570
rect 42359 3794 42393 4570
rect 39559 3701 39727 3735
rect 39931 3701 40099 3735
rect 40303 3701 40471 3735
rect 40675 3701 40843 3735
rect 41047 3701 41215 3735
rect 41419 3701 41587 3735
rect 41791 3701 41959 3735
rect 42163 3701 42331 3735
rect 39559 3593 39727 3627
rect 39931 3593 40099 3627
rect 40303 3593 40471 3627
rect 40675 3593 40843 3627
rect 41047 3593 41215 3627
rect 41419 3593 41587 3627
rect 41791 3593 41959 3627
rect 42163 3593 42331 3627
rect 39497 2758 39531 3534
rect 39755 2758 39789 3534
rect 39869 2758 39903 3534
rect 40127 2758 40161 3534
rect 40241 2758 40275 3534
rect 40499 2758 40533 3534
rect 40613 2758 40647 3534
rect 40871 2758 40905 3534
rect 40985 2758 41019 3534
rect 41243 2758 41277 3534
rect 41357 2758 41391 3534
rect 41615 2758 41649 3534
rect 41729 2758 41763 3534
rect 41987 2758 42021 3534
rect 42101 2758 42135 3534
rect 42359 2758 42393 3534
rect 39559 2665 39727 2699
rect 39931 2665 40099 2699
rect 40303 2665 40471 2699
rect 40675 2665 40843 2699
rect 41047 2665 41215 2699
rect 41419 2665 41587 2699
rect 41791 2665 41959 2699
rect 42163 2665 42331 2699
rect 43155 4378 43193 4775
rect 43290 4596 43305 4658
rect 43305 4596 43339 4658
rect 43339 4596 43354 4658
rect 43290 4196 43305 4258
rect 43305 4196 43339 4258
rect 43339 4196 43354 4258
rect 43290 3796 43305 3858
rect 43305 3796 43339 3858
rect 43339 3796 43354 3858
rect 43155 3387 43193 3784
rect 43290 3396 43305 3458
rect 43305 3396 43339 3458
rect 43339 3396 43354 3458
rect 39559 2007 39727 2041
rect 39931 2007 40099 2041
rect 40303 2007 40471 2041
rect 40675 2007 40843 2041
rect 41047 2007 41215 2041
rect 41419 2007 41587 2041
rect 41791 2007 41959 2041
rect 42163 2007 42331 2041
rect 42535 2007 42703 2041
rect 42907 2007 43075 2041
rect 43279 2007 43447 2041
rect 43651 2007 43819 2041
rect 44023 2007 44191 2041
rect 44395 2007 44563 2041
rect 44767 2007 44935 2041
rect 45139 2007 45307 2041
rect 45511 2007 45679 2041
rect 45883 2007 46051 2041
rect 46255 2007 46423 2041
rect 46627 2007 46795 2041
rect 46999 2007 47167 2041
rect 47371 2007 47539 2041
rect 47743 2007 47911 2041
rect 48115 2007 48283 2041
rect 39497 1781 39531 1957
rect 39755 1781 39789 1957
rect 39869 1781 39903 1957
rect 40127 1781 40161 1957
rect 40241 1781 40275 1957
rect 40499 1781 40533 1957
rect 40613 1781 40647 1957
rect 40871 1781 40905 1957
rect 40985 1781 41019 1957
rect 41243 1781 41277 1957
rect 41357 1781 41391 1957
rect 41615 1781 41649 1957
rect 41729 1781 41763 1957
rect 41987 1781 42021 1957
rect 42101 1781 42135 1957
rect 42359 1781 42393 1957
rect 42473 1781 42507 1957
rect 42731 1781 42765 1957
rect 42845 1781 42879 1957
rect 43103 1781 43137 1957
rect 43217 1781 43251 1957
rect 43475 1781 43509 1957
rect 43589 1781 43623 1957
rect 43847 1781 43881 1957
rect 43961 1781 43995 1957
rect 44219 1781 44253 1957
rect 44333 1781 44367 1957
rect 44591 1781 44625 1957
rect 44705 1781 44739 1957
rect 44963 1781 44997 1957
rect 45077 1781 45111 1957
rect 45335 1781 45369 1957
rect 45449 1781 45483 1957
rect 45707 1781 45741 1957
rect 45821 1781 45855 1957
rect 46079 1781 46113 1957
rect 46193 1781 46227 1957
rect 46451 1781 46485 1957
rect 46565 1781 46599 1957
rect 46823 1781 46857 1957
rect 46937 1781 46971 1957
rect 47195 1781 47229 1957
rect 47309 1781 47343 1957
rect 47567 1781 47601 1957
rect 47681 1781 47715 1957
rect 47939 1781 47973 1957
rect 48053 1781 48087 1957
rect 48311 1781 48345 1957
rect 39559 1697 39727 1731
rect 39931 1697 40099 1731
rect 40303 1697 40471 1731
rect 40675 1697 40843 1731
rect 41047 1697 41215 1731
rect 41419 1697 41587 1731
rect 41791 1697 41959 1731
rect 42163 1697 42331 1731
rect 42535 1697 42703 1731
rect 42907 1697 43075 1731
rect 43279 1697 43447 1731
rect 43651 1697 43819 1731
rect 44023 1697 44191 1731
rect 44395 1697 44563 1731
rect 44767 1697 44935 1731
rect 45139 1697 45307 1731
rect 45511 1697 45679 1731
rect 45883 1697 46051 1731
rect 46255 1697 46423 1731
rect 46627 1697 46795 1731
rect 46999 1697 47167 1731
rect 47371 1697 47539 1731
rect 47743 1697 47911 1731
rect 48115 1697 48283 1731
rect 39559 1589 39727 1623
rect 39931 1589 40099 1623
rect 40303 1589 40471 1623
rect 40675 1589 40843 1623
rect 41047 1589 41215 1623
rect 41419 1589 41587 1623
rect 41791 1589 41959 1623
rect 42163 1589 42331 1623
rect 42535 1589 42703 1623
rect 42907 1589 43075 1623
rect 43279 1589 43447 1623
rect 43651 1589 43819 1623
rect 44023 1589 44191 1623
rect 44395 1589 44563 1623
rect 44767 1589 44935 1623
rect 45139 1589 45307 1623
rect 45511 1589 45679 1623
rect 45883 1589 46051 1623
rect 46255 1589 46423 1623
rect 46627 1589 46795 1623
rect 46999 1589 47167 1623
rect 47371 1589 47539 1623
rect 47743 1589 47911 1623
rect 48115 1589 48283 1623
rect 39497 1363 39531 1539
rect 39755 1363 39789 1539
rect 39869 1363 39903 1539
rect 40127 1363 40161 1539
rect 40241 1363 40275 1539
rect 40499 1363 40533 1539
rect 40613 1363 40647 1539
rect 40871 1363 40905 1539
rect 40985 1363 41019 1539
rect 41243 1363 41277 1539
rect 41357 1363 41391 1539
rect 41615 1363 41649 1539
rect 41729 1363 41763 1539
rect 41987 1363 42021 1539
rect 42101 1363 42135 1539
rect 42359 1363 42393 1539
rect 42473 1363 42507 1539
rect 42731 1363 42765 1539
rect 42845 1363 42879 1539
rect 43103 1363 43137 1539
rect 43217 1363 43251 1539
rect 43475 1363 43509 1539
rect 43589 1363 43623 1539
rect 43847 1363 43881 1539
rect 43961 1363 43995 1539
rect 44219 1363 44253 1539
rect 44333 1363 44367 1539
rect 44591 1363 44625 1539
rect 44705 1363 44739 1539
rect 44963 1363 44997 1539
rect 45077 1363 45111 1539
rect 45335 1363 45369 1539
rect 45449 1363 45483 1539
rect 45707 1363 45741 1539
rect 45821 1363 45855 1539
rect 46079 1363 46113 1539
rect 46193 1363 46227 1539
rect 46451 1363 46485 1539
rect 46565 1363 46599 1539
rect 46823 1363 46857 1539
rect 46937 1363 46971 1539
rect 47195 1363 47229 1539
rect 47309 1363 47343 1539
rect 47567 1363 47601 1539
rect 47681 1363 47715 1539
rect 47939 1363 47973 1539
rect 48053 1363 48087 1539
rect 48311 1363 48345 1539
rect 39559 1279 39727 1313
rect 39931 1279 40099 1313
rect 40303 1279 40471 1313
rect 40675 1279 40843 1313
rect 41047 1279 41215 1313
rect 41419 1279 41587 1313
rect 41791 1279 41959 1313
rect 42163 1279 42331 1313
rect 42535 1279 42703 1313
rect 42907 1279 43075 1313
rect 43279 1279 43447 1313
rect 43651 1279 43819 1313
rect 44023 1279 44191 1313
rect 44395 1279 44563 1313
rect 44767 1279 44935 1313
rect 45139 1279 45307 1313
rect 45511 1279 45679 1313
rect 45883 1279 46051 1313
rect 46255 1279 46423 1313
rect 46627 1279 46795 1313
rect 46999 1279 47167 1313
rect 47371 1279 47539 1313
rect 47743 1279 47911 1313
rect 48115 1279 48283 1313
rect 39559 1171 39727 1205
rect 39931 1171 40099 1205
rect 40303 1171 40471 1205
rect 40675 1171 40843 1205
rect 41047 1171 41215 1205
rect 41419 1171 41587 1205
rect 41791 1171 41959 1205
rect 42163 1171 42331 1205
rect 42535 1171 42703 1205
rect 42907 1171 43075 1205
rect 43279 1171 43447 1205
rect 43651 1171 43819 1205
rect 44023 1171 44191 1205
rect 44395 1171 44563 1205
rect 44767 1171 44935 1205
rect 45139 1171 45307 1205
rect 45511 1171 45679 1205
rect 45883 1171 46051 1205
rect 46255 1171 46423 1205
rect 46627 1171 46795 1205
rect 46999 1171 47167 1205
rect 47371 1171 47539 1205
rect 47743 1171 47911 1205
rect 48115 1171 48283 1205
rect 39497 945 39531 1121
rect 39755 945 39789 1121
rect 39869 945 39903 1121
rect 40127 945 40161 1121
rect 40241 945 40275 1121
rect 40499 945 40533 1121
rect 40613 945 40647 1121
rect 40871 945 40905 1121
rect 40985 945 41019 1121
rect 41243 945 41277 1121
rect 41357 945 41391 1121
rect 41615 945 41649 1121
rect 41729 945 41763 1121
rect 41987 945 42021 1121
rect 42101 945 42135 1121
rect 42359 945 42393 1121
rect 42473 945 42507 1121
rect 42731 945 42765 1121
rect 42845 945 42879 1121
rect 43103 945 43137 1121
rect 43217 945 43251 1121
rect 43475 945 43509 1121
rect 43589 945 43623 1121
rect 43847 945 43881 1121
rect 43961 945 43995 1121
rect 44219 945 44253 1121
rect 44333 945 44367 1121
rect 44591 945 44625 1121
rect 44705 945 44739 1121
rect 44963 945 44997 1121
rect 45077 945 45111 1121
rect 45335 945 45369 1121
rect 45449 945 45483 1121
rect 45707 945 45741 1121
rect 45821 945 45855 1121
rect 46079 945 46113 1121
rect 46193 945 46227 1121
rect 46451 945 46485 1121
rect 46565 945 46599 1121
rect 46823 945 46857 1121
rect 46937 945 46971 1121
rect 47195 945 47229 1121
rect 47309 945 47343 1121
rect 47567 945 47601 1121
rect 47681 945 47715 1121
rect 47939 945 47973 1121
rect 48053 945 48087 1121
rect 48311 945 48345 1121
rect 39559 861 39727 895
rect 39931 861 40099 895
rect 40303 861 40471 895
rect 40675 861 40843 895
rect 41047 861 41215 895
rect 41419 861 41587 895
rect 41791 861 41959 895
rect 42163 861 42331 895
rect 42535 861 42703 895
rect 42907 861 43075 895
rect 43279 861 43447 895
rect 43651 861 43819 895
rect 44023 861 44191 895
rect 44395 861 44563 895
rect 44767 861 44935 895
rect 45139 861 45307 895
rect 45511 861 45679 895
rect 45883 861 46051 895
rect 46255 861 46423 895
rect 46627 861 46795 895
rect 46999 861 47167 895
rect 47371 861 47539 895
rect 47743 861 47911 895
rect 48115 861 48283 895
rect 39559 753 39727 787
rect 39931 753 40099 787
rect 40303 753 40471 787
rect 40675 753 40843 787
rect 41047 753 41215 787
rect 41419 753 41587 787
rect 41791 753 41959 787
rect 42163 753 42331 787
rect 42535 753 42703 787
rect 42907 753 43075 787
rect 43279 753 43447 787
rect 43651 753 43819 787
rect 44023 753 44191 787
rect 44395 753 44563 787
rect 44767 753 44935 787
rect 45139 753 45307 787
rect 45511 753 45679 787
rect 45883 753 46051 787
rect 46255 753 46423 787
rect 46627 753 46795 787
rect 46999 753 47167 787
rect 47371 753 47539 787
rect 47743 753 47911 787
rect 48115 753 48283 787
rect 39497 527 39531 703
rect 39755 527 39789 703
rect 39869 527 39903 703
rect 40127 527 40161 703
rect 40241 527 40275 703
rect 40499 527 40533 703
rect 40613 527 40647 703
rect 40871 527 40905 703
rect 40985 527 41019 703
rect 41243 527 41277 703
rect 41357 527 41391 703
rect 41615 527 41649 703
rect 41729 527 41763 703
rect 41987 527 42021 703
rect 42101 527 42135 703
rect 42359 527 42393 703
rect 42473 527 42507 703
rect 42731 527 42765 703
rect 42845 527 42879 703
rect 43103 527 43137 703
rect 43217 527 43251 703
rect 43475 527 43509 703
rect 43589 527 43623 703
rect 43847 527 43881 703
rect 43961 527 43995 703
rect 44219 527 44253 703
rect 44333 527 44367 703
rect 44591 527 44625 703
rect 44705 527 44739 703
rect 44963 527 44997 703
rect 45077 527 45111 703
rect 45335 527 45369 703
rect 45449 527 45483 703
rect 45707 527 45741 703
rect 45821 527 45855 703
rect 46079 527 46113 703
rect 46193 527 46227 703
rect 46451 527 46485 703
rect 46565 527 46599 703
rect 46823 527 46857 703
rect 46937 527 46971 703
rect 47195 527 47229 703
rect 47309 527 47343 703
rect 47567 527 47601 703
rect 47681 527 47715 703
rect 47939 527 47973 703
rect 48053 527 48087 703
rect 48311 527 48345 703
rect 39559 443 39727 477
rect 39931 443 40099 477
rect 40303 443 40471 477
rect 40675 443 40843 477
rect 41047 443 41215 477
rect 41419 443 41587 477
rect 41791 443 41959 477
rect 42163 443 42331 477
rect 42535 443 42703 477
rect 42907 443 43075 477
rect 43279 443 43447 477
rect 43651 443 43819 477
rect 44023 443 44191 477
rect 44395 443 44563 477
rect 44767 443 44935 477
rect 45139 443 45307 477
rect 45511 443 45679 477
rect 45883 443 46051 477
rect 46255 443 46423 477
rect 46627 443 46795 477
rect 46999 443 47167 477
rect 47371 443 47539 477
rect 47743 443 47911 477
rect 48115 443 48283 477
rect 39498 375 39568 386
rect 40166 375 40236 394
rect 40910 375 40980 394
rect 41654 375 41724 394
rect 42398 375 42468 394
rect 43142 375 43212 394
rect 43886 375 43956 394
rect 44630 375 44700 394
rect 45374 375 45444 394
rect 46118 375 46188 394
rect 46862 375 46932 394
rect 47606 375 47676 394
rect 48268 375 48338 390
rect 39498 341 39568 375
rect 40166 341 40236 375
rect 40910 341 40980 375
rect 41654 341 41724 375
rect 42398 341 42468 375
rect 43142 341 43212 375
rect 43886 341 43956 375
rect 44630 341 44700 375
rect 45374 341 45444 375
rect 46118 341 46188 375
rect 46862 341 46932 375
rect 47606 341 47676 375
rect 48268 341 48338 375
rect 39498 316 39568 341
rect 40166 324 40236 341
rect 40910 324 40980 341
rect 41654 324 41724 341
rect 42398 324 42468 341
rect 43142 324 43212 341
rect 43886 324 43956 341
rect 44630 324 44700 341
rect 45374 324 45444 341
rect 46118 324 46188 341
rect 46862 324 46932 341
rect 47606 324 47676 341
rect 48268 320 48338 341
<< metal1 >>
rect 35518 10928 35528 11896
rect 36446 10928 36456 11896
rect 35850 7216 36126 10928
rect 38230 9324 38240 9524
rect 38440 9324 38450 9524
rect 38974 9324 38984 9524
rect 39184 9324 39194 9524
rect 39718 9324 39728 9524
rect 39928 9324 39938 9524
rect 40462 9324 40472 9524
rect 40672 9324 40682 9524
rect 41206 9324 41216 9524
rect 41416 9324 41426 9524
rect 41950 9324 41960 9524
rect 42160 9324 42170 9524
rect 42694 9324 42704 9524
rect 42904 9324 42914 9524
rect 43438 9324 43448 9524
rect 43648 9324 43658 9524
rect 43810 9324 43820 9524
rect 44020 9324 44030 9524
rect 44554 9324 44564 9524
rect 44764 9324 44774 9524
rect 45298 9324 45308 9524
rect 45508 9324 45518 9524
rect 46042 9324 46052 9524
rect 46252 9324 46262 9524
rect 46786 9324 46796 9524
rect 46996 9324 47006 9524
rect 47530 9324 47540 9524
rect 47740 9324 47750 9524
rect 48274 9324 48284 9524
rect 48484 9324 48494 9524
rect 49018 9324 49028 9524
rect 49228 9324 49238 9524
rect 49762 9324 49772 9524
rect 49972 9324 49982 9524
rect 38312 9248 38370 9324
rect 39056 9248 39114 9324
rect 39800 9248 39858 9324
rect 40544 9248 40602 9324
rect 41288 9248 41346 9324
rect 42032 9248 42090 9324
rect 42776 9248 42834 9324
rect 43500 9314 43578 9324
rect 43520 9248 43578 9314
rect 43930 9248 43982 9324
rect 44636 9248 44694 9324
rect 45380 9248 45438 9324
rect 46124 9248 46182 9324
rect 46868 9248 46926 9324
rect 47612 9248 47670 9324
rect 48356 9248 48414 9324
rect 49100 9248 49158 9324
rect 49826 9308 49902 9324
rect 49826 9248 49884 9308
rect 38294 9242 38388 9248
rect 38294 9172 38306 9242
rect 38376 9172 38388 9242
rect 38294 9166 38388 9172
rect 39038 9242 39132 9248
rect 39038 9172 39050 9242
rect 39120 9172 39132 9242
rect 39038 9166 39132 9172
rect 39782 9242 39876 9248
rect 39782 9172 39794 9242
rect 39864 9172 39876 9242
rect 39782 9166 39876 9172
rect 40526 9242 40620 9248
rect 40526 9172 40538 9242
rect 40608 9172 40620 9242
rect 40526 9166 40620 9172
rect 41270 9242 41364 9248
rect 41270 9172 41282 9242
rect 41352 9172 41364 9242
rect 41270 9166 41364 9172
rect 42014 9242 42108 9248
rect 42014 9172 42026 9242
rect 42096 9172 42108 9242
rect 42014 9166 42108 9172
rect 42758 9242 42852 9248
rect 42758 9172 42770 9242
rect 42840 9172 42852 9242
rect 42758 9166 42852 9172
rect 43502 9242 43596 9248
rect 43502 9172 43514 9242
rect 43584 9172 43596 9242
rect 43502 9166 43596 9172
rect 43874 9242 43982 9248
rect 43874 9172 43886 9242
rect 43956 9172 43982 9242
rect 43874 9166 43982 9172
rect 44618 9242 44712 9248
rect 44618 9172 44630 9242
rect 44700 9172 44712 9242
rect 44618 9166 44712 9172
rect 45362 9242 45456 9248
rect 45362 9172 45374 9242
rect 45444 9172 45456 9242
rect 45362 9166 45456 9172
rect 46106 9242 46200 9248
rect 46106 9172 46118 9242
rect 46188 9172 46200 9242
rect 46106 9166 46200 9172
rect 46850 9242 46944 9248
rect 46850 9172 46862 9242
rect 46932 9172 46944 9242
rect 46850 9166 46944 9172
rect 47594 9242 47688 9248
rect 47594 9172 47606 9242
rect 47676 9172 47688 9242
rect 47594 9166 47688 9172
rect 48338 9242 48432 9248
rect 48338 9172 48350 9242
rect 48420 9172 48432 9242
rect 48338 9166 48432 9172
rect 49082 9242 49176 9248
rect 49082 9172 49094 9242
rect 49164 9172 49176 9242
rect 49082 9166 49176 9172
rect 49772 9242 49884 9248
rect 49772 9172 49784 9242
rect 49854 9172 49884 9242
rect 49772 9166 49884 9172
rect 38002 9076 38070 9136
rect 38240 9129 38250 9136
rect 38240 9083 38251 9129
rect 38240 9076 38250 9083
rect 38002 9030 38050 9076
rect 38312 9042 38370 9166
rect 38432 9129 38442 9136
rect 38431 9083 38442 9129
rect 38612 9129 38622 9136
rect 38804 9129 38814 9136
rect 38432 9076 38442 9083
rect 38612 9083 38623 9129
rect 38803 9083 38814 9129
rect 38984 9129 38994 9136
rect 38612 9076 38622 9083
rect 38804 9076 38814 9083
rect 38984 9083 38995 9129
rect 38984 9076 38994 9083
rect 39056 9042 39114 9166
rect 39176 9129 39186 9136
rect 39175 9083 39186 9129
rect 39176 9076 39186 9083
rect 39356 9076 39558 9136
rect 39728 9129 39738 9136
rect 39728 9083 39739 9129
rect 39728 9076 39738 9083
rect 39428 9042 39486 9076
rect 39800 9042 39858 9166
rect 39920 9129 39930 9136
rect 39919 9083 39930 9129
rect 40100 9129 40110 9136
rect 40292 9129 40302 9136
rect 39920 9076 39930 9083
rect 40100 9083 40111 9129
rect 40291 9083 40302 9129
rect 40472 9129 40482 9136
rect 40100 9076 40110 9083
rect 40292 9076 40302 9083
rect 40472 9083 40483 9129
rect 40472 9076 40482 9083
rect 40544 9042 40602 9166
rect 40664 9129 40674 9136
rect 40663 9083 40674 9129
rect 40664 9076 40674 9083
rect 40844 9076 41046 9136
rect 41216 9129 41226 9136
rect 41216 9083 41227 9129
rect 41216 9076 41226 9083
rect 40916 9042 40974 9076
rect 41288 9042 41346 9166
rect 41408 9129 41418 9136
rect 41407 9083 41418 9129
rect 41588 9129 41598 9136
rect 41780 9129 41790 9136
rect 41408 9076 41418 9083
rect 41588 9083 41599 9129
rect 41779 9083 41790 9129
rect 41960 9129 41970 9136
rect 41588 9076 41598 9083
rect 41780 9076 41790 9083
rect 41960 9083 41971 9129
rect 41960 9076 41970 9083
rect 42032 9042 42090 9166
rect 42152 9129 42162 9136
rect 42151 9083 42162 9129
rect 42152 9076 42162 9083
rect 42332 9076 42534 9136
rect 42704 9129 42714 9136
rect 42704 9083 42715 9129
rect 42704 9076 42714 9083
rect 42404 9042 42462 9076
rect 42776 9042 42834 9166
rect 42896 9129 42906 9136
rect 42895 9083 42906 9129
rect 43076 9129 43086 9136
rect 43268 9129 43278 9136
rect 42896 9076 42906 9083
rect 43076 9083 43087 9129
rect 43267 9083 43278 9129
rect 43448 9129 43458 9136
rect 43076 9076 43086 9083
rect 43268 9076 43278 9083
rect 43448 9083 43459 9129
rect 43448 9076 43458 9083
rect 43520 9042 43578 9166
rect 43640 9129 43650 9136
rect 43639 9083 43650 9129
rect 43640 9076 43650 9083
rect 43820 9076 43892 9136
rect 38002 8654 38009 9030
rect 38043 8654 38050 9030
rect 38002 8602 38050 8654
rect 38261 9030 38421 9042
rect 38261 8654 38267 9030
rect 38301 8654 38381 9030
rect 38415 8654 38421 9030
rect 38261 8642 38421 8654
rect 38633 9030 38793 9042
rect 38633 8654 38639 9030
rect 38673 8654 38753 9030
rect 38787 8654 38793 9030
rect 38633 8642 38793 8654
rect 39005 9030 39165 9042
rect 39005 8654 39011 9030
rect 39045 8654 39125 9030
rect 39159 8654 39165 9030
rect 39005 8642 39165 8654
rect 39377 9030 39537 9042
rect 39377 8654 39383 9030
rect 39417 8654 39497 9030
rect 39531 8654 39537 9030
rect 39377 8642 39537 8654
rect 39749 9030 39909 9042
rect 39749 8654 39755 9030
rect 39789 8654 39869 9030
rect 39903 8654 39909 9030
rect 39749 8642 39909 8654
rect 40121 9030 40281 9042
rect 40121 8654 40127 9030
rect 40161 8654 40241 9030
rect 40275 8654 40281 9030
rect 40121 8642 40281 8654
rect 40493 9030 40653 9042
rect 40493 8654 40499 9030
rect 40533 8654 40613 9030
rect 40647 8654 40653 9030
rect 40493 8642 40653 8654
rect 40865 9030 41025 9042
rect 40865 8654 40871 9030
rect 40905 8654 40985 9030
rect 41019 8654 41025 9030
rect 40865 8642 41025 8654
rect 41237 9030 41397 9042
rect 41237 8654 41243 9030
rect 41277 8654 41357 9030
rect 41391 8654 41397 9030
rect 41237 8642 41397 8654
rect 41609 9030 41769 9042
rect 41609 8654 41615 9030
rect 41649 8654 41729 9030
rect 41763 8654 41769 9030
rect 41609 8642 41769 8654
rect 41981 9030 42141 9042
rect 41981 8654 41987 9030
rect 42021 8654 42101 9030
rect 42135 8654 42141 9030
rect 41981 8642 42141 8654
rect 42353 9030 42513 9042
rect 42353 8654 42359 9030
rect 42393 8654 42473 9030
rect 42507 8654 42513 9030
rect 42353 8642 42513 8654
rect 42725 9030 42885 9042
rect 42725 8654 42731 9030
rect 42765 8654 42845 9030
rect 42879 8654 42885 9030
rect 42725 8642 42885 8654
rect 43097 9030 43257 9042
rect 43097 8654 43103 9030
rect 43137 8654 43217 9030
rect 43251 8654 43257 9030
rect 43097 8642 43257 8654
rect 43469 9030 43629 9042
rect 43469 8654 43475 9030
rect 43509 8654 43589 9030
rect 43623 8654 43629 9030
rect 43469 8642 43629 8654
rect 43840 9030 43892 9076
rect 43840 8654 43847 9030
rect 43881 8654 43892 9030
rect 38002 8601 38090 8602
rect 38002 8596 38251 8601
rect 38002 8452 38070 8596
rect 38240 8555 38251 8596
rect 38240 8493 38250 8555
rect 38240 8452 38251 8493
rect 38002 8447 38251 8452
rect 38002 8446 38088 8447
rect 38002 8394 38050 8446
rect 38306 8406 38376 8642
rect 38431 8596 38623 8601
rect 38431 8555 38442 8596
rect 38432 8493 38442 8555
rect 38431 8452 38442 8493
rect 38612 8555 38623 8596
rect 38612 8493 38622 8555
rect 38612 8452 38623 8493
rect 38431 8447 38623 8452
rect 38678 8406 38748 8642
rect 38803 8596 38995 8601
rect 38803 8555 38814 8596
rect 38804 8493 38814 8555
rect 38803 8452 38814 8493
rect 38984 8555 38995 8596
rect 38984 8493 38994 8555
rect 38984 8452 38995 8493
rect 38803 8447 38995 8452
rect 39050 8406 39120 8642
rect 39175 8600 39367 8601
rect 39422 8600 39492 8642
rect 39547 8600 39739 8601
rect 39175 8596 39739 8600
rect 39175 8555 39186 8596
rect 39176 8493 39186 8555
rect 39175 8452 39186 8493
rect 39356 8452 39558 8596
rect 39728 8555 39739 8596
rect 39728 8493 39738 8555
rect 39728 8452 39739 8493
rect 39175 8448 39739 8452
rect 39175 8447 39367 8448
rect 39422 8406 39492 8448
rect 39547 8447 39739 8448
rect 39794 8406 39864 8642
rect 39919 8596 40111 8601
rect 39919 8555 39930 8596
rect 39920 8493 39930 8555
rect 39919 8452 39930 8493
rect 40100 8555 40111 8596
rect 40100 8493 40110 8555
rect 40100 8452 40111 8493
rect 39919 8447 40111 8452
rect 40166 8406 40236 8642
rect 40291 8596 40483 8601
rect 40291 8555 40302 8596
rect 40292 8493 40302 8555
rect 40291 8452 40302 8493
rect 40472 8555 40483 8596
rect 40472 8493 40482 8555
rect 40472 8452 40483 8493
rect 40291 8447 40483 8452
rect 40538 8406 40608 8642
rect 40910 8602 40980 8642
rect 40718 8601 41136 8602
rect 40663 8596 41227 8601
rect 40663 8555 40674 8596
rect 40664 8493 40674 8555
rect 40663 8452 40674 8493
rect 40844 8452 41046 8596
rect 41216 8555 41227 8596
rect 41216 8493 41226 8555
rect 41216 8452 41227 8493
rect 40663 8447 41227 8452
rect 40718 8446 41136 8447
rect 40910 8406 40980 8446
rect 41282 8406 41352 8642
rect 41407 8596 41599 8601
rect 41407 8555 41418 8596
rect 41408 8493 41418 8555
rect 41407 8452 41418 8493
rect 41588 8555 41599 8596
rect 41588 8493 41598 8555
rect 41588 8452 41599 8493
rect 41407 8447 41599 8452
rect 41654 8406 41724 8642
rect 41779 8596 41971 8601
rect 41779 8555 41790 8596
rect 41780 8493 41790 8555
rect 41779 8452 41790 8493
rect 41960 8555 41971 8596
rect 41960 8493 41970 8555
rect 41960 8452 41971 8493
rect 41779 8447 41971 8452
rect 42026 8406 42096 8642
rect 42398 8602 42468 8642
rect 42246 8601 42622 8602
rect 42151 8596 42715 8601
rect 42151 8555 42162 8596
rect 42152 8493 42162 8555
rect 42151 8452 42162 8493
rect 42332 8452 42534 8596
rect 42704 8555 42715 8596
rect 42704 8493 42714 8555
rect 42704 8452 42715 8493
rect 42151 8447 42715 8452
rect 42246 8446 42622 8447
rect 42398 8406 42468 8446
rect 42770 8406 42840 8642
rect 42895 8596 43087 8601
rect 42895 8555 42906 8596
rect 42896 8493 42906 8555
rect 42895 8452 42906 8493
rect 43076 8555 43087 8596
rect 43076 8493 43086 8555
rect 43076 8452 43087 8493
rect 42895 8447 43087 8452
rect 43142 8406 43212 8642
rect 43267 8596 43459 8601
rect 43267 8555 43278 8596
rect 43268 8493 43278 8555
rect 43267 8452 43278 8493
rect 43448 8555 43459 8596
rect 43448 8493 43458 8555
rect 43448 8452 43459 8493
rect 43267 8447 43459 8452
rect 43514 8406 43584 8642
rect 43840 8602 43892 8654
rect 43734 8601 43892 8602
rect 43639 8596 43892 8601
rect 43639 8555 43650 8596
rect 43640 8493 43650 8555
rect 43639 8452 43650 8493
rect 43820 8452 43892 8596
rect 43639 8447 43892 8452
rect 43734 8446 43892 8447
rect 38002 8018 38009 8394
rect 38043 8018 38050 8394
rect 38002 7966 38050 8018
rect 38261 8394 38421 8406
rect 38261 8018 38267 8394
rect 38301 8018 38381 8394
rect 38415 8018 38421 8394
rect 38261 8006 38421 8018
rect 38633 8394 38793 8406
rect 38633 8018 38639 8394
rect 38673 8018 38753 8394
rect 38787 8018 38793 8394
rect 38633 8006 38793 8018
rect 39005 8394 39165 8406
rect 39005 8018 39011 8394
rect 39045 8018 39125 8394
rect 39159 8018 39165 8394
rect 39005 8006 39165 8018
rect 39377 8394 39537 8406
rect 39377 8018 39383 8394
rect 39417 8018 39497 8394
rect 39531 8018 39537 8394
rect 39377 8006 39537 8018
rect 39749 8394 39909 8406
rect 39749 8018 39755 8394
rect 39789 8018 39869 8394
rect 39903 8018 39909 8394
rect 39749 8006 39909 8018
rect 40121 8394 40281 8406
rect 40121 8018 40127 8394
rect 40161 8018 40241 8394
rect 40275 8018 40281 8394
rect 40121 8006 40281 8018
rect 40493 8394 40653 8406
rect 40493 8018 40499 8394
rect 40533 8018 40613 8394
rect 40647 8018 40653 8394
rect 40493 8006 40653 8018
rect 40865 8394 41025 8406
rect 40865 8018 40871 8394
rect 40905 8018 40985 8394
rect 41019 8018 41025 8394
rect 40865 8006 41025 8018
rect 41237 8394 41397 8406
rect 41237 8018 41243 8394
rect 41277 8018 41357 8394
rect 41391 8018 41397 8394
rect 41237 8006 41397 8018
rect 41609 8394 41769 8406
rect 41609 8018 41615 8394
rect 41649 8018 41729 8394
rect 41763 8018 41769 8394
rect 41609 8006 41769 8018
rect 41981 8394 42141 8406
rect 41981 8018 41987 8394
rect 42021 8018 42101 8394
rect 42135 8018 42141 8394
rect 41981 8006 42141 8018
rect 42353 8394 42513 8406
rect 42353 8018 42359 8394
rect 42393 8018 42473 8394
rect 42507 8018 42513 8394
rect 42353 8006 42513 8018
rect 42725 8394 42885 8406
rect 42725 8018 42731 8394
rect 42765 8018 42845 8394
rect 42879 8018 42885 8394
rect 42725 8006 42885 8018
rect 43097 8394 43257 8406
rect 43097 8018 43103 8394
rect 43137 8018 43217 8394
rect 43251 8018 43257 8394
rect 43097 8006 43257 8018
rect 43469 8394 43629 8406
rect 43469 8018 43475 8394
rect 43509 8018 43589 8394
rect 43623 8018 43629 8394
rect 43469 8006 43629 8018
rect 43840 8394 43892 8446
rect 43840 8018 43847 8394
rect 43881 8018 43892 8394
rect 38002 7965 38092 7966
rect 38002 7960 38251 7965
rect 38002 7816 38070 7960
rect 38240 7919 38251 7960
rect 38240 7857 38250 7919
rect 38240 7816 38251 7857
rect 38002 7811 38251 7816
rect 38002 7806 38092 7811
rect 38002 7758 38050 7806
rect 38306 7770 38376 8006
rect 38431 7960 38623 7965
rect 38431 7919 38442 7960
rect 38432 7857 38442 7919
rect 38431 7816 38442 7857
rect 38612 7919 38623 7960
rect 38612 7857 38622 7919
rect 38612 7816 38623 7857
rect 38431 7811 38623 7816
rect 38678 7770 38748 8006
rect 38803 7960 38995 7965
rect 38803 7919 38814 7960
rect 38804 7857 38814 7919
rect 38803 7816 38814 7857
rect 38984 7919 38995 7960
rect 38984 7857 38994 7919
rect 38984 7816 38995 7857
rect 38803 7811 38995 7816
rect 39050 7770 39120 8006
rect 39175 7962 39367 7965
rect 39422 7962 39492 8006
rect 39547 7962 39739 7965
rect 39175 7960 39739 7962
rect 39175 7919 39186 7960
rect 39176 7857 39186 7919
rect 39175 7816 39186 7857
rect 39356 7816 39558 7960
rect 39728 7919 39739 7960
rect 39728 7857 39738 7919
rect 39728 7816 39739 7857
rect 39175 7811 39739 7816
rect 39216 7810 39692 7811
rect 39422 7770 39492 7810
rect 39794 7770 39864 8006
rect 39919 7960 40111 7965
rect 39919 7919 39930 7960
rect 39920 7857 39930 7919
rect 39919 7816 39930 7857
rect 40100 7919 40111 7960
rect 40100 7857 40110 7919
rect 40100 7816 40111 7857
rect 39919 7811 40111 7816
rect 40166 7770 40236 8006
rect 40291 7960 40483 7965
rect 40291 7919 40302 7960
rect 40292 7857 40302 7919
rect 40291 7816 40302 7857
rect 40472 7919 40483 7960
rect 40472 7857 40482 7919
rect 40472 7816 40483 7857
rect 40291 7811 40483 7816
rect 40538 7770 40608 8006
rect 40910 7966 40980 8006
rect 40738 7965 41156 7966
rect 40663 7960 41227 7965
rect 40663 7919 40674 7960
rect 40664 7857 40674 7919
rect 40663 7816 40674 7857
rect 40844 7816 41046 7960
rect 41216 7919 41227 7960
rect 41216 7857 41226 7919
rect 41216 7816 41227 7857
rect 40663 7811 41227 7816
rect 40738 7810 41156 7811
rect 40910 7770 40980 7810
rect 41282 7770 41352 8006
rect 41407 7960 41599 7965
rect 41407 7919 41418 7960
rect 41408 7857 41418 7919
rect 41407 7816 41418 7857
rect 41588 7919 41599 7960
rect 41588 7857 41598 7919
rect 41588 7816 41599 7857
rect 41407 7811 41599 7816
rect 41654 7770 41724 8006
rect 41779 7960 41971 7965
rect 41779 7919 41790 7960
rect 41780 7857 41790 7919
rect 41779 7816 41790 7857
rect 41960 7919 41971 7960
rect 41960 7857 41970 7919
rect 41960 7816 41971 7857
rect 41779 7811 41971 7816
rect 42026 7770 42096 8006
rect 42398 7966 42468 8006
rect 42234 7965 42610 7966
rect 42151 7960 42715 7965
rect 42151 7919 42162 7960
rect 42152 7857 42162 7919
rect 42151 7816 42162 7857
rect 42332 7816 42534 7960
rect 42704 7919 42715 7960
rect 42704 7857 42714 7919
rect 42704 7816 42715 7857
rect 42151 7811 42715 7816
rect 42234 7810 42610 7811
rect 42398 7770 42468 7810
rect 42770 7770 42840 8006
rect 42895 7960 43087 7965
rect 42895 7919 42906 7960
rect 42896 7857 42906 7919
rect 42895 7816 42906 7857
rect 43076 7919 43087 7960
rect 43076 7857 43086 7919
rect 43076 7816 43087 7857
rect 42895 7811 43087 7816
rect 43142 7770 43212 8006
rect 43267 7960 43459 7965
rect 43267 7919 43278 7960
rect 43268 7857 43278 7919
rect 43267 7816 43278 7857
rect 43448 7919 43459 7960
rect 43448 7857 43458 7919
rect 43448 7816 43459 7857
rect 43267 7811 43459 7816
rect 43514 7770 43584 8006
rect 43840 7966 43892 8018
rect 43750 7965 43892 7966
rect 43639 7960 43892 7965
rect 43639 7919 43650 7960
rect 43640 7857 43650 7919
rect 43639 7816 43650 7857
rect 43820 7816 43892 7960
rect 43639 7811 43892 7816
rect 43750 7810 43892 7811
rect 38002 7382 38009 7758
rect 38043 7382 38050 7758
rect 38002 7336 38050 7382
rect 38261 7758 38421 7770
rect 38261 7382 38267 7758
rect 38301 7382 38381 7758
rect 38415 7382 38421 7758
rect 38261 7370 38421 7382
rect 38633 7758 38793 7770
rect 38633 7382 38639 7758
rect 38673 7382 38753 7758
rect 38787 7382 38793 7758
rect 38633 7370 38793 7382
rect 39005 7758 39165 7770
rect 39005 7382 39011 7758
rect 39045 7382 39125 7758
rect 39159 7382 39165 7758
rect 39005 7370 39165 7382
rect 39377 7758 39537 7770
rect 39377 7382 39383 7758
rect 39417 7382 39497 7758
rect 39531 7382 39537 7758
rect 39377 7370 39537 7382
rect 39749 7758 39909 7770
rect 39749 7382 39755 7758
rect 39789 7382 39869 7758
rect 39903 7382 39909 7758
rect 39749 7370 39909 7382
rect 40121 7758 40281 7770
rect 40121 7382 40127 7758
rect 40161 7382 40241 7758
rect 40275 7382 40281 7758
rect 40121 7370 40281 7382
rect 40493 7758 40653 7770
rect 40493 7382 40499 7758
rect 40533 7382 40613 7758
rect 40647 7382 40653 7758
rect 40493 7370 40653 7382
rect 40865 7758 41025 7770
rect 40865 7382 40871 7758
rect 40905 7382 40985 7758
rect 41019 7382 41025 7758
rect 40865 7370 41025 7382
rect 41237 7758 41397 7770
rect 41237 7382 41243 7758
rect 41277 7382 41357 7758
rect 41391 7382 41397 7758
rect 41237 7370 41397 7382
rect 41609 7758 41769 7770
rect 41609 7382 41615 7758
rect 41649 7382 41729 7758
rect 41763 7382 41769 7758
rect 41609 7370 41769 7382
rect 41981 7758 42141 7770
rect 41981 7382 41987 7758
rect 42021 7382 42101 7758
rect 42135 7382 42141 7758
rect 41981 7370 42141 7382
rect 42353 7758 42513 7770
rect 42353 7382 42359 7758
rect 42393 7382 42473 7758
rect 42507 7382 42513 7758
rect 42353 7370 42513 7382
rect 42725 7758 42885 7770
rect 42725 7382 42731 7758
rect 42765 7382 42845 7758
rect 42879 7382 42885 7758
rect 42725 7370 42885 7382
rect 43097 7758 43257 7770
rect 43097 7382 43103 7758
rect 43137 7382 43217 7758
rect 43251 7382 43257 7758
rect 43097 7370 43257 7382
rect 43469 7758 43629 7770
rect 43469 7382 43475 7758
rect 43509 7382 43589 7758
rect 43623 7382 43629 7758
rect 43469 7370 43629 7382
rect 43840 7758 43892 7810
rect 43840 7382 43847 7758
rect 43881 7382 43892 7758
rect 38002 7276 38070 7336
rect 38240 7329 38250 7336
rect 38432 7329 38442 7336
rect 38240 7283 38251 7329
rect 38431 7283 38442 7329
rect 38612 7329 38622 7336
rect 38240 7276 38250 7283
rect 38432 7276 38442 7283
rect 38612 7283 38623 7329
rect 38612 7276 38622 7283
rect 35692 6594 35702 7216
rect 36308 6594 36318 7216
rect 38684 7028 38742 7370
rect 39428 7336 39486 7370
rect 38804 7329 38814 7336
rect 38803 7283 38814 7329
rect 38984 7329 38994 7336
rect 39176 7329 39186 7336
rect 38804 7276 38814 7283
rect 38984 7283 38995 7329
rect 39175 7283 39186 7329
rect 38984 7276 38994 7283
rect 39176 7276 39186 7283
rect 39356 7276 39558 7336
rect 39728 7329 39738 7336
rect 39920 7329 39930 7336
rect 39728 7283 39739 7329
rect 39919 7283 39930 7329
rect 40100 7329 40110 7336
rect 39728 7276 39738 7283
rect 39920 7276 39930 7283
rect 40100 7283 40111 7329
rect 40100 7276 40110 7283
rect 39302 7274 39632 7276
rect 40172 7028 40230 7370
rect 40916 7336 40974 7370
rect 40292 7329 40302 7336
rect 40291 7283 40302 7329
rect 40472 7329 40482 7336
rect 40664 7329 40674 7336
rect 40292 7276 40302 7283
rect 40472 7283 40483 7329
rect 40663 7283 40674 7329
rect 40472 7276 40482 7283
rect 40664 7276 40674 7283
rect 40844 7276 41046 7336
rect 41216 7329 41226 7336
rect 41408 7329 41418 7336
rect 41216 7283 41227 7329
rect 41407 7283 41418 7329
rect 41588 7329 41598 7336
rect 41216 7276 41226 7283
rect 41408 7276 41418 7283
rect 41588 7283 41599 7329
rect 41588 7276 41598 7283
rect 41660 7028 41718 7370
rect 42404 7336 42462 7370
rect 41780 7329 41790 7336
rect 41779 7283 41790 7329
rect 41960 7329 41970 7336
rect 42152 7329 42162 7336
rect 41780 7276 41790 7283
rect 41960 7283 41971 7329
rect 42151 7283 42162 7329
rect 41960 7276 41970 7283
rect 42152 7276 42162 7283
rect 42332 7276 42534 7336
rect 42704 7329 42714 7336
rect 42896 7329 42906 7336
rect 42704 7283 42715 7329
rect 42895 7283 42906 7329
rect 43076 7329 43086 7336
rect 42704 7276 42714 7283
rect 42896 7276 42906 7283
rect 43076 7283 43087 7329
rect 43076 7276 43086 7283
rect 43148 7028 43206 7370
rect 43840 7336 43892 7382
rect 43930 9042 43982 9166
rect 44016 9076 44022 9136
rect 44192 9129 44202 9136
rect 44384 9129 44394 9136
rect 44192 9083 44203 9129
rect 44383 9083 44394 9129
rect 44564 9129 44574 9136
rect 44192 9076 44202 9083
rect 44384 9076 44394 9083
rect 44564 9083 44575 9129
rect 44564 9076 44574 9083
rect 44636 9042 44694 9166
rect 44756 9129 44766 9136
rect 44755 9083 44766 9129
rect 44936 9129 44946 9136
rect 45128 9129 45138 9136
rect 44756 9076 44766 9083
rect 44936 9083 44947 9129
rect 45127 9083 45138 9129
rect 45308 9129 45318 9136
rect 44936 9076 44946 9083
rect 45128 9076 45138 9083
rect 45308 9083 45319 9129
rect 45308 9076 45318 9083
rect 45380 9042 45438 9166
rect 45500 9129 45510 9136
rect 45499 9083 45510 9129
rect 45680 9129 45690 9136
rect 45872 9129 45882 9136
rect 45500 9076 45510 9083
rect 45680 9083 45691 9129
rect 45871 9083 45882 9129
rect 46052 9129 46062 9136
rect 45680 9076 45690 9083
rect 45872 9076 45882 9083
rect 46052 9083 46063 9129
rect 46052 9076 46062 9083
rect 46124 9042 46182 9166
rect 46244 9129 46254 9136
rect 46243 9083 46254 9129
rect 46424 9129 46434 9136
rect 46616 9129 46626 9136
rect 46244 9076 46254 9083
rect 46424 9083 46435 9129
rect 46615 9083 46626 9129
rect 46796 9129 46806 9136
rect 46424 9076 46434 9083
rect 46616 9076 46626 9083
rect 46796 9083 46807 9129
rect 46796 9076 46806 9083
rect 46868 9042 46926 9166
rect 46988 9129 46998 9136
rect 46987 9083 46998 9129
rect 47168 9129 47178 9136
rect 47360 9129 47370 9136
rect 46988 9076 46998 9083
rect 47168 9083 47179 9129
rect 47359 9083 47370 9129
rect 47540 9129 47550 9136
rect 47168 9076 47178 9083
rect 47360 9076 47370 9083
rect 47540 9083 47551 9129
rect 47540 9076 47550 9083
rect 47612 9042 47670 9166
rect 47732 9129 47742 9136
rect 47731 9083 47742 9129
rect 47912 9129 47922 9136
rect 48104 9129 48114 9136
rect 47732 9076 47742 9083
rect 47912 9083 47923 9129
rect 48103 9083 48114 9129
rect 48284 9129 48294 9136
rect 47912 9076 47922 9083
rect 48104 9076 48114 9083
rect 48284 9083 48295 9129
rect 48284 9076 48294 9083
rect 48356 9042 48414 9166
rect 48476 9129 48486 9136
rect 48475 9083 48486 9129
rect 48656 9129 48666 9136
rect 48848 9129 48858 9136
rect 48476 9076 48486 9083
rect 48656 9083 48667 9129
rect 48847 9083 48858 9129
rect 49028 9129 49038 9136
rect 48656 9076 48666 9083
rect 48848 9076 48858 9083
rect 49028 9083 49039 9129
rect 49028 9076 49038 9083
rect 49100 9042 49158 9166
rect 49220 9129 49230 9136
rect 49219 9083 49230 9129
rect 49400 9129 49410 9136
rect 49592 9129 49602 9136
rect 49220 9076 49230 9083
rect 49400 9083 49411 9129
rect 49591 9083 49602 9129
rect 49772 9129 49782 9136
rect 49400 9076 49410 9083
rect 49592 9076 49602 9083
rect 49772 9083 49783 9129
rect 49772 9076 49782 9083
rect 49826 9042 49884 9166
rect 43930 9030 44001 9042
rect 43930 8654 43961 9030
rect 43995 8654 44001 9030
rect 43930 8642 44001 8654
rect 44213 9030 44373 9042
rect 44213 8654 44219 9030
rect 44253 8654 44333 9030
rect 44367 8654 44373 9030
rect 44213 8642 44373 8654
rect 44585 9030 44745 9042
rect 44585 8654 44591 9030
rect 44625 8654 44705 9030
rect 44739 8654 44745 9030
rect 44585 8642 44745 8654
rect 44957 9030 45117 9042
rect 44957 8654 44963 9030
rect 44997 8654 45077 9030
rect 45111 8654 45117 9030
rect 44957 8642 45117 8654
rect 45329 9030 45489 9042
rect 45329 8654 45335 9030
rect 45369 8654 45449 9030
rect 45483 8654 45489 9030
rect 45329 8642 45489 8654
rect 45701 9030 45861 9042
rect 45701 8654 45707 9030
rect 45741 8654 45821 9030
rect 45855 8654 45861 9030
rect 45701 8642 45861 8654
rect 46073 9030 46233 9042
rect 46073 8654 46079 9030
rect 46113 8654 46193 9030
rect 46227 8654 46233 9030
rect 46073 8642 46233 8654
rect 46445 9030 46605 9042
rect 46445 8654 46451 9030
rect 46485 8654 46565 9030
rect 46599 8654 46605 9030
rect 46445 8642 46605 8654
rect 46817 9030 46977 9042
rect 46817 8654 46823 9030
rect 46857 8654 46937 9030
rect 46971 8654 46977 9030
rect 46817 8642 46977 8654
rect 47189 9030 47349 9042
rect 47189 8654 47195 9030
rect 47229 8654 47309 9030
rect 47343 8654 47349 9030
rect 47189 8642 47349 8654
rect 47561 9030 47721 9042
rect 47561 8654 47567 9030
rect 47601 8654 47681 9030
rect 47715 8654 47721 9030
rect 47561 8642 47721 8654
rect 47933 9030 48093 9042
rect 47933 8654 47939 9030
rect 47973 8654 48053 9030
rect 48087 8654 48093 9030
rect 47933 8642 48093 8654
rect 48305 9030 48465 9042
rect 48305 8654 48311 9030
rect 48345 8654 48425 9030
rect 48459 8654 48465 9030
rect 48305 8642 48465 8654
rect 48677 9030 48837 9042
rect 48677 8654 48683 9030
rect 48717 8654 48797 9030
rect 48831 8654 48837 9030
rect 48677 8642 48837 8654
rect 49049 9030 49209 9042
rect 49049 8654 49055 9030
rect 49089 8654 49169 9030
rect 49203 8654 49209 9030
rect 49049 8642 49209 8654
rect 49421 9030 49581 9042
rect 49421 8654 49427 9030
rect 49461 8654 49541 9030
rect 49575 8654 49581 9030
rect 49421 8642 49581 8654
rect 49793 9030 49884 9042
rect 49793 8654 49799 9030
rect 49833 8654 49884 9030
rect 49793 8642 49884 8654
rect 43930 8406 43982 8642
rect 44010 8601 44136 8602
rect 44010 8596 44203 8601
rect 44010 8452 44022 8596
rect 44192 8555 44203 8596
rect 44192 8493 44202 8555
rect 44192 8452 44203 8493
rect 44010 8447 44203 8452
rect 44010 8446 44136 8447
rect 44258 8406 44328 8642
rect 44383 8596 44575 8601
rect 44383 8555 44394 8596
rect 44384 8493 44394 8555
rect 44383 8452 44394 8493
rect 44564 8555 44575 8596
rect 44564 8493 44574 8555
rect 44564 8452 44575 8493
rect 44383 8447 44575 8452
rect 44630 8406 44700 8642
rect 44755 8596 44947 8601
rect 44755 8555 44766 8596
rect 44756 8493 44766 8555
rect 44755 8452 44766 8493
rect 44936 8555 44947 8596
rect 44936 8493 44946 8555
rect 44936 8452 44947 8493
rect 44755 8447 44947 8452
rect 45002 8406 45072 8642
rect 45127 8596 45319 8601
rect 45127 8555 45138 8596
rect 45128 8493 45138 8555
rect 45127 8452 45138 8493
rect 45308 8555 45319 8596
rect 45308 8493 45318 8555
rect 45308 8452 45319 8493
rect 45127 8447 45319 8452
rect 45374 8406 45444 8642
rect 45499 8596 45691 8601
rect 45499 8555 45510 8596
rect 45500 8493 45510 8555
rect 45499 8452 45510 8493
rect 45680 8555 45691 8596
rect 45680 8493 45690 8555
rect 45680 8452 45691 8493
rect 45499 8447 45691 8452
rect 45746 8406 45816 8642
rect 45871 8596 46063 8601
rect 45871 8555 45882 8596
rect 45872 8493 45882 8555
rect 45871 8452 45882 8493
rect 46052 8555 46063 8596
rect 46052 8493 46062 8555
rect 46052 8452 46063 8493
rect 45871 8447 46063 8452
rect 46118 8406 46188 8642
rect 46243 8596 46435 8601
rect 46243 8555 46254 8596
rect 46244 8493 46254 8555
rect 46243 8452 46254 8493
rect 46424 8555 46435 8596
rect 46424 8493 46434 8555
rect 46424 8452 46435 8493
rect 46243 8447 46435 8452
rect 46490 8406 46560 8642
rect 46615 8596 46807 8601
rect 46615 8555 46626 8596
rect 46616 8493 46626 8555
rect 46615 8452 46626 8493
rect 46796 8555 46807 8596
rect 46796 8493 46806 8555
rect 46796 8452 46807 8493
rect 46615 8447 46807 8452
rect 46862 8406 46932 8642
rect 46987 8596 47179 8601
rect 46987 8555 46998 8596
rect 46988 8493 46998 8555
rect 46987 8452 46998 8493
rect 47168 8555 47179 8596
rect 47168 8493 47178 8555
rect 47168 8452 47179 8493
rect 46987 8447 47179 8452
rect 47234 8406 47304 8642
rect 47359 8596 47551 8601
rect 47359 8555 47370 8596
rect 47360 8493 47370 8555
rect 47359 8452 47370 8493
rect 47540 8555 47551 8596
rect 47540 8493 47550 8555
rect 47540 8452 47551 8493
rect 47359 8447 47551 8452
rect 47606 8406 47676 8642
rect 47731 8596 47923 8601
rect 47731 8555 47742 8596
rect 47732 8493 47742 8555
rect 47731 8452 47742 8493
rect 47912 8555 47923 8596
rect 47912 8493 47922 8555
rect 47912 8452 47923 8493
rect 47731 8447 47923 8452
rect 47978 8406 48048 8642
rect 48103 8596 48295 8601
rect 48103 8555 48114 8596
rect 48104 8493 48114 8555
rect 48103 8452 48114 8493
rect 48284 8555 48295 8596
rect 48284 8493 48294 8555
rect 48284 8452 48295 8493
rect 48103 8447 48295 8452
rect 48350 8406 48420 8642
rect 48475 8596 48667 8601
rect 48475 8555 48486 8596
rect 48476 8493 48486 8555
rect 48475 8452 48486 8493
rect 48656 8555 48667 8596
rect 48656 8493 48666 8555
rect 48656 8452 48667 8493
rect 48475 8447 48667 8452
rect 48722 8406 48792 8642
rect 48847 8596 49039 8601
rect 48847 8555 48858 8596
rect 48848 8493 48858 8555
rect 48847 8452 48858 8493
rect 49028 8555 49039 8596
rect 49028 8493 49038 8555
rect 49028 8452 49039 8493
rect 48847 8447 49039 8452
rect 49094 8406 49164 8642
rect 49219 8596 49411 8601
rect 49219 8555 49230 8596
rect 49220 8493 49230 8555
rect 49219 8452 49230 8493
rect 49400 8555 49411 8596
rect 49400 8493 49410 8555
rect 49400 8452 49411 8493
rect 49219 8447 49411 8452
rect 49466 8406 49536 8642
rect 49591 8596 49783 8601
rect 49591 8555 49602 8596
rect 49592 8493 49602 8555
rect 49591 8452 49602 8493
rect 49772 8555 49783 8596
rect 49772 8493 49782 8555
rect 49772 8452 49783 8493
rect 49591 8447 49783 8452
rect 49826 8406 49884 8642
rect 43930 8394 44001 8406
rect 43930 8018 43961 8394
rect 43995 8018 44001 8394
rect 43930 8006 44001 8018
rect 44213 8394 44373 8406
rect 44213 8018 44219 8394
rect 44253 8018 44333 8394
rect 44367 8018 44373 8394
rect 44213 8006 44373 8018
rect 44585 8394 44745 8406
rect 44585 8018 44591 8394
rect 44625 8018 44705 8394
rect 44739 8018 44745 8394
rect 44585 8006 44745 8018
rect 44957 8394 45117 8406
rect 44957 8018 44963 8394
rect 44997 8018 45077 8394
rect 45111 8018 45117 8394
rect 44957 8006 45117 8018
rect 45329 8394 45489 8406
rect 45329 8018 45335 8394
rect 45369 8018 45449 8394
rect 45483 8018 45489 8394
rect 45329 8006 45489 8018
rect 45701 8394 45861 8406
rect 45701 8018 45707 8394
rect 45741 8018 45821 8394
rect 45855 8018 45861 8394
rect 45701 8006 45861 8018
rect 46073 8394 46233 8406
rect 46073 8018 46079 8394
rect 46113 8018 46193 8394
rect 46227 8018 46233 8394
rect 46073 8006 46233 8018
rect 46445 8394 46605 8406
rect 46445 8018 46451 8394
rect 46485 8018 46565 8394
rect 46599 8018 46605 8394
rect 46445 8006 46605 8018
rect 46817 8394 46977 8406
rect 46817 8018 46823 8394
rect 46857 8018 46937 8394
rect 46971 8018 46977 8394
rect 46817 8006 46977 8018
rect 47189 8394 47349 8406
rect 47189 8018 47195 8394
rect 47229 8018 47309 8394
rect 47343 8018 47349 8394
rect 47189 8006 47349 8018
rect 47561 8394 47721 8406
rect 47561 8018 47567 8394
rect 47601 8018 47681 8394
rect 47715 8018 47721 8394
rect 47561 8006 47721 8018
rect 47933 8394 48093 8406
rect 47933 8018 47939 8394
rect 47973 8018 48053 8394
rect 48087 8018 48093 8394
rect 47933 8006 48093 8018
rect 48305 8394 48465 8406
rect 48305 8018 48311 8394
rect 48345 8018 48425 8394
rect 48459 8018 48465 8394
rect 48305 8006 48465 8018
rect 48677 8394 48837 8406
rect 48677 8018 48683 8394
rect 48717 8018 48797 8394
rect 48831 8018 48837 8394
rect 48677 8006 48837 8018
rect 49049 8394 49209 8406
rect 49049 8018 49055 8394
rect 49089 8018 49169 8394
rect 49203 8018 49209 8394
rect 49049 8006 49209 8018
rect 49421 8394 49581 8406
rect 49421 8018 49427 8394
rect 49461 8018 49541 8394
rect 49575 8018 49581 8394
rect 49421 8006 49581 8018
rect 49793 8394 49884 8406
rect 49793 8018 49799 8394
rect 49833 8018 49884 8394
rect 49793 8006 49884 8018
rect 43930 7770 43982 8006
rect 44010 7965 44152 7966
rect 44010 7960 44203 7965
rect 44010 7816 44022 7960
rect 44192 7919 44203 7960
rect 44192 7857 44202 7919
rect 44192 7816 44203 7857
rect 44010 7811 44203 7816
rect 44010 7810 44152 7811
rect 44258 7770 44328 8006
rect 44383 7960 44575 7965
rect 44383 7919 44394 7960
rect 44384 7857 44394 7919
rect 44383 7816 44394 7857
rect 44564 7919 44575 7960
rect 44564 7857 44574 7919
rect 44564 7816 44575 7857
rect 44383 7811 44575 7816
rect 44630 7770 44700 8006
rect 44755 7960 44947 7965
rect 44755 7919 44766 7960
rect 44756 7857 44766 7919
rect 44755 7816 44766 7857
rect 44936 7919 44947 7960
rect 44936 7857 44946 7919
rect 44936 7816 44947 7857
rect 44755 7811 44947 7816
rect 45002 7770 45072 8006
rect 45127 7960 45319 7965
rect 45127 7919 45138 7960
rect 45128 7857 45138 7919
rect 45127 7816 45138 7857
rect 45308 7919 45319 7960
rect 45308 7857 45318 7919
rect 45308 7816 45319 7857
rect 45127 7811 45319 7816
rect 45374 7770 45444 8006
rect 45499 7960 45691 7965
rect 45499 7919 45510 7960
rect 45500 7857 45510 7919
rect 45499 7816 45510 7857
rect 45680 7919 45691 7960
rect 45680 7857 45690 7919
rect 45680 7816 45691 7857
rect 45499 7811 45691 7816
rect 45746 7770 45816 8006
rect 45871 7960 46063 7965
rect 45871 7919 45882 7960
rect 45872 7857 45882 7919
rect 45871 7816 45882 7857
rect 46052 7919 46063 7960
rect 46052 7857 46062 7919
rect 46052 7816 46063 7857
rect 45871 7811 46063 7816
rect 46118 7770 46188 8006
rect 46243 7960 46435 7965
rect 46243 7919 46254 7960
rect 46244 7857 46254 7919
rect 46243 7816 46254 7857
rect 46424 7919 46435 7960
rect 46424 7857 46434 7919
rect 46424 7816 46435 7857
rect 46243 7811 46435 7816
rect 46490 7770 46560 8006
rect 46615 7960 46807 7965
rect 46615 7919 46626 7960
rect 46616 7857 46626 7919
rect 46615 7816 46626 7857
rect 46796 7919 46807 7960
rect 46796 7857 46806 7919
rect 46796 7816 46807 7857
rect 46615 7811 46807 7816
rect 46862 7770 46932 8006
rect 46987 7960 47179 7965
rect 46987 7919 46998 7960
rect 46988 7857 46998 7919
rect 46987 7816 46998 7857
rect 47168 7919 47179 7960
rect 47168 7857 47178 7919
rect 47168 7816 47179 7857
rect 46987 7811 47179 7816
rect 47234 7770 47304 8006
rect 47359 7960 47551 7965
rect 47359 7919 47370 7960
rect 47360 7857 47370 7919
rect 47359 7816 47370 7857
rect 47540 7919 47551 7960
rect 47540 7857 47550 7919
rect 47540 7816 47551 7857
rect 47359 7811 47551 7816
rect 47606 7770 47676 8006
rect 47731 7960 47923 7965
rect 47731 7919 47742 7960
rect 47732 7857 47742 7919
rect 47731 7816 47742 7857
rect 47912 7919 47923 7960
rect 47912 7857 47922 7919
rect 47912 7816 47923 7857
rect 47731 7811 47923 7816
rect 47978 7770 48048 8006
rect 48103 7960 48295 7965
rect 48103 7919 48114 7960
rect 48104 7857 48114 7919
rect 48103 7816 48114 7857
rect 48284 7919 48295 7960
rect 48284 7857 48294 7919
rect 48284 7816 48295 7857
rect 48103 7811 48295 7816
rect 48350 7770 48420 8006
rect 48475 7960 48667 7965
rect 48475 7919 48486 7960
rect 48476 7857 48486 7919
rect 48475 7816 48486 7857
rect 48656 7919 48667 7960
rect 48656 7857 48666 7919
rect 48656 7816 48667 7857
rect 48475 7811 48667 7816
rect 48722 7770 48792 8006
rect 48847 7960 49039 7965
rect 48847 7919 48858 7960
rect 48848 7857 48858 7919
rect 48847 7816 48858 7857
rect 49028 7919 49039 7960
rect 49028 7857 49038 7919
rect 49028 7816 49039 7857
rect 48847 7811 49039 7816
rect 49094 7770 49164 8006
rect 49219 7960 49411 7965
rect 49219 7919 49230 7960
rect 49220 7857 49230 7919
rect 49219 7816 49230 7857
rect 49400 7919 49411 7960
rect 49400 7857 49410 7919
rect 49400 7816 49411 7857
rect 49219 7811 49411 7816
rect 49466 7770 49536 8006
rect 49591 7960 49783 7965
rect 49591 7919 49602 7960
rect 49592 7857 49602 7919
rect 49591 7816 49602 7857
rect 49772 7919 49783 7960
rect 49772 7857 49782 7919
rect 49772 7816 49783 7857
rect 49591 7811 49783 7816
rect 49826 7770 49884 8006
rect 43930 7758 44001 7770
rect 43930 7382 43961 7758
rect 43995 7382 44001 7758
rect 43930 7370 44001 7382
rect 44213 7758 44373 7770
rect 44213 7382 44219 7758
rect 44253 7382 44333 7758
rect 44367 7382 44373 7758
rect 44213 7370 44373 7382
rect 44585 7758 44745 7770
rect 44585 7382 44591 7758
rect 44625 7382 44705 7758
rect 44739 7382 44745 7758
rect 44585 7370 44745 7382
rect 44957 7758 45117 7770
rect 44957 7382 44963 7758
rect 44997 7382 45077 7758
rect 45111 7382 45117 7758
rect 44957 7370 45117 7382
rect 45329 7758 45489 7770
rect 45329 7382 45335 7758
rect 45369 7382 45449 7758
rect 45483 7382 45489 7758
rect 45329 7370 45489 7382
rect 45701 7758 45861 7770
rect 45701 7382 45707 7758
rect 45741 7382 45821 7758
rect 45855 7382 45861 7758
rect 45701 7370 45861 7382
rect 46073 7758 46233 7770
rect 46073 7382 46079 7758
rect 46113 7382 46193 7758
rect 46227 7382 46233 7758
rect 46073 7370 46233 7382
rect 46445 7758 46605 7770
rect 46445 7382 46451 7758
rect 46485 7382 46565 7758
rect 46599 7382 46605 7758
rect 46445 7370 46605 7382
rect 46817 7758 46977 7770
rect 46817 7382 46823 7758
rect 46857 7382 46937 7758
rect 46971 7382 46977 7758
rect 46817 7370 46977 7382
rect 47189 7758 47349 7770
rect 47189 7382 47195 7758
rect 47229 7382 47309 7758
rect 47343 7382 47349 7758
rect 47189 7370 47349 7382
rect 47561 7758 47721 7770
rect 47561 7382 47567 7758
rect 47601 7382 47681 7758
rect 47715 7382 47721 7758
rect 47561 7370 47721 7382
rect 47933 7758 48093 7770
rect 47933 7382 47939 7758
rect 47973 7382 48053 7758
rect 48087 7382 48093 7758
rect 47933 7370 48093 7382
rect 48305 7758 48465 7770
rect 48305 7382 48311 7758
rect 48345 7382 48425 7758
rect 48459 7382 48465 7758
rect 48305 7370 48465 7382
rect 48677 7758 48837 7770
rect 48677 7382 48683 7758
rect 48717 7382 48797 7758
rect 48831 7382 48837 7758
rect 48677 7370 48837 7382
rect 49049 7758 49209 7770
rect 49049 7382 49055 7758
rect 49089 7382 49169 7758
rect 49203 7382 49209 7758
rect 49049 7370 49209 7382
rect 49421 7758 49581 7770
rect 49421 7382 49427 7758
rect 49461 7382 49541 7758
rect 49575 7382 49581 7758
rect 49421 7370 49581 7382
rect 49793 7758 49884 7770
rect 49793 7382 49799 7758
rect 49833 7382 49884 7758
rect 49793 7370 49884 7382
rect 43268 7329 43278 7336
rect 43267 7283 43278 7329
rect 43448 7329 43458 7336
rect 43640 7329 43650 7336
rect 43268 7276 43278 7283
rect 43448 7283 43459 7329
rect 43639 7283 43650 7329
rect 43448 7276 43458 7283
rect 43640 7276 43650 7283
rect 43820 7276 43892 7336
rect 44008 7276 44022 7336
rect 44192 7329 44202 7336
rect 44192 7283 44203 7329
rect 44192 7276 44202 7283
rect 38684 6964 43206 7028
rect 44258 6968 44328 7370
rect 44384 7329 44394 7336
rect 44383 7283 44394 7329
rect 44564 7329 44574 7336
rect 44756 7329 44766 7336
rect 44384 7276 44394 7283
rect 44564 7283 44575 7329
rect 44755 7283 44766 7329
rect 44936 7329 44946 7336
rect 44564 7276 44574 7283
rect 44756 7276 44766 7283
rect 44936 7283 44947 7329
rect 44936 7276 44946 7283
rect 45002 6968 45072 7370
rect 45128 7329 45138 7336
rect 45127 7283 45138 7329
rect 45308 7329 45318 7336
rect 45500 7329 45510 7336
rect 45128 7276 45138 7283
rect 45308 7283 45319 7329
rect 45499 7283 45510 7329
rect 45680 7329 45690 7336
rect 45308 7276 45318 7283
rect 45500 7276 45510 7283
rect 45680 7283 45691 7329
rect 45680 7276 45690 7283
rect 45746 6968 45816 7370
rect 45872 7329 45882 7336
rect 45871 7283 45882 7329
rect 46052 7329 46062 7336
rect 46244 7329 46254 7336
rect 45872 7276 45882 7283
rect 46052 7283 46063 7329
rect 46243 7283 46254 7329
rect 46424 7329 46434 7336
rect 46052 7276 46062 7283
rect 46244 7276 46254 7283
rect 46424 7283 46435 7329
rect 46424 7276 46434 7283
rect 46490 6968 46560 7370
rect 46616 7329 46626 7336
rect 46615 7283 46626 7329
rect 46796 7329 46806 7336
rect 46988 7329 46998 7336
rect 46616 7276 46626 7283
rect 46796 7283 46807 7329
rect 46987 7283 46998 7329
rect 47168 7329 47178 7336
rect 46796 7276 46806 7283
rect 46988 7276 46998 7283
rect 47168 7283 47179 7329
rect 47168 7276 47178 7283
rect 47234 6968 47304 7370
rect 47360 7329 47370 7336
rect 47359 7283 47370 7329
rect 47540 7329 47550 7336
rect 47732 7329 47742 7336
rect 47360 7276 47370 7283
rect 47540 7283 47551 7329
rect 47731 7283 47742 7329
rect 47912 7329 47922 7336
rect 47540 7276 47550 7283
rect 47732 7276 47742 7283
rect 47912 7283 47923 7329
rect 47912 7276 47922 7283
rect 47978 6968 48048 7370
rect 48104 7329 48114 7336
rect 48103 7283 48114 7329
rect 48284 7329 48294 7336
rect 48476 7329 48486 7336
rect 48104 7276 48114 7283
rect 48284 7283 48295 7329
rect 48475 7283 48486 7329
rect 48656 7329 48666 7336
rect 48284 7276 48294 7283
rect 48476 7276 48486 7283
rect 48656 7283 48667 7329
rect 48656 7276 48666 7283
rect 48722 6968 48792 7370
rect 48848 7329 48858 7336
rect 48847 7283 48858 7329
rect 49028 7329 49038 7336
rect 49220 7329 49230 7336
rect 48848 7276 48858 7283
rect 49028 7283 49039 7329
rect 49219 7283 49230 7329
rect 49400 7329 49410 7336
rect 49028 7276 49038 7283
rect 49220 7276 49230 7283
rect 49400 7283 49411 7329
rect 49400 7276 49410 7283
rect 49466 6968 49536 7370
rect 49592 7329 49602 7336
rect 49591 7283 49602 7329
rect 49772 7329 49782 7336
rect 49592 7276 49602 7283
rect 49772 7283 49783 7329
rect 49772 7276 49782 7283
rect 39444 6860 39498 6964
rect 39840 6860 39910 6964
rect 40172 6860 40230 6964
rect 40584 6860 40654 6964
rect 40916 6860 40974 6964
rect 41328 6860 41398 6964
rect 41660 6860 41718 6964
rect 42072 6860 42142 6964
rect 42392 6860 42446 6964
rect 39444 6854 39550 6860
rect 39444 6784 39468 6854
rect 39538 6784 39550 6854
rect 39444 6778 39550 6784
rect 39828 6854 39922 6860
rect 39828 6784 39840 6854
rect 39910 6784 39922 6854
rect 39828 6778 39922 6784
rect 40172 6854 40294 6860
rect 40172 6784 40212 6854
rect 40282 6784 40294 6854
rect 40172 6778 40294 6784
rect 40572 6854 40666 6860
rect 40572 6784 40584 6854
rect 40654 6784 40666 6854
rect 40572 6778 40666 6784
rect 40916 6854 41038 6860
rect 40916 6784 40956 6854
rect 41026 6784 41038 6854
rect 40916 6778 41038 6784
rect 41316 6854 41410 6860
rect 41316 6784 41328 6854
rect 41398 6784 41410 6854
rect 41316 6778 41410 6784
rect 41660 6854 41782 6860
rect 41660 6784 41700 6854
rect 41770 6784 41782 6854
rect 41660 6778 41782 6784
rect 42060 6854 42154 6860
rect 42060 6784 42072 6854
rect 42142 6784 42154 6854
rect 42060 6778 42154 6784
rect 42322 6854 42446 6860
rect 42322 6784 42334 6854
rect 42404 6784 42446 6854
rect 42322 6778 42446 6784
rect 39444 6654 39498 6778
rect 39548 6741 39558 6750
rect 39547 6695 39558 6741
rect 39728 6741 39738 6750
rect 39920 6741 39930 6750
rect 39548 6686 39558 6695
rect 39728 6695 39739 6741
rect 39919 6695 39930 6741
rect 40100 6741 40110 6750
rect 39728 6686 39738 6695
rect 39920 6686 39930 6695
rect 40100 6695 40111 6741
rect 40100 6686 40110 6695
rect 40172 6654 40230 6778
rect 40292 6741 40302 6750
rect 40291 6695 40302 6741
rect 40472 6741 40482 6750
rect 40664 6741 40674 6750
rect 40292 6686 40302 6695
rect 40472 6695 40483 6741
rect 40663 6695 40674 6741
rect 40844 6741 40854 6750
rect 40472 6686 40482 6695
rect 40664 6686 40674 6695
rect 40844 6695 40855 6741
rect 40844 6686 40854 6695
rect 40916 6654 40974 6778
rect 41036 6741 41046 6750
rect 41035 6695 41046 6741
rect 41216 6741 41226 6750
rect 41408 6741 41418 6750
rect 41036 6686 41046 6695
rect 41216 6695 41227 6741
rect 41407 6695 41418 6741
rect 41588 6741 41598 6750
rect 41216 6686 41226 6695
rect 41408 6686 41418 6695
rect 41588 6695 41599 6741
rect 41588 6686 41598 6695
rect 41660 6654 41718 6778
rect 41780 6741 41790 6750
rect 41779 6695 41790 6741
rect 41960 6741 41970 6750
rect 42152 6741 42162 6750
rect 41780 6686 41790 6695
rect 41960 6695 41971 6741
rect 42151 6695 42162 6741
rect 42332 6741 42342 6750
rect 41960 6686 41970 6695
rect 42152 6686 42162 6695
rect 42332 6695 42343 6741
rect 42332 6686 42342 6695
rect 42392 6654 42446 6778
rect 44144 6696 44154 6968
rect 44436 6696 44446 6968
rect 44888 6696 44898 6968
rect 45180 6696 45190 6968
rect 45632 6696 45642 6968
rect 45924 6696 45934 6968
rect 46376 6696 46386 6968
rect 46668 6696 46678 6968
rect 47120 6696 47130 6968
rect 47412 6696 47422 6968
rect 47864 6696 47874 6968
rect 48156 6696 48166 6968
rect 48608 6696 48618 6968
rect 48900 6696 48910 6968
rect 49352 6696 49362 6968
rect 49644 6696 49654 6968
rect 39444 6642 39537 6654
rect 39444 5866 39497 6642
rect 39531 5866 39537 6642
rect 39444 5854 39537 5866
rect 39749 6642 39909 6654
rect 39749 5866 39755 6642
rect 39789 5866 39869 6642
rect 39903 5866 39909 6642
rect 39749 5854 39909 5866
rect 40121 6642 40281 6654
rect 40121 5866 40127 6642
rect 40161 5866 40241 6642
rect 40275 5866 40281 6642
rect 40121 5854 40281 5866
rect 40493 6642 40653 6654
rect 40493 5866 40499 6642
rect 40533 5866 40613 6642
rect 40647 5866 40653 6642
rect 40493 5854 40653 5866
rect 40865 6642 41025 6654
rect 40865 5866 40871 6642
rect 40905 5866 40985 6642
rect 41019 5866 41025 6642
rect 40865 5854 41025 5866
rect 41237 6642 41397 6654
rect 41237 5866 41243 6642
rect 41277 5866 41357 6642
rect 41391 5866 41397 6642
rect 41237 5854 41397 5866
rect 41609 6642 41769 6654
rect 41609 5866 41615 6642
rect 41649 5866 41729 6642
rect 41763 5866 41769 6642
rect 41609 5854 41769 5866
rect 41981 6642 42141 6654
rect 41981 5866 41987 6642
rect 42021 5866 42101 6642
rect 42135 5866 42141 6642
rect 41981 5854 42141 5866
rect 42353 6642 42446 6654
rect 42353 5866 42359 6642
rect 42393 5866 42446 6642
rect 42353 5854 42446 5866
rect 39444 5618 39492 5854
rect 39547 5808 39739 5813
rect 39547 5767 39558 5808
rect 39548 5705 39558 5767
rect 39547 5664 39558 5705
rect 39728 5767 39739 5808
rect 39728 5705 39738 5767
rect 39728 5664 39739 5705
rect 39547 5659 39739 5664
rect 39794 5618 39864 5854
rect 39919 5808 40111 5813
rect 39919 5767 39930 5808
rect 39920 5705 39930 5767
rect 39919 5664 39930 5705
rect 40100 5767 40111 5808
rect 40100 5705 40110 5767
rect 40100 5664 40111 5705
rect 39919 5659 40111 5664
rect 40166 5618 40236 5854
rect 40291 5808 40483 5813
rect 40291 5767 40302 5808
rect 40292 5705 40302 5767
rect 40291 5664 40302 5705
rect 40472 5767 40483 5808
rect 40472 5705 40482 5767
rect 40472 5664 40483 5705
rect 40291 5659 40483 5664
rect 40538 5618 40608 5854
rect 40663 5808 40855 5813
rect 40663 5767 40674 5808
rect 40664 5705 40674 5767
rect 40663 5664 40674 5705
rect 40844 5767 40855 5808
rect 40844 5705 40854 5767
rect 40844 5664 40855 5705
rect 40663 5659 40855 5664
rect 40910 5618 40980 5854
rect 41035 5808 41227 5813
rect 41035 5767 41046 5808
rect 41036 5705 41046 5767
rect 41035 5664 41046 5705
rect 41216 5767 41227 5808
rect 41216 5705 41226 5767
rect 41216 5664 41227 5705
rect 41035 5659 41227 5664
rect 41282 5618 41352 5854
rect 41407 5808 41599 5813
rect 41407 5767 41418 5808
rect 41408 5705 41418 5767
rect 41407 5664 41418 5705
rect 41588 5767 41599 5808
rect 41588 5705 41598 5767
rect 41588 5664 41599 5705
rect 41407 5659 41599 5664
rect 41654 5618 41724 5854
rect 41779 5808 41971 5813
rect 41779 5767 41790 5808
rect 41780 5705 41790 5767
rect 41779 5664 41790 5705
rect 41960 5767 41971 5808
rect 41960 5705 41970 5767
rect 41960 5664 41971 5705
rect 41779 5659 41971 5664
rect 42026 5618 42096 5854
rect 42151 5808 42343 5813
rect 42151 5767 42162 5808
rect 42152 5705 42162 5767
rect 42151 5664 42162 5705
rect 42332 5767 42343 5808
rect 42332 5705 42342 5767
rect 42332 5664 42343 5705
rect 42151 5659 42343 5664
rect 42392 5618 42446 5854
rect 39444 5606 39537 5618
rect 39444 4830 39497 5606
rect 39531 4830 39537 5606
rect 39444 4818 39537 4830
rect 39749 5606 39909 5618
rect 39749 4830 39755 5606
rect 39789 4830 39869 5606
rect 39903 4830 39909 5606
rect 39749 4818 39909 4830
rect 40121 5606 40281 5618
rect 40121 4830 40127 5606
rect 40161 4830 40241 5606
rect 40275 4830 40281 5606
rect 40121 4818 40281 4830
rect 40493 5606 40653 5618
rect 40493 4830 40499 5606
rect 40533 4830 40613 5606
rect 40647 4830 40653 5606
rect 40493 4818 40653 4830
rect 40865 5606 41025 5618
rect 40865 4830 40871 5606
rect 40905 4830 40985 5606
rect 41019 4830 41025 5606
rect 40865 4818 41025 4830
rect 41237 5606 41397 5618
rect 41237 4830 41243 5606
rect 41277 4830 41357 5606
rect 41391 4830 41397 5606
rect 41237 4818 41397 4830
rect 41609 5606 41769 5618
rect 41609 4830 41615 5606
rect 41649 4830 41729 5606
rect 41763 4830 41769 5606
rect 41609 4818 41769 4830
rect 41981 5606 42141 5618
rect 41981 4830 41987 5606
rect 42021 4830 42101 5606
rect 42135 4830 42141 5606
rect 41981 4818 42141 4830
rect 42353 5606 42446 5618
rect 42353 4830 42359 5606
rect 42393 4830 42446 5606
rect 43026 4980 43036 5252
rect 43318 4980 43328 5252
rect 42353 4818 42446 4830
rect 39444 4582 39492 4818
rect 39547 4772 39739 4777
rect 39547 4731 39558 4772
rect 39548 4669 39558 4731
rect 39547 4628 39558 4669
rect 39728 4731 39739 4772
rect 39728 4669 39738 4731
rect 39728 4628 39739 4669
rect 39547 4623 39739 4628
rect 39794 4582 39864 4818
rect 39919 4772 40111 4777
rect 39919 4731 39930 4772
rect 39920 4669 39930 4731
rect 39919 4628 39930 4669
rect 40100 4731 40111 4772
rect 40100 4669 40110 4731
rect 40100 4628 40111 4669
rect 39919 4623 40111 4628
rect 40166 4582 40236 4818
rect 40291 4772 40483 4777
rect 40291 4731 40302 4772
rect 40292 4669 40302 4731
rect 40291 4628 40302 4669
rect 40472 4731 40483 4772
rect 40472 4669 40482 4731
rect 40472 4628 40483 4669
rect 40291 4623 40483 4628
rect 40538 4582 40608 4818
rect 40663 4772 40855 4777
rect 40663 4731 40674 4772
rect 40664 4669 40674 4731
rect 40663 4628 40674 4669
rect 40844 4731 40855 4772
rect 40844 4669 40854 4731
rect 40844 4628 40855 4669
rect 40663 4623 40855 4628
rect 40910 4582 40980 4818
rect 41035 4772 41227 4777
rect 41035 4731 41046 4772
rect 41036 4669 41046 4731
rect 41035 4628 41046 4669
rect 41216 4731 41227 4772
rect 41216 4669 41226 4731
rect 41216 4628 41227 4669
rect 41035 4623 41227 4628
rect 41282 4582 41352 4818
rect 41407 4772 41599 4777
rect 41407 4731 41418 4772
rect 41408 4669 41418 4731
rect 41407 4628 41418 4669
rect 41588 4731 41599 4772
rect 41588 4669 41598 4731
rect 41588 4628 41599 4669
rect 41407 4623 41599 4628
rect 41654 4582 41724 4818
rect 41779 4772 41971 4777
rect 41779 4731 41790 4772
rect 41780 4669 41790 4731
rect 41779 4628 41790 4669
rect 41960 4731 41971 4772
rect 41960 4669 41970 4731
rect 41960 4628 41971 4669
rect 41779 4623 41971 4628
rect 42026 4582 42096 4818
rect 42151 4772 42343 4777
rect 42151 4731 42162 4772
rect 42152 4669 42162 4731
rect 42151 4628 42162 4669
rect 42332 4731 42343 4772
rect 42332 4669 42342 4731
rect 42332 4628 42343 4669
rect 42151 4623 42343 4628
rect 42392 4582 42446 4818
rect 39444 4570 39537 4582
rect 39444 3794 39497 4570
rect 39531 3794 39537 4570
rect 39444 3782 39537 3794
rect 39749 4570 39909 4582
rect 39749 3794 39755 4570
rect 39789 3794 39869 4570
rect 39903 3794 39909 4570
rect 39749 3782 39909 3794
rect 40121 4570 40281 4582
rect 40121 3794 40127 4570
rect 40161 3794 40241 4570
rect 40275 3794 40281 4570
rect 40121 3782 40281 3794
rect 40493 4570 40653 4582
rect 40493 3794 40499 4570
rect 40533 3794 40613 4570
rect 40647 3794 40653 4570
rect 40493 3782 40653 3794
rect 40865 4570 41025 4582
rect 40865 3794 40871 4570
rect 40905 3794 40985 4570
rect 41019 3794 41025 4570
rect 40865 3782 41025 3794
rect 41237 4570 41397 4582
rect 41237 3794 41243 4570
rect 41277 3794 41357 4570
rect 41391 3794 41397 4570
rect 41237 3782 41397 3794
rect 41609 4570 41769 4582
rect 41609 3794 41615 4570
rect 41649 3794 41729 4570
rect 41763 3794 41769 4570
rect 41609 3782 41769 3794
rect 41981 4570 42141 4582
rect 41981 3794 41987 4570
rect 42021 3794 42101 4570
rect 42135 3794 42141 4570
rect 41981 3782 42141 3794
rect 42353 4570 42446 4582
rect 42353 3794 42359 4570
rect 42393 3794 42446 4570
rect 43138 4775 43210 4980
rect 43138 4378 43155 4775
rect 43193 4378 43210 4775
rect 43450 4664 43460 4712
rect 43278 4658 43460 4664
rect 43278 4596 43290 4658
rect 43354 4596 43460 4658
rect 43278 4590 43460 4596
rect 43450 4548 43460 4590
rect 43612 4548 43622 4712
rect 43138 4360 43210 4378
rect 43450 4264 43460 4312
rect 43278 4258 43460 4264
rect 43278 4196 43290 4258
rect 43354 4196 43460 4258
rect 43278 4190 43460 4196
rect 43450 4148 43460 4190
rect 43612 4148 43622 4312
rect 43450 3864 43460 3912
rect 43278 3858 43460 3864
rect 42353 3782 42446 3794
rect 39444 3546 39492 3782
rect 39547 3736 39739 3741
rect 39547 3695 39558 3736
rect 39548 3633 39558 3695
rect 39547 3592 39558 3633
rect 39728 3695 39739 3736
rect 39728 3633 39738 3695
rect 39728 3592 39739 3633
rect 39547 3587 39739 3592
rect 39794 3546 39864 3782
rect 39919 3736 40111 3741
rect 39919 3695 39930 3736
rect 39920 3633 39930 3695
rect 39919 3592 39930 3633
rect 40100 3695 40111 3736
rect 40100 3633 40110 3695
rect 40100 3592 40111 3633
rect 39919 3587 40111 3592
rect 40166 3546 40236 3782
rect 40291 3736 40483 3741
rect 40291 3695 40302 3736
rect 40292 3633 40302 3695
rect 40291 3592 40302 3633
rect 40472 3695 40483 3736
rect 40472 3633 40482 3695
rect 40472 3592 40483 3633
rect 40291 3587 40483 3592
rect 40538 3546 40608 3782
rect 40663 3736 40855 3741
rect 40663 3695 40674 3736
rect 40664 3633 40674 3695
rect 40663 3592 40674 3633
rect 40844 3695 40855 3736
rect 40844 3633 40854 3695
rect 40844 3592 40855 3633
rect 40663 3587 40855 3592
rect 40910 3546 40980 3782
rect 41035 3736 41227 3741
rect 41035 3695 41046 3736
rect 41036 3633 41046 3695
rect 41035 3592 41046 3633
rect 41216 3695 41227 3736
rect 41216 3633 41226 3695
rect 41216 3592 41227 3633
rect 41035 3587 41227 3592
rect 41282 3546 41352 3782
rect 41407 3736 41599 3741
rect 41407 3695 41418 3736
rect 41408 3633 41418 3695
rect 41407 3592 41418 3633
rect 41588 3695 41599 3736
rect 41588 3633 41598 3695
rect 41588 3592 41599 3633
rect 41407 3587 41599 3592
rect 41654 3546 41724 3782
rect 41779 3736 41971 3741
rect 41779 3695 41790 3736
rect 41780 3633 41790 3695
rect 41779 3592 41790 3633
rect 41960 3695 41971 3736
rect 41960 3633 41970 3695
rect 41960 3592 41971 3633
rect 41779 3587 41971 3592
rect 42026 3546 42096 3782
rect 42151 3736 42343 3741
rect 42151 3695 42162 3736
rect 42152 3633 42162 3695
rect 42151 3592 42162 3633
rect 42332 3695 42343 3736
rect 42332 3633 42342 3695
rect 42332 3592 42343 3633
rect 42151 3587 42343 3592
rect 42392 3546 42446 3782
rect 39444 3534 39537 3546
rect 39444 2758 39497 3534
rect 39531 2758 39537 3534
rect 39444 2746 39537 2758
rect 39749 3534 39909 3546
rect 39749 2758 39755 3534
rect 39789 2758 39869 3534
rect 39903 2758 39909 3534
rect 39749 2746 39909 2758
rect 40121 3534 40281 3546
rect 40121 2758 40127 3534
rect 40161 2758 40241 3534
rect 40275 2758 40281 3534
rect 40121 2746 40281 2758
rect 40493 3534 40653 3546
rect 40493 2758 40499 3534
rect 40533 2758 40613 3534
rect 40647 2758 40653 3534
rect 40493 2746 40653 2758
rect 40865 3534 41025 3546
rect 40865 2758 40871 3534
rect 40905 2758 40985 3534
rect 41019 2758 41025 3534
rect 40865 2746 41025 2758
rect 41237 3534 41397 3546
rect 41237 2758 41243 3534
rect 41277 2758 41357 3534
rect 41391 2758 41397 3534
rect 41237 2746 41397 2758
rect 41609 3534 41769 3546
rect 41609 2758 41615 3534
rect 41649 2758 41729 3534
rect 41763 2758 41769 3534
rect 41609 2746 41769 2758
rect 41981 3534 42141 3546
rect 41981 2758 41987 3534
rect 42021 2758 42101 3534
rect 42135 2758 42141 3534
rect 41981 2746 42141 2758
rect 42353 3534 42446 3546
rect 42353 2758 42359 3534
rect 42393 2758 42446 3534
rect 43138 3784 43210 3800
rect 43278 3796 43290 3858
rect 43354 3796 43460 3858
rect 43278 3790 43460 3796
rect 43138 3387 43155 3784
rect 43193 3387 43210 3784
rect 43450 3748 43460 3790
rect 43612 3748 43622 3912
rect 43450 3464 43460 3512
rect 43278 3458 43460 3464
rect 43278 3396 43290 3458
rect 43354 3396 43460 3458
rect 43278 3390 43460 3396
rect 42353 2746 42446 2758
rect 39548 2705 39558 2710
rect 39547 2659 39558 2705
rect 39728 2705 39738 2710
rect 39548 2656 39558 2659
rect 39728 2659 39739 2705
rect 39728 2656 39738 2659
rect 39794 2062 39864 2746
rect 39920 2705 39930 2710
rect 39919 2659 39930 2705
rect 40100 2705 40110 2710
rect 40292 2705 40302 2710
rect 39920 2656 39930 2659
rect 40100 2659 40111 2705
rect 40291 2659 40302 2705
rect 40472 2705 40482 2710
rect 40100 2656 40110 2659
rect 40292 2656 40302 2659
rect 40472 2659 40483 2705
rect 40472 2656 40482 2659
rect 40538 2370 40608 2746
rect 40664 2705 40674 2710
rect 40663 2659 40674 2705
rect 40844 2705 40854 2710
rect 41036 2705 41046 2710
rect 40664 2656 40674 2659
rect 40844 2659 40855 2705
rect 41035 2659 41046 2705
rect 41216 2705 41226 2710
rect 40844 2656 40854 2659
rect 41036 2656 41046 2659
rect 41216 2659 41227 2705
rect 41216 2656 41226 2659
rect 41282 2370 41352 2746
rect 41408 2705 41418 2710
rect 41407 2659 41418 2705
rect 41588 2705 41598 2710
rect 41780 2705 41790 2710
rect 41408 2656 41418 2659
rect 41588 2659 41599 2705
rect 41779 2659 41790 2705
rect 41960 2705 41970 2710
rect 41588 2656 41598 2659
rect 41780 2656 41790 2659
rect 41960 2659 41971 2705
rect 41960 2656 41970 2659
rect 40528 2190 40538 2370
rect 41352 2190 41362 2370
rect 39546 2052 40112 2062
rect 39546 2006 39558 2052
rect 39547 2001 39558 2006
rect 39548 1996 39558 2001
rect 39728 2006 39930 2052
rect 39728 2001 39739 2006
rect 39728 1996 39738 2001
rect 39442 1969 39516 1970
rect 39794 1969 39864 2006
rect 39919 2001 39930 2006
rect 39920 1996 39930 2001
rect 40100 2006 40112 2052
rect 40292 2047 40302 2052
rect 40100 2001 40111 2006
rect 40291 2001 40302 2047
rect 40472 2047 40482 2052
rect 40100 1996 40110 2001
rect 40292 1996 40302 2001
rect 40472 2001 40483 2047
rect 40472 1996 40482 2001
rect 40166 1969 40236 1970
rect 40538 1969 40608 2190
rect 40664 2047 40674 2052
rect 40663 2001 40674 2047
rect 40844 2047 40854 2052
rect 41036 2047 41046 2052
rect 40664 1996 40674 2001
rect 40844 2001 40855 2047
rect 41035 2001 41046 2047
rect 41216 2047 41226 2052
rect 40844 1996 40854 2001
rect 41036 1996 41046 2001
rect 41216 2001 41227 2047
rect 41216 1996 41226 2001
rect 40910 1969 40980 1970
rect 41282 1969 41352 2190
rect 42026 2062 42096 2746
rect 42152 2705 42162 2710
rect 42151 2659 42162 2705
rect 42332 2705 42342 2710
rect 42152 2656 42162 2659
rect 42332 2659 42343 2705
rect 42332 2656 42342 2659
rect 42654 2514 42664 2786
rect 42946 2514 42956 2786
rect 41778 2052 42344 2062
rect 41408 2047 41418 2052
rect 41407 2001 41418 2047
rect 41588 2047 41598 2052
rect 41408 1996 41418 2001
rect 41588 2001 41599 2047
rect 41778 2006 41790 2052
rect 41779 2001 41790 2006
rect 41588 1996 41598 2001
rect 41780 1996 41790 2001
rect 41960 2006 42162 2052
rect 41960 2001 41971 2006
rect 41960 1996 41970 2001
rect 41654 1969 41724 1970
rect 42026 1969 42096 2006
rect 42151 2001 42162 2006
rect 42152 1996 42162 2001
rect 42332 2006 42344 2052
rect 42524 2047 42534 2052
rect 42332 2001 42343 2006
rect 42523 2001 42534 2047
rect 42704 2047 42714 2052
rect 42332 1996 42342 2001
rect 42524 1996 42534 2001
rect 42704 2001 42715 2047
rect 42704 1996 42714 2001
rect 42398 1969 42468 1970
rect 42770 1969 42840 2514
rect 43138 2440 43210 3387
rect 43450 3348 43460 3390
rect 43612 3348 43622 3512
rect 43398 2514 43408 2786
rect 43690 2514 43700 2786
rect 44142 2514 44152 2786
rect 44434 2514 44444 2786
rect 44886 2514 44896 2786
rect 45178 2514 45188 2786
rect 45630 2514 45640 2786
rect 45922 2514 45932 2786
rect 46374 2514 46384 2786
rect 46666 2514 46676 2786
rect 47118 2514 47128 2786
rect 47410 2514 47420 2786
rect 47862 2514 47872 2786
rect 48154 2514 48164 2786
rect 43034 2190 43044 2440
rect 43294 2190 43304 2440
rect 42896 2047 42906 2052
rect 42895 2001 42906 2047
rect 43076 2047 43086 2052
rect 43268 2047 43278 2052
rect 42896 1996 42906 2001
rect 43076 2001 43087 2047
rect 43267 2001 43278 2047
rect 43448 2047 43458 2052
rect 43076 1996 43086 2001
rect 43268 1996 43278 2001
rect 43448 2001 43459 2047
rect 43448 1996 43458 2001
rect 43142 1969 43212 1970
rect 43514 1969 43584 2514
rect 43640 2047 43650 2052
rect 43639 2001 43650 2047
rect 43820 2047 43830 2052
rect 44012 2047 44022 2052
rect 43640 1996 43650 2001
rect 43820 2001 43831 2047
rect 44011 2001 44022 2047
rect 44192 2047 44202 2052
rect 43820 1996 43830 2001
rect 44012 1996 44022 2001
rect 44192 2001 44203 2047
rect 44192 1996 44202 2001
rect 43886 1969 43956 1970
rect 44258 1969 44328 2514
rect 44384 2047 44394 2052
rect 44383 2001 44394 2047
rect 44564 2047 44574 2052
rect 44756 2047 44766 2052
rect 44384 1996 44394 2001
rect 44564 2001 44575 2047
rect 44755 2001 44766 2047
rect 44936 2047 44946 2052
rect 44564 1996 44574 2001
rect 44756 1996 44766 2001
rect 44936 2001 44947 2047
rect 44936 1996 44946 2001
rect 44630 1969 44700 1970
rect 45002 1969 45072 2514
rect 45128 2047 45138 2052
rect 45127 2001 45138 2047
rect 45308 2047 45318 2052
rect 45500 2047 45510 2052
rect 45128 1996 45138 2001
rect 45308 2001 45319 2047
rect 45499 2001 45510 2047
rect 45680 2047 45690 2052
rect 45308 1996 45318 2001
rect 45500 1996 45510 2001
rect 45680 2001 45691 2047
rect 45680 1996 45690 2001
rect 45374 1969 45444 1970
rect 45746 1969 45816 2514
rect 45872 2047 45882 2052
rect 45871 2001 45882 2047
rect 46052 2047 46062 2052
rect 46244 2047 46254 2052
rect 45872 1996 45882 2001
rect 46052 2001 46063 2047
rect 46243 2001 46254 2047
rect 46424 2047 46434 2052
rect 46052 1996 46062 2001
rect 46244 1996 46254 2001
rect 46424 2001 46435 2047
rect 46424 1996 46434 2001
rect 46118 1969 46188 1970
rect 46490 1969 46560 2514
rect 46616 2047 46626 2052
rect 46615 2001 46626 2047
rect 46796 2047 46806 2052
rect 46988 2047 46998 2052
rect 46616 1996 46626 2001
rect 46796 2001 46807 2047
rect 46987 2001 46998 2047
rect 47168 2047 47178 2052
rect 46796 1996 46806 2001
rect 46988 1996 46998 2001
rect 47168 2001 47179 2047
rect 47168 1996 47178 2001
rect 46862 1969 46932 1970
rect 47234 1969 47304 2514
rect 47360 2047 47370 2052
rect 47359 2001 47370 2047
rect 47540 2047 47550 2052
rect 47732 2047 47742 2052
rect 47360 1996 47370 2001
rect 47540 2001 47551 2047
rect 47731 2001 47742 2047
rect 47912 2047 47922 2052
rect 47540 1996 47550 2001
rect 47732 1996 47742 2001
rect 47912 2001 47923 2047
rect 47912 1996 47922 2001
rect 47606 1969 47676 1970
rect 47978 1969 48048 2514
rect 48104 2047 48114 2052
rect 48103 2001 48114 2047
rect 48284 2047 48294 2052
rect 48104 1996 48114 2001
rect 48284 2001 48295 2047
rect 48284 1996 48294 2001
rect 48326 1969 48400 1982
rect 39442 1957 39537 1969
rect 39442 1781 39497 1957
rect 39531 1781 39537 1957
rect 39442 1769 39537 1781
rect 39749 1957 39909 1969
rect 39749 1781 39755 1957
rect 39789 1781 39869 1957
rect 39903 1781 39909 1957
rect 39749 1769 39909 1781
rect 40121 1957 40281 1969
rect 40121 1781 40127 1957
rect 40161 1781 40241 1957
rect 40275 1781 40281 1957
rect 40121 1769 40281 1781
rect 40493 1957 40653 1969
rect 40493 1781 40499 1957
rect 40533 1781 40613 1957
rect 40647 1781 40653 1957
rect 40493 1769 40653 1781
rect 40865 1957 41025 1969
rect 40865 1781 40871 1957
rect 40905 1781 40985 1957
rect 41019 1781 41025 1957
rect 40865 1769 41025 1781
rect 41237 1957 41397 1969
rect 41237 1781 41243 1957
rect 41277 1781 41357 1957
rect 41391 1781 41397 1957
rect 41237 1769 41397 1781
rect 41609 1957 41769 1969
rect 41609 1781 41615 1957
rect 41649 1781 41729 1957
rect 41763 1781 41769 1957
rect 41609 1769 41769 1781
rect 41981 1957 42141 1969
rect 41981 1781 41987 1957
rect 42021 1781 42101 1957
rect 42135 1781 42141 1957
rect 41981 1769 42141 1781
rect 42353 1957 42513 1969
rect 42353 1781 42359 1957
rect 42393 1781 42473 1957
rect 42507 1781 42513 1957
rect 42353 1769 42513 1781
rect 42725 1957 42885 1969
rect 42725 1781 42731 1957
rect 42765 1781 42845 1957
rect 42879 1781 42885 1957
rect 42725 1769 42885 1781
rect 43097 1957 43257 1969
rect 43097 1781 43103 1957
rect 43137 1781 43217 1957
rect 43251 1781 43257 1957
rect 43097 1769 43257 1781
rect 43469 1957 43629 1969
rect 43469 1781 43475 1957
rect 43509 1781 43589 1957
rect 43623 1781 43629 1957
rect 43469 1769 43629 1781
rect 43841 1957 44001 1969
rect 43841 1781 43847 1957
rect 43881 1781 43961 1957
rect 43995 1781 44001 1957
rect 43841 1769 44001 1781
rect 44213 1957 44373 1969
rect 44213 1781 44219 1957
rect 44253 1781 44333 1957
rect 44367 1781 44373 1957
rect 44213 1769 44373 1781
rect 44585 1957 44745 1969
rect 44585 1781 44591 1957
rect 44625 1781 44705 1957
rect 44739 1781 44745 1957
rect 44585 1769 44745 1781
rect 44957 1957 45117 1969
rect 44957 1781 44963 1957
rect 44997 1781 45077 1957
rect 45111 1781 45117 1957
rect 44957 1769 45117 1781
rect 45329 1957 45489 1969
rect 45329 1781 45335 1957
rect 45369 1781 45449 1957
rect 45483 1781 45489 1957
rect 45329 1769 45489 1781
rect 45701 1957 45861 1969
rect 45701 1781 45707 1957
rect 45741 1781 45821 1957
rect 45855 1781 45861 1957
rect 45701 1769 45861 1781
rect 46073 1957 46233 1969
rect 46073 1781 46079 1957
rect 46113 1781 46193 1957
rect 46227 1781 46233 1957
rect 46073 1769 46233 1781
rect 46445 1957 46605 1969
rect 46445 1781 46451 1957
rect 46485 1781 46565 1957
rect 46599 1781 46605 1957
rect 46445 1769 46605 1781
rect 46817 1957 46977 1969
rect 46817 1781 46823 1957
rect 46857 1781 46937 1957
rect 46971 1781 46977 1957
rect 46817 1769 46977 1781
rect 47189 1957 47349 1969
rect 47189 1781 47195 1957
rect 47229 1781 47309 1957
rect 47343 1781 47349 1957
rect 47189 1769 47349 1781
rect 47561 1957 47721 1969
rect 47561 1781 47567 1957
rect 47601 1781 47681 1957
rect 47715 1781 47721 1957
rect 47561 1769 47721 1781
rect 47933 1957 48093 1969
rect 47933 1781 47939 1957
rect 47973 1781 48053 1957
rect 48087 1781 48093 1957
rect 47933 1769 48093 1781
rect 48305 1957 48400 1969
rect 48305 1781 48311 1957
rect 48345 1781 48400 1957
rect 48305 1769 48400 1781
rect 39442 1551 39516 1769
rect 39794 1738 39864 1769
rect 39546 1732 40112 1738
rect 39546 1588 39558 1732
rect 39728 1588 39930 1732
rect 40100 1588 40112 1732
rect 39546 1582 40112 1588
rect 39794 1551 39864 1582
rect 40166 1551 40236 1769
rect 40291 1732 40483 1737
rect 40291 1691 40302 1732
rect 40292 1629 40302 1691
rect 40291 1588 40302 1629
rect 40472 1691 40483 1732
rect 40472 1629 40482 1691
rect 40472 1588 40483 1629
rect 40291 1583 40483 1588
rect 40538 1551 40608 1769
rect 40663 1732 40855 1737
rect 40663 1691 40674 1732
rect 40664 1629 40674 1691
rect 40663 1588 40674 1629
rect 40844 1691 40855 1732
rect 40844 1629 40854 1691
rect 40844 1588 40855 1629
rect 40663 1583 40855 1588
rect 40910 1551 40980 1769
rect 41035 1732 41227 1737
rect 41035 1691 41046 1732
rect 41036 1629 41046 1691
rect 41035 1588 41046 1629
rect 41216 1691 41227 1732
rect 41216 1629 41226 1691
rect 41216 1588 41227 1629
rect 41035 1583 41227 1588
rect 41282 1551 41352 1769
rect 41407 1732 41599 1737
rect 41407 1691 41418 1732
rect 41408 1629 41418 1691
rect 41407 1588 41418 1629
rect 41588 1691 41599 1732
rect 41588 1629 41598 1691
rect 41588 1588 41599 1629
rect 41407 1583 41599 1588
rect 41654 1551 41724 1769
rect 42026 1738 42096 1769
rect 41778 1732 42344 1738
rect 41778 1588 41790 1732
rect 41960 1588 42162 1732
rect 42332 1588 42344 1732
rect 41778 1582 42344 1588
rect 42026 1551 42096 1582
rect 42398 1551 42468 1769
rect 42523 1732 42715 1737
rect 42523 1691 42534 1732
rect 42524 1629 42534 1691
rect 42523 1588 42534 1629
rect 42704 1691 42715 1732
rect 42704 1629 42714 1691
rect 42704 1588 42715 1629
rect 42523 1583 42715 1588
rect 42770 1551 42840 1769
rect 42895 1732 43087 1737
rect 42895 1691 42906 1732
rect 42896 1629 42906 1691
rect 42895 1588 42906 1629
rect 43076 1691 43087 1732
rect 43076 1629 43086 1691
rect 43076 1588 43087 1629
rect 42895 1583 43087 1588
rect 43142 1551 43212 1769
rect 43267 1732 43459 1737
rect 43267 1691 43278 1732
rect 43268 1629 43278 1691
rect 43267 1588 43278 1629
rect 43448 1691 43459 1732
rect 43448 1629 43458 1691
rect 43448 1588 43459 1629
rect 43267 1583 43459 1588
rect 43514 1551 43584 1769
rect 43639 1732 43831 1737
rect 43639 1691 43650 1732
rect 43640 1629 43650 1691
rect 43639 1588 43650 1629
rect 43820 1691 43831 1732
rect 43820 1629 43830 1691
rect 43820 1588 43831 1629
rect 43639 1583 43831 1588
rect 43886 1551 43956 1769
rect 44011 1732 44203 1737
rect 44011 1691 44022 1732
rect 44012 1629 44022 1691
rect 44011 1588 44022 1629
rect 44192 1691 44203 1732
rect 44192 1629 44202 1691
rect 44192 1588 44203 1629
rect 44011 1583 44203 1588
rect 44258 1551 44328 1769
rect 44383 1732 44575 1737
rect 44383 1691 44394 1732
rect 44384 1629 44394 1691
rect 44383 1588 44394 1629
rect 44564 1691 44575 1732
rect 44564 1629 44574 1691
rect 44564 1588 44575 1629
rect 44383 1583 44575 1588
rect 44630 1551 44700 1769
rect 44755 1732 44947 1737
rect 44755 1691 44766 1732
rect 44756 1629 44766 1691
rect 44755 1588 44766 1629
rect 44936 1691 44947 1732
rect 44936 1629 44946 1691
rect 44936 1588 44947 1629
rect 44755 1583 44947 1588
rect 45002 1551 45072 1769
rect 45127 1732 45319 1737
rect 45127 1691 45138 1732
rect 45128 1629 45138 1691
rect 45127 1588 45138 1629
rect 45308 1691 45319 1732
rect 45308 1629 45318 1691
rect 45308 1588 45319 1629
rect 45127 1583 45319 1588
rect 45374 1551 45444 1769
rect 45499 1732 45691 1737
rect 45499 1691 45510 1732
rect 45500 1629 45510 1691
rect 45499 1588 45510 1629
rect 45680 1691 45691 1732
rect 45680 1629 45690 1691
rect 45680 1588 45691 1629
rect 45499 1583 45691 1588
rect 45746 1551 45816 1769
rect 45871 1732 46063 1737
rect 45871 1691 45882 1732
rect 45872 1629 45882 1691
rect 45871 1588 45882 1629
rect 46052 1691 46063 1732
rect 46052 1629 46062 1691
rect 46052 1588 46063 1629
rect 45871 1583 46063 1588
rect 46118 1551 46188 1769
rect 46243 1732 46435 1737
rect 46243 1691 46254 1732
rect 46244 1629 46254 1691
rect 46243 1588 46254 1629
rect 46424 1691 46435 1732
rect 46424 1629 46434 1691
rect 46424 1588 46435 1629
rect 46243 1583 46435 1588
rect 46490 1551 46560 1769
rect 46615 1732 46807 1737
rect 46615 1691 46626 1732
rect 46616 1629 46626 1691
rect 46615 1588 46626 1629
rect 46796 1691 46807 1732
rect 46796 1629 46806 1691
rect 46796 1588 46807 1629
rect 46615 1583 46807 1588
rect 46862 1551 46932 1769
rect 46987 1732 47179 1737
rect 46987 1691 46998 1732
rect 46988 1629 46998 1691
rect 46987 1588 46998 1629
rect 47168 1691 47179 1732
rect 47168 1629 47178 1691
rect 47168 1588 47179 1629
rect 46987 1583 47179 1588
rect 47234 1551 47304 1769
rect 47359 1732 47551 1737
rect 47359 1691 47370 1732
rect 47360 1629 47370 1691
rect 47359 1588 47370 1629
rect 47540 1691 47551 1732
rect 47540 1629 47550 1691
rect 47540 1588 47551 1629
rect 47359 1583 47551 1588
rect 47606 1551 47676 1769
rect 47731 1732 47923 1737
rect 47731 1691 47742 1732
rect 47732 1629 47742 1691
rect 47731 1588 47742 1629
rect 47912 1691 47923 1732
rect 47912 1629 47922 1691
rect 47912 1588 47923 1629
rect 47731 1583 47923 1588
rect 47978 1551 48048 1769
rect 48103 1732 48295 1737
rect 48103 1691 48114 1732
rect 48104 1629 48114 1691
rect 48103 1588 48114 1629
rect 48284 1691 48295 1732
rect 48284 1629 48294 1691
rect 48284 1588 48295 1629
rect 48103 1583 48295 1588
rect 48326 1551 48400 1769
rect 39442 1539 39537 1551
rect 39442 1363 39497 1539
rect 39531 1363 39537 1539
rect 39442 1351 39537 1363
rect 39749 1539 39909 1551
rect 39749 1363 39755 1539
rect 39789 1363 39869 1539
rect 39903 1363 39909 1539
rect 39749 1351 39909 1363
rect 40121 1539 40281 1551
rect 40121 1363 40127 1539
rect 40161 1363 40241 1539
rect 40275 1363 40281 1539
rect 40121 1351 40281 1363
rect 40493 1539 40653 1551
rect 40493 1363 40499 1539
rect 40533 1363 40613 1539
rect 40647 1363 40653 1539
rect 40493 1351 40653 1363
rect 40865 1539 41025 1551
rect 40865 1363 40871 1539
rect 40905 1363 40985 1539
rect 41019 1363 41025 1539
rect 40865 1351 41025 1363
rect 41237 1539 41397 1551
rect 41237 1363 41243 1539
rect 41277 1363 41357 1539
rect 41391 1363 41397 1539
rect 41237 1351 41397 1363
rect 41609 1539 41769 1551
rect 41609 1363 41615 1539
rect 41649 1363 41729 1539
rect 41763 1363 41769 1539
rect 41609 1351 41769 1363
rect 41981 1539 42141 1551
rect 41981 1363 41987 1539
rect 42021 1363 42101 1539
rect 42135 1363 42141 1539
rect 41981 1351 42141 1363
rect 42353 1539 42513 1551
rect 42353 1363 42359 1539
rect 42393 1363 42473 1539
rect 42507 1363 42513 1539
rect 42353 1351 42513 1363
rect 42725 1539 42885 1551
rect 42725 1363 42731 1539
rect 42765 1363 42845 1539
rect 42879 1363 42885 1539
rect 42725 1351 42885 1363
rect 43097 1539 43257 1551
rect 43097 1363 43103 1539
rect 43137 1363 43217 1539
rect 43251 1363 43257 1539
rect 43097 1351 43257 1363
rect 43469 1539 43629 1551
rect 43469 1363 43475 1539
rect 43509 1363 43589 1539
rect 43623 1363 43629 1539
rect 43469 1351 43629 1363
rect 43841 1539 44001 1551
rect 43841 1363 43847 1539
rect 43881 1363 43961 1539
rect 43995 1363 44001 1539
rect 43841 1351 44001 1363
rect 44213 1539 44373 1551
rect 44213 1363 44219 1539
rect 44253 1363 44333 1539
rect 44367 1363 44373 1539
rect 44213 1351 44373 1363
rect 44585 1539 44745 1551
rect 44585 1363 44591 1539
rect 44625 1363 44705 1539
rect 44739 1363 44745 1539
rect 44585 1351 44745 1363
rect 44957 1539 45117 1551
rect 44957 1363 44963 1539
rect 44997 1363 45077 1539
rect 45111 1363 45117 1539
rect 44957 1351 45117 1363
rect 45329 1539 45489 1551
rect 45329 1363 45335 1539
rect 45369 1363 45449 1539
rect 45483 1363 45489 1539
rect 45329 1351 45489 1363
rect 45701 1539 45861 1551
rect 45701 1363 45707 1539
rect 45741 1363 45821 1539
rect 45855 1363 45861 1539
rect 45701 1351 45861 1363
rect 46073 1539 46233 1551
rect 46073 1363 46079 1539
rect 46113 1363 46193 1539
rect 46227 1363 46233 1539
rect 46073 1351 46233 1363
rect 46445 1539 46605 1551
rect 46445 1363 46451 1539
rect 46485 1363 46565 1539
rect 46599 1363 46605 1539
rect 46445 1351 46605 1363
rect 46817 1539 46977 1551
rect 46817 1363 46823 1539
rect 46857 1363 46937 1539
rect 46971 1363 46977 1539
rect 46817 1351 46977 1363
rect 47189 1539 47349 1551
rect 47189 1363 47195 1539
rect 47229 1363 47309 1539
rect 47343 1363 47349 1539
rect 47189 1351 47349 1363
rect 47561 1539 47721 1551
rect 47561 1363 47567 1539
rect 47601 1363 47681 1539
rect 47715 1363 47721 1539
rect 47561 1351 47721 1363
rect 47933 1539 48093 1551
rect 47933 1363 47939 1539
rect 47973 1363 48053 1539
rect 48087 1363 48093 1539
rect 47933 1351 48093 1363
rect 48305 1539 48400 1551
rect 48305 1363 48311 1539
rect 48345 1363 48400 1539
rect 48305 1351 48400 1363
rect 39442 1133 39516 1351
rect 39794 1320 39864 1351
rect 39546 1314 40112 1320
rect 39546 1170 39558 1314
rect 39728 1170 39930 1314
rect 40100 1170 40112 1314
rect 39546 1164 40112 1170
rect 39794 1133 39864 1164
rect 40166 1133 40236 1351
rect 40291 1314 40483 1319
rect 40291 1273 40302 1314
rect 40292 1211 40302 1273
rect 40291 1170 40302 1211
rect 40472 1273 40483 1314
rect 40472 1211 40482 1273
rect 40472 1170 40483 1211
rect 40291 1165 40483 1170
rect 40538 1133 40608 1351
rect 40663 1314 40855 1319
rect 40663 1273 40674 1314
rect 40664 1211 40674 1273
rect 40663 1170 40674 1211
rect 40844 1273 40855 1314
rect 40844 1211 40854 1273
rect 40844 1170 40855 1211
rect 40663 1165 40855 1170
rect 40910 1133 40980 1351
rect 41035 1314 41227 1319
rect 41035 1273 41046 1314
rect 41036 1211 41046 1273
rect 41035 1170 41046 1211
rect 41216 1273 41227 1314
rect 41216 1211 41226 1273
rect 41216 1170 41227 1211
rect 41035 1165 41227 1170
rect 41282 1133 41352 1351
rect 41407 1314 41599 1319
rect 41407 1273 41418 1314
rect 41408 1211 41418 1273
rect 41407 1170 41418 1211
rect 41588 1273 41599 1314
rect 41588 1211 41598 1273
rect 41588 1170 41599 1211
rect 41407 1165 41599 1170
rect 41654 1133 41724 1351
rect 42026 1320 42096 1351
rect 41778 1314 42344 1320
rect 41778 1170 41790 1314
rect 41960 1170 42162 1314
rect 42332 1170 42344 1314
rect 41778 1164 42344 1170
rect 42026 1133 42096 1164
rect 42398 1133 42468 1351
rect 42523 1314 42715 1319
rect 42523 1273 42534 1314
rect 42524 1211 42534 1273
rect 42523 1170 42534 1211
rect 42704 1273 42715 1314
rect 42704 1211 42714 1273
rect 42704 1170 42715 1211
rect 42523 1165 42715 1170
rect 42770 1133 42840 1351
rect 42895 1314 43087 1319
rect 42895 1273 42906 1314
rect 42896 1211 42906 1273
rect 42895 1170 42906 1211
rect 43076 1273 43087 1314
rect 43076 1211 43086 1273
rect 43076 1170 43087 1211
rect 42895 1165 43087 1170
rect 43142 1133 43212 1351
rect 43267 1314 43459 1319
rect 43267 1273 43278 1314
rect 43268 1211 43278 1273
rect 43267 1170 43278 1211
rect 43448 1273 43459 1314
rect 43448 1211 43458 1273
rect 43448 1170 43459 1211
rect 43267 1165 43459 1170
rect 43514 1133 43584 1351
rect 43639 1314 43831 1319
rect 43639 1273 43650 1314
rect 43640 1211 43650 1273
rect 43639 1170 43650 1211
rect 43820 1273 43831 1314
rect 43820 1211 43830 1273
rect 43820 1170 43831 1211
rect 43639 1165 43831 1170
rect 43886 1133 43956 1351
rect 44011 1314 44203 1319
rect 44011 1273 44022 1314
rect 44012 1211 44022 1273
rect 44011 1170 44022 1211
rect 44192 1273 44203 1314
rect 44192 1211 44202 1273
rect 44192 1170 44203 1211
rect 44011 1165 44203 1170
rect 44258 1133 44328 1351
rect 44383 1314 44575 1319
rect 44383 1273 44394 1314
rect 44384 1211 44394 1273
rect 44383 1170 44394 1211
rect 44564 1273 44575 1314
rect 44564 1211 44574 1273
rect 44564 1170 44575 1211
rect 44383 1165 44575 1170
rect 44630 1133 44700 1351
rect 44755 1314 44947 1319
rect 44755 1273 44766 1314
rect 44756 1211 44766 1273
rect 44755 1170 44766 1211
rect 44936 1273 44947 1314
rect 44936 1211 44946 1273
rect 44936 1170 44947 1211
rect 44755 1165 44947 1170
rect 45002 1133 45072 1351
rect 45127 1314 45319 1319
rect 45127 1273 45138 1314
rect 45128 1211 45138 1273
rect 45127 1170 45138 1211
rect 45308 1273 45319 1314
rect 45308 1211 45318 1273
rect 45308 1170 45319 1211
rect 45127 1165 45319 1170
rect 45374 1133 45444 1351
rect 45499 1314 45691 1319
rect 45499 1273 45510 1314
rect 45500 1211 45510 1273
rect 45499 1170 45510 1211
rect 45680 1273 45691 1314
rect 45680 1211 45690 1273
rect 45680 1170 45691 1211
rect 45499 1165 45691 1170
rect 45746 1133 45816 1351
rect 45871 1314 46063 1319
rect 45871 1273 45882 1314
rect 45872 1211 45882 1273
rect 45871 1170 45882 1211
rect 46052 1273 46063 1314
rect 46052 1211 46062 1273
rect 46052 1170 46063 1211
rect 45871 1165 46063 1170
rect 46118 1133 46188 1351
rect 46243 1314 46435 1319
rect 46243 1273 46254 1314
rect 46244 1211 46254 1273
rect 46243 1170 46254 1211
rect 46424 1273 46435 1314
rect 46424 1211 46434 1273
rect 46424 1170 46435 1211
rect 46243 1165 46435 1170
rect 46490 1133 46560 1351
rect 46615 1314 46807 1319
rect 46615 1273 46626 1314
rect 46616 1211 46626 1273
rect 46615 1170 46626 1211
rect 46796 1273 46807 1314
rect 46796 1211 46806 1273
rect 46796 1170 46807 1211
rect 46615 1165 46807 1170
rect 46862 1133 46932 1351
rect 46987 1314 47179 1319
rect 46987 1273 46998 1314
rect 46988 1211 46998 1273
rect 46987 1170 46998 1211
rect 47168 1273 47179 1314
rect 47168 1211 47178 1273
rect 47168 1170 47179 1211
rect 46987 1165 47179 1170
rect 47234 1133 47304 1351
rect 47359 1314 47551 1319
rect 47359 1273 47370 1314
rect 47360 1211 47370 1273
rect 47359 1170 47370 1211
rect 47540 1273 47551 1314
rect 47540 1211 47550 1273
rect 47540 1170 47551 1211
rect 47359 1165 47551 1170
rect 47606 1133 47676 1351
rect 47731 1314 47923 1319
rect 47731 1273 47742 1314
rect 47732 1211 47742 1273
rect 47731 1170 47742 1211
rect 47912 1273 47923 1314
rect 47912 1211 47922 1273
rect 47912 1170 47923 1211
rect 47731 1165 47923 1170
rect 47978 1133 48048 1351
rect 48103 1314 48295 1319
rect 48103 1273 48114 1314
rect 48104 1211 48114 1273
rect 48103 1170 48114 1211
rect 48284 1273 48295 1314
rect 48284 1211 48294 1273
rect 48284 1170 48295 1211
rect 48103 1165 48295 1170
rect 48326 1133 48400 1351
rect 39442 1121 39537 1133
rect 39442 945 39497 1121
rect 39531 945 39537 1121
rect 39442 933 39537 945
rect 39749 1121 39909 1133
rect 39749 945 39755 1121
rect 39789 945 39869 1121
rect 39903 945 39909 1121
rect 39749 933 39909 945
rect 40121 1121 40281 1133
rect 40121 945 40127 1121
rect 40161 945 40241 1121
rect 40275 945 40281 1121
rect 40121 933 40281 945
rect 40493 1121 40653 1133
rect 40493 945 40499 1121
rect 40533 945 40613 1121
rect 40647 945 40653 1121
rect 40493 933 40653 945
rect 40865 1121 41025 1133
rect 40865 945 40871 1121
rect 40905 945 40985 1121
rect 41019 945 41025 1121
rect 40865 933 41025 945
rect 41237 1121 41397 1133
rect 41237 945 41243 1121
rect 41277 945 41357 1121
rect 41391 945 41397 1121
rect 41237 933 41397 945
rect 41609 1121 41769 1133
rect 41609 945 41615 1121
rect 41649 945 41729 1121
rect 41763 945 41769 1121
rect 41609 933 41769 945
rect 41981 1121 42141 1133
rect 41981 945 41987 1121
rect 42021 945 42101 1121
rect 42135 945 42141 1121
rect 41981 933 42141 945
rect 42353 1121 42513 1133
rect 42353 945 42359 1121
rect 42393 945 42473 1121
rect 42507 945 42513 1121
rect 42353 933 42513 945
rect 42725 1121 42885 1133
rect 42725 945 42731 1121
rect 42765 945 42845 1121
rect 42879 945 42885 1121
rect 42725 933 42885 945
rect 43097 1121 43257 1133
rect 43097 945 43103 1121
rect 43137 945 43217 1121
rect 43251 945 43257 1121
rect 43097 933 43257 945
rect 43469 1121 43629 1133
rect 43469 945 43475 1121
rect 43509 945 43589 1121
rect 43623 945 43629 1121
rect 43469 933 43629 945
rect 43841 1121 44001 1133
rect 43841 945 43847 1121
rect 43881 945 43961 1121
rect 43995 945 44001 1121
rect 43841 933 44001 945
rect 44213 1121 44373 1133
rect 44213 945 44219 1121
rect 44253 945 44333 1121
rect 44367 945 44373 1121
rect 44213 933 44373 945
rect 44585 1121 44745 1133
rect 44585 945 44591 1121
rect 44625 945 44705 1121
rect 44739 945 44745 1121
rect 44585 933 44745 945
rect 44957 1121 45117 1133
rect 44957 945 44963 1121
rect 44997 945 45077 1121
rect 45111 945 45117 1121
rect 44957 933 45117 945
rect 45329 1121 45489 1133
rect 45329 945 45335 1121
rect 45369 945 45449 1121
rect 45483 945 45489 1121
rect 45329 933 45489 945
rect 45701 1121 45861 1133
rect 45701 945 45707 1121
rect 45741 945 45821 1121
rect 45855 945 45861 1121
rect 45701 933 45861 945
rect 46073 1121 46233 1133
rect 46073 945 46079 1121
rect 46113 945 46193 1121
rect 46227 945 46233 1121
rect 46073 933 46233 945
rect 46445 1121 46605 1133
rect 46445 945 46451 1121
rect 46485 945 46565 1121
rect 46599 945 46605 1121
rect 46445 933 46605 945
rect 46817 1121 46977 1133
rect 46817 945 46823 1121
rect 46857 945 46937 1121
rect 46971 945 46977 1121
rect 46817 933 46977 945
rect 47189 1121 47349 1133
rect 47189 945 47195 1121
rect 47229 945 47309 1121
rect 47343 945 47349 1121
rect 47189 933 47349 945
rect 47561 1121 47721 1133
rect 47561 945 47567 1121
rect 47601 945 47681 1121
rect 47715 945 47721 1121
rect 47561 933 47721 945
rect 47933 1121 48093 1133
rect 47933 945 47939 1121
rect 47973 945 48053 1121
rect 48087 945 48093 1121
rect 47933 933 48093 945
rect 48305 1121 48400 1133
rect 48305 945 48311 1121
rect 48345 945 48400 1121
rect 48305 933 48400 945
rect 39442 715 39516 933
rect 39794 902 39864 933
rect 39546 896 40112 902
rect 39546 752 39558 896
rect 39728 752 39930 896
rect 40100 752 40112 896
rect 39546 746 40112 752
rect 39794 715 39864 746
rect 40166 715 40236 933
rect 40291 896 40483 901
rect 40291 855 40302 896
rect 40292 793 40302 855
rect 40291 752 40302 793
rect 40472 855 40483 896
rect 40472 793 40482 855
rect 40472 752 40483 793
rect 40291 747 40483 752
rect 40538 715 40608 933
rect 40663 896 40855 901
rect 40663 855 40674 896
rect 40664 793 40674 855
rect 40663 752 40674 793
rect 40844 855 40855 896
rect 40844 793 40854 855
rect 40844 752 40855 793
rect 40663 747 40855 752
rect 40910 715 40980 933
rect 41035 896 41227 901
rect 41035 855 41046 896
rect 41036 793 41046 855
rect 41035 752 41046 793
rect 41216 855 41227 896
rect 41216 793 41226 855
rect 41216 752 41227 793
rect 41035 747 41227 752
rect 41282 715 41352 933
rect 41407 896 41599 901
rect 41407 855 41418 896
rect 41408 793 41418 855
rect 41407 752 41418 793
rect 41588 855 41599 896
rect 41588 793 41598 855
rect 41588 752 41599 793
rect 41407 747 41599 752
rect 41654 715 41724 933
rect 42026 902 42096 933
rect 41778 896 42344 902
rect 41778 752 41790 896
rect 41960 752 42162 896
rect 42332 752 42344 896
rect 41778 746 42344 752
rect 42026 715 42096 746
rect 42398 715 42468 933
rect 42523 896 42715 901
rect 42523 855 42534 896
rect 42524 793 42534 855
rect 42523 752 42534 793
rect 42704 855 42715 896
rect 42704 793 42714 855
rect 42704 752 42715 793
rect 42523 747 42715 752
rect 42770 715 42840 933
rect 42895 896 43087 901
rect 42895 855 42906 896
rect 42896 793 42906 855
rect 42895 752 42906 793
rect 43076 855 43087 896
rect 43076 793 43086 855
rect 43076 752 43087 793
rect 42895 747 43087 752
rect 43142 715 43212 933
rect 43267 896 43459 901
rect 43267 855 43278 896
rect 43268 793 43278 855
rect 43267 752 43278 793
rect 43448 855 43459 896
rect 43448 793 43458 855
rect 43448 752 43459 793
rect 43267 747 43459 752
rect 43514 715 43584 933
rect 43639 896 43831 901
rect 43639 855 43650 896
rect 43640 793 43650 855
rect 43639 752 43650 793
rect 43820 855 43831 896
rect 43820 793 43830 855
rect 43820 752 43831 793
rect 43639 747 43831 752
rect 43886 715 43956 933
rect 44011 896 44203 901
rect 44011 855 44022 896
rect 44012 793 44022 855
rect 44011 752 44022 793
rect 44192 855 44203 896
rect 44192 793 44202 855
rect 44192 752 44203 793
rect 44011 747 44203 752
rect 44258 715 44328 933
rect 44383 896 44575 901
rect 44383 855 44394 896
rect 44384 793 44394 855
rect 44383 752 44394 793
rect 44564 855 44575 896
rect 44564 793 44574 855
rect 44564 752 44575 793
rect 44383 747 44575 752
rect 44630 715 44700 933
rect 44755 896 44947 901
rect 44755 855 44766 896
rect 44756 793 44766 855
rect 44755 752 44766 793
rect 44936 855 44947 896
rect 44936 793 44946 855
rect 44936 752 44947 793
rect 44755 747 44947 752
rect 45002 715 45072 933
rect 45127 896 45319 901
rect 45127 855 45138 896
rect 45128 793 45138 855
rect 45127 752 45138 793
rect 45308 855 45319 896
rect 45308 793 45318 855
rect 45308 752 45319 793
rect 45127 747 45319 752
rect 45374 715 45444 933
rect 45499 896 45691 901
rect 45499 855 45510 896
rect 45500 793 45510 855
rect 45499 752 45510 793
rect 45680 855 45691 896
rect 45680 793 45690 855
rect 45680 752 45691 793
rect 45499 747 45691 752
rect 45746 715 45816 933
rect 45871 896 46063 901
rect 45871 855 45882 896
rect 45872 793 45882 855
rect 45871 752 45882 793
rect 46052 855 46063 896
rect 46052 793 46062 855
rect 46052 752 46063 793
rect 45871 747 46063 752
rect 46118 715 46188 933
rect 46243 896 46435 901
rect 46243 855 46254 896
rect 46244 793 46254 855
rect 46243 752 46254 793
rect 46424 855 46435 896
rect 46424 793 46434 855
rect 46424 752 46435 793
rect 46243 747 46435 752
rect 46490 715 46560 933
rect 46615 896 46807 901
rect 46615 855 46626 896
rect 46616 793 46626 855
rect 46615 752 46626 793
rect 46796 855 46807 896
rect 46796 793 46806 855
rect 46796 752 46807 793
rect 46615 747 46807 752
rect 46862 715 46932 933
rect 46987 896 47179 901
rect 46987 855 46998 896
rect 46988 793 46998 855
rect 46987 752 46998 793
rect 47168 855 47179 896
rect 47168 793 47178 855
rect 47168 752 47179 793
rect 46987 747 47179 752
rect 47234 715 47304 933
rect 47359 896 47551 901
rect 47359 855 47370 896
rect 47360 793 47370 855
rect 47359 752 47370 793
rect 47540 855 47551 896
rect 47540 793 47550 855
rect 47540 752 47551 793
rect 47359 747 47551 752
rect 47606 715 47676 933
rect 47731 896 47923 901
rect 47731 855 47742 896
rect 47732 793 47742 855
rect 47731 752 47742 793
rect 47912 855 47923 896
rect 47912 793 47922 855
rect 47912 752 47923 793
rect 47731 747 47923 752
rect 47978 715 48048 933
rect 48103 896 48295 901
rect 48103 855 48114 896
rect 48104 793 48114 855
rect 48103 752 48114 793
rect 48284 855 48295 896
rect 48284 793 48294 855
rect 48284 752 48295 793
rect 48103 747 48295 752
rect 48326 715 48400 933
rect 39442 703 39537 715
rect 39442 527 39497 703
rect 39531 527 39537 703
rect 39442 515 39537 527
rect 39749 703 39909 715
rect 39749 527 39755 703
rect 39789 527 39869 703
rect 39903 527 39909 703
rect 39749 515 39909 527
rect 40121 703 40281 715
rect 40121 527 40127 703
rect 40161 527 40241 703
rect 40275 527 40281 703
rect 40121 515 40281 527
rect 40493 703 40653 715
rect 40493 527 40499 703
rect 40533 527 40613 703
rect 40647 527 40653 703
rect 40493 515 40653 527
rect 40865 703 41025 715
rect 40865 527 40871 703
rect 40905 527 40985 703
rect 41019 527 41025 703
rect 40865 515 41025 527
rect 41237 703 41397 715
rect 41237 527 41243 703
rect 41277 527 41357 703
rect 41391 527 41397 703
rect 41237 515 41397 527
rect 41609 703 41769 715
rect 41609 527 41615 703
rect 41649 527 41729 703
rect 41763 527 41769 703
rect 41609 515 41769 527
rect 41981 703 42141 715
rect 41981 527 41987 703
rect 42021 527 42101 703
rect 42135 527 42141 703
rect 41981 515 42141 527
rect 42353 703 42513 715
rect 42353 527 42359 703
rect 42393 527 42473 703
rect 42507 527 42513 703
rect 42353 515 42513 527
rect 42725 703 42885 715
rect 42725 527 42731 703
rect 42765 527 42845 703
rect 42879 527 42885 703
rect 42725 515 42885 527
rect 43097 703 43257 715
rect 43097 527 43103 703
rect 43137 527 43217 703
rect 43251 527 43257 703
rect 43097 515 43257 527
rect 43469 703 43629 715
rect 43469 527 43475 703
rect 43509 527 43589 703
rect 43623 527 43629 703
rect 43469 515 43629 527
rect 43841 703 44001 715
rect 43841 527 43847 703
rect 43881 527 43961 703
rect 43995 527 44001 703
rect 43841 515 44001 527
rect 44213 703 44373 715
rect 44213 527 44219 703
rect 44253 527 44333 703
rect 44367 527 44373 703
rect 44213 515 44373 527
rect 44585 703 44745 715
rect 44585 527 44591 703
rect 44625 527 44705 703
rect 44739 527 44745 703
rect 44585 515 44745 527
rect 44957 703 45117 715
rect 44957 527 44963 703
rect 44997 527 45077 703
rect 45111 527 45117 703
rect 44957 515 45117 527
rect 45329 703 45489 715
rect 45329 527 45335 703
rect 45369 527 45449 703
rect 45483 527 45489 703
rect 45329 515 45489 527
rect 45701 703 45861 715
rect 45701 527 45707 703
rect 45741 527 45821 703
rect 45855 527 45861 703
rect 45701 515 45861 527
rect 46073 703 46233 715
rect 46073 527 46079 703
rect 46113 527 46193 703
rect 46227 527 46233 703
rect 46073 515 46233 527
rect 46445 703 46605 715
rect 46445 527 46451 703
rect 46485 527 46565 703
rect 46599 527 46605 703
rect 46445 515 46605 527
rect 46817 703 46977 715
rect 46817 527 46823 703
rect 46857 527 46937 703
rect 46971 527 46977 703
rect 46817 515 46977 527
rect 47189 703 47349 715
rect 47189 527 47195 703
rect 47229 527 47309 703
rect 47343 527 47349 703
rect 47189 515 47349 527
rect 47561 703 47721 715
rect 47561 527 47567 703
rect 47601 527 47681 703
rect 47715 527 47721 703
rect 47561 515 47721 527
rect 47933 703 48093 715
rect 47933 527 47939 703
rect 47973 527 48053 703
rect 48087 527 48093 703
rect 47933 515 48093 527
rect 48305 703 48400 715
rect 48305 527 48311 703
rect 48345 527 48400 703
rect 48305 515 48400 527
rect 39442 392 39516 515
rect 39548 483 39558 488
rect 39547 478 39558 483
rect 39546 432 39558 478
rect 39728 483 39738 488
rect 39728 478 39739 483
rect 39794 478 39864 515
rect 40166 514 40236 515
rect 40538 514 40608 515
rect 40910 514 40980 515
rect 41282 514 41352 515
rect 41654 514 41724 515
rect 39920 483 39930 488
rect 39919 478 39930 483
rect 39728 432 39930 478
rect 40100 483 40110 488
rect 40100 478 40111 483
rect 40100 432 40112 478
rect 39546 420 40112 432
rect 40172 400 40230 514
rect 40292 483 40302 488
rect 40291 437 40302 483
rect 40472 483 40482 488
rect 40664 483 40674 488
rect 40292 432 40302 437
rect 40472 437 40483 483
rect 40663 437 40674 483
rect 40844 483 40854 488
rect 40472 432 40482 437
rect 40664 432 40674 437
rect 40844 437 40855 483
rect 40844 432 40854 437
rect 40916 400 40974 514
rect 41036 483 41046 488
rect 41035 437 41046 483
rect 41216 483 41226 488
rect 41408 483 41418 488
rect 41036 432 41046 437
rect 41216 437 41227 483
rect 41407 437 41418 483
rect 41588 483 41598 488
rect 41216 432 41226 437
rect 41408 432 41418 437
rect 41588 437 41599 483
rect 41588 432 41598 437
rect 41660 400 41718 514
rect 41780 483 41790 488
rect 41779 478 41790 483
rect 41778 432 41790 478
rect 41960 483 41970 488
rect 41960 478 41971 483
rect 42026 478 42096 515
rect 42398 514 42468 515
rect 42770 514 42840 515
rect 43142 514 43212 515
rect 43514 514 43584 515
rect 43886 514 43956 515
rect 44258 514 44328 515
rect 44630 514 44700 515
rect 45002 514 45072 515
rect 45374 514 45444 515
rect 45746 514 45816 515
rect 46118 514 46188 515
rect 46490 514 46560 515
rect 46862 514 46932 515
rect 47234 514 47304 515
rect 47606 514 47676 515
rect 47978 514 48048 515
rect 42152 483 42162 488
rect 42151 478 42162 483
rect 41960 432 42162 478
rect 42332 483 42342 488
rect 42332 478 42343 483
rect 42332 432 42344 478
rect 41778 420 42344 432
rect 42404 400 42462 514
rect 42524 483 42534 488
rect 42523 437 42534 483
rect 42704 483 42714 488
rect 42896 483 42906 488
rect 42524 432 42534 437
rect 42704 437 42715 483
rect 42895 437 42906 483
rect 43076 483 43086 488
rect 42704 432 42714 437
rect 42896 432 42906 437
rect 43076 437 43087 483
rect 43076 432 43086 437
rect 43148 400 43206 514
rect 43268 483 43278 488
rect 43267 437 43278 483
rect 43448 483 43458 488
rect 43640 483 43650 488
rect 43268 432 43278 437
rect 43448 437 43459 483
rect 43639 437 43650 483
rect 43820 483 43830 488
rect 43448 432 43458 437
rect 43640 432 43650 437
rect 43820 437 43831 483
rect 43820 432 43830 437
rect 43892 400 43950 514
rect 44012 483 44022 488
rect 44011 437 44022 483
rect 44192 483 44202 488
rect 44384 483 44394 488
rect 44012 432 44022 437
rect 44192 437 44203 483
rect 44383 437 44394 483
rect 44564 483 44574 488
rect 44192 432 44202 437
rect 44384 432 44394 437
rect 44564 437 44575 483
rect 44564 432 44574 437
rect 44636 400 44694 514
rect 44756 483 44766 488
rect 44755 437 44766 483
rect 44936 483 44946 488
rect 45128 483 45138 488
rect 44756 432 44766 437
rect 44936 437 44947 483
rect 45127 437 45138 483
rect 45308 483 45318 488
rect 44936 432 44946 437
rect 45128 432 45138 437
rect 45308 437 45319 483
rect 45308 432 45318 437
rect 45380 400 45438 514
rect 45500 483 45510 488
rect 45499 437 45510 483
rect 45680 483 45690 488
rect 45872 483 45882 488
rect 45500 432 45510 437
rect 45680 437 45691 483
rect 45871 437 45882 483
rect 46052 483 46062 488
rect 45680 432 45690 437
rect 45872 432 45882 437
rect 46052 437 46063 483
rect 46052 432 46062 437
rect 46124 400 46182 514
rect 46244 483 46254 488
rect 46243 437 46254 483
rect 46424 483 46434 488
rect 46616 483 46626 488
rect 46244 432 46254 437
rect 46424 437 46435 483
rect 46615 437 46626 483
rect 46796 483 46806 488
rect 46424 432 46434 437
rect 46616 432 46626 437
rect 46796 437 46807 483
rect 46796 432 46806 437
rect 46868 400 46926 514
rect 46988 483 46998 488
rect 46987 437 46998 483
rect 47168 483 47178 488
rect 47360 483 47370 488
rect 46988 432 46998 437
rect 47168 437 47179 483
rect 47359 437 47370 483
rect 47540 483 47550 488
rect 47168 432 47178 437
rect 47360 432 47370 437
rect 47540 437 47551 483
rect 47540 432 47550 437
rect 47612 400 47670 514
rect 47732 483 47742 488
rect 47731 437 47742 483
rect 47912 483 47922 488
rect 48104 483 48114 488
rect 47732 432 47742 437
rect 47912 437 47923 483
rect 48103 437 48114 483
rect 48284 483 48294 488
rect 47912 432 47922 437
rect 48104 432 48114 437
rect 48284 437 48295 483
rect 48284 432 48294 437
rect 40154 394 40248 400
rect 39442 386 39580 392
rect 39442 316 39498 386
rect 39568 316 39580 386
rect 40154 324 40166 394
rect 40236 324 40248 394
rect 40154 318 40248 324
rect 40898 394 40992 400
rect 40898 324 40910 394
rect 40980 324 40992 394
rect 40898 318 40992 324
rect 41642 394 41736 400
rect 41642 324 41654 394
rect 41724 324 41736 394
rect 41642 318 41736 324
rect 42386 394 42480 400
rect 42386 324 42398 394
rect 42468 324 42480 394
rect 42386 318 42480 324
rect 43130 394 43224 400
rect 43130 324 43142 394
rect 43212 324 43224 394
rect 43130 318 43224 324
rect 43874 394 43968 400
rect 43874 324 43886 394
rect 43956 324 43968 394
rect 43874 318 43968 324
rect 44618 394 44712 400
rect 44618 324 44630 394
rect 44700 324 44712 394
rect 44618 318 44712 324
rect 45362 394 45456 400
rect 45362 324 45374 394
rect 45444 324 45456 394
rect 45362 318 45456 324
rect 46106 394 46200 400
rect 46106 324 46118 394
rect 46188 324 46200 394
rect 46106 318 46200 324
rect 46850 394 46944 400
rect 46850 324 46862 394
rect 46932 324 46944 394
rect 46850 318 46944 324
rect 47594 394 47688 400
rect 48326 396 48400 515
rect 47594 324 47606 394
rect 47676 324 47688 394
rect 47594 318 47688 324
rect 48256 390 48400 396
rect 48256 320 48268 390
rect 48338 320 48400 390
rect 39442 310 39580 316
rect 39442 278 39516 310
rect 40172 278 40230 318
rect 40916 278 40974 318
rect 41660 278 41718 318
rect 42404 278 42462 318
rect 43148 278 43206 318
rect 43892 278 43950 318
rect 44636 278 44694 318
rect 45380 278 45438 318
rect 46124 278 46182 318
rect 46868 278 46926 318
rect 47612 278 47670 318
rect 48256 314 48400 320
rect 48326 290 48400 314
rect 48326 278 48414 290
rect 39368 78 39378 278
rect 39578 78 39588 278
rect 40092 78 40102 278
rect 40302 78 40312 278
rect 40836 78 40846 278
rect 41046 78 41056 278
rect 41580 78 41590 278
rect 41790 78 41800 278
rect 42324 78 42334 278
rect 42534 78 42544 278
rect 43068 78 43078 278
rect 43278 78 43288 278
rect 43812 78 43822 278
rect 44022 78 44032 278
rect 44556 78 44566 278
rect 44766 78 44776 278
rect 45300 78 45310 278
rect 45510 78 45520 278
rect 46044 78 46054 278
rect 46254 78 46264 278
rect 46788 78 46798 278
rect 46998 78 47008 278
rect 47532 78 47542 278
rect 47742 78 47752 278
rect 48276 78 48286 278
rect 48486 78 48496 278
<< via1 >>
rect 35528 10928 36446 11896
rect 38240 9324 38440 9524
rect 38984 9324 39184 9524
rect 39728 9324 39928 9524
rect 40472 9324 40672 9524
rect 41216 9324 41416 9524
rect 41960 9324 42160 9524
rect 42704 9324 42904 9524
rect 43448 9324 43648 9524
rect 43820 9324 44020 9524
rect 44564 9324 44764 9524
rect 45308 9324 45508 9524
rect 46052 9324 46252 9524
rect 46796 9324 46996 9524
rect 47540 9324 47740 9524
rect 48284 9324 48484 9524
rect 49028 9324 49228 9524
rect 49772 9324 49972 9524
rect 38070 9123 38240 9136
rect 38070 9089 38071 9123
rect 38071 9089 38239 9123
rect 38239 9089 38240 9123
rect 38070 9076 38240 9089
rect 38442 9123 38612 9136
rect 38442 9089 38443 9123
rect 38443 9089 38611 9123
rect 38611 9089 38612 9123
rect 38442 9076 38612 9089
rect 38814 9123 38984 9136
rect 38814 9089 38815 9123
rect 38815 9089 38983 9123
rect 38983 9089 38984 9123
rect 38814 9076 38984 9089
rect 39186 9123 39356 9136
rect 39186 9089 39187 9123
rect 39187 9089 39355 9123
rect 39355 9089 39356 9123
rect 39186 9076 39356 9089
rect 39558 9123 39728 9136
rect 39558 9089 39559 9123
rect 39559 9089 39727 9123
rect 39727 9089 39728 9123
rect 39558 9076 39728 9089
rect 39930 9123 40100 9136
rect 39930 9089 39931 9123
rect 39931 9089 40099 9123
rect 40099 9089 40100 9123
rect 39930 9076 40100 9089
rect 40302 9123 40472 9136
rect 40302 9089 40303 9123
rect 40303 9089 40471 9123
rect 40471 9089 40472 9123
rect 40302 9076 40472 9089
rect 40674 9123 40844 9136
rect 40674 9089 40675 9123
rect 40675 9089 40843 9123
rect 40843 9089 40844 9123
rect 40674 9076 40844 9089
rect 41046 9123 41216 9136
rect 41046 9089 41047 9123
rect 41047 9089 41215 9123
rect 41215 9089 41216 9123
rect 41046 9076 41216 9089
rect 41418 9123 41588 9136
rect 41418 9089 41419 9123
rect 41419 9089 41587 9123
rect 41587 9089 41588 9123
rect 41418 9076 41588 9089
rect 41790 9123 41960 9136
rect 41790 9089 41791 9123
rect 41791 9089 41959 9123
rect 41959 9089 41960 9123
rect 41790 9076 41960 9089
rect 42162 9123 42332 9136
rect 42162 9089 42163 9123
rect 42163 9089 42331 9123
rect 42331 9089 42332 9123
rect 42162 9076 42332 9089
rect 42534 9123 42704 9136
rect 42534 9089 42535 9123
rect 42535 9089 42703 9123
rect 42703 9089 42704 9123
rect 42534 9076 42704 9089
rect 42906 9123 43076 9136
rect 42906 9089 42907 9123
rect 42907 9089 43075 9123
rect 43075 9089 43076 9123
rect 42906 9076 43076 9089
rect 43278 9123 43448 9136
rect 43278 9089 43279 9123
rect 43279 9089 43447 9123
rect 43447 9089 43448 9123
rect 43278 9076 43448 9089
rect 43650 9123 43820 9136
rect 43650 9089 43651 9123
rect 43651 9089 43819 9123
rect 43819 9089 43820 9123
rect 43650 9076 43820 9089
rect 38070 8595 38240 8596
rect 38070 8561 38071 8595
rect 38071 8561 38239 8595
rect 38239 8561 38240 8595
rect 38070 8487 38240 8561
rect 38070 8453 38071 8487
rect 38071 8453 38239 8487
rect 38239 8453 38240 8487
rect 38070 8452 38240 8453
rect 38442 8595 38612 8596
rect 38442 8561 38443 8595
rect 38443 8561 38611 8595
rect 38611 8561 38612 8595
rect 38442 8487 38612 8561
rect 38442 8453 38443 8487
rect 38443 8453 38611 8487
rect 38611 8453 38612 8487
rect 38442 8452 38612 8453
rect 38814 8595 38984 8596
rect 38814 8561 38815 8595
rect 38815 8561 38983 8595
rect 38983 8561 38984 8595
rect 38814 8487 38984 8561
rect 38814 8453 38815 8487
rect 38815 8453 38983 8487
rect 38983 8453 38984 8487
rect 38814 8452 38984 8453
rect 39186 8595 39356 8596
rect 39186 8561 39187 8595
rect 39187 8561 39355 8595
rect 39355 8561 39356 8595
rect 39186 8487 39356 8561
rect 39186 8453 39187 8487
rect 39187 8453 39355 8487
rect 39355 8453 39356 8487
rect 39186 8452 39356 8453
rect 39558 8595 39728 8596
rect 39558 8561 39559 8595
rect 39559 8561 39727 8595
rect 39727 8561 39728 8595
rect 39558 8487 39728 8561
rect 39558 8453 39559 8487
rect 39559 8453 39727 8487
rect 39727 8453 39728 8487
rect 39558 8452 39728 8453
rect 39930 8595 40100 8596
rect 39930 8561 39931 8595
rect 39931 8561 40099 8595
rect 40099 8561 40100 8595
rect 39930 8487 40100 8561
rect 39930 8453 39931 8487
rect 39931 8453 40099 8487
rect 40099 8453 40100 8487
rect 39930 8452 40100 8453
rect 40302 8595 40472 8596
rect 40302 8561 40303 8595
rect 40303 8561 40471 8595
rect 40471 8561 40472 8595
rect 40302 8487 40472 8561
rect 40302 8453 40303 8487
rect 40303 8453 40471 8487
rect 40471 8453 40472 8487
rect 40302 8452 40472 8453
rect 40674 8595 40844 8596
rect 40674 8561 40675 8595
rect 40675 8561 40843 8595
rect 40843 8561 40844 8595
rect 40674 8487 40844 8561
rect 40674 8453 40675 8487
rect 40675 8453 40843 8487
rect 40843 8453 40844 8487
rect 40674 8452 40844 8453
rect 41046 8595 41216 8596
rect 41046 8561 41047 8595
rect 41047 8561 41215 8595
rect 41215 8561 41216 8595
rect 41046 8487 41216 8561
rect 41046 8453 41047 8487
rect 41047 8453 41215 8487
rect 41215 8453 41216 8487
rect 41046 8452 41216 8453
rect 41418 8595 41588 8596
rect 41418 8561 41419 8595
rect 41419 8561 41587 8595
rect 41587 8561 41588 8595
rect 41418 8487 41588 8561
rect 41418 8453 41419 8487
rect 41419 8453 41587 8487
rect 41587 8453 41588 8487
rect 41418 8452 41588 8453
rect 41790 8595 41960 8596
rect 41790 8561 41791 8595
rect 41791 8561 41959 8595
rect 41959 8561 41960 8595
rect 41790 8487 41960 8561
rect 41790 8453 41791 8487
rect 41791 8453 41959 8487
rect 41959 8453 41960 8487
rect 41790 8452 41960 8453
rect 42162 8595 42332 8596
rect 42162 8561 42163 8595
rect 42163 8561 42331 8595
rect 42331 8561 42332 8595
rect 42162 8487 42332 8561
rect 42162 8453 42163 8487
rect 42163 8453 42331 8487
rect 42331 8453 42332 8487
rect 42162 8452 42332 8453
rect 42534 8595 42704 8596
rect 42534 8561 42535 8595
rect 42535 8561 42703 8595
rect 42703 8561 42704 8595
rect 42534 8487 42704 8561
rect 42534 8453 42535 8487
rect 42535 8453 42703 8487
rect 42703 8453 42704 8487
rect 42534 8452 42704 8453
rect 42906 8595 43076 8596
rect 42906 8561 42907 8595
rect 42907 8561 43075 8595
rect 43075 8561 43076 8595
rect 42906 8487 43076 8561
rect 42906 8453 42907 8487
rect 42907 8453 43075 8487
rect 43075 8453 43076 8487
rect 42906 8452 43076 8453
rect 43278 8595 43448 8596
rect 43278 8561 43279 8595
rect 43279 8561 43447 8595
rect 43447 8561 43448 8595
rect 43278 8487 43448 8561
rect 43278 8453 43279 8487
rect 43279 8453 43447 8487
rect 43447 8453 43448 8487
rect 43278 8452 43448 8453
rect 43650 8595 43820 8596
rect 43650 8561 43651 8595
rect 43651 8561 43819 8595
rect 43819 8561 43820 8595
rect 43650 8487 43820 8561
rect 43650 8453 43651 8487
rect 43651 8453 43819 8487
rect 43819 8453 43820 8487
rect 43650 8452 43820 8453
rect 38070 7959 38240 7960
rect 38070 7925 38071 7959
rect 38071 7925 38239 7959
rect 38239 7925 38240 7959
rect 38070 7851 38240 7925
rect 38070 7817 38071 7851
rect 38071 7817 38239 7851
rect 38239 7817 38240 7851
rect 38070 7816 38240 7817
rect 38442 7959 38612 7960
rect 38442 7925 38443 7959
rect 38443 7925 38611 7959
rect 38611 7925 38612 7959
rect 38442 7851 38612 7925
rect 38442 7817 38443 7851
rect 38443 7817 38611 7851
rect 38611 7817 38612 7851
rect 38442 7816 38612 7817
rect 38814 7959 38984 7960
rect 38814 7925 38815 7959
rect 38815 7925 38983 7959
rect 38983 7925 38984 7959
rect 38814 7851 38984 7925
rect 38814 7817 38815 7851
rect 38815 7817 38983 7851
rect 38983 7817 38984 7851
rect 38814 7816 38984 7817
rect 39186 7959 39356 7960
rect 39186 7925 39187 7959
rect 39187 7925 39355 7959
rect 39355 7925 39356 7959
rect 39186 7851 39356 7925
rect 39186 7817 39187 7851
rect 39187 7817 39355 7851
rect 39355 7817 39356 7851
rect 39186 7816 39356 7817
rect 39558 7959 39728 7960
rect 39558 7925 39559 7959
rect 39559 7925 39727 7959
rect 39727 7925 39728 7959
rect 39558 7851 39728 7925
rect 39558 7817 39559 7851
rect 39559 7817 39727 7851
rect 39727 7817 39728 7851
rect 39558 7816 39728 7817
rect 39930 7959 40100 7960
rect 39930 7925 39931 7959
rect 39931 7925 40099 7959
rect 40099 7925 40100 7959
rect 39930 7851 40100 7925
rect 39930 7817 39931 7851
rect 39931 7817 40099 7851
rect 40099 7817 40100 7851
rect 39930 7816 40100 7817
rect 40302 7959 40472 7960
rect 40302 7925 40303 7959
rect 40303 7925 40471 7959
rect 40471 7925 40472 7959
rect 40302 7851 40472 7925
rect 40302 7817 40303 7851
rect 40303 7817 40471 7851
rect 40471 7817 40472 7851
rect 40302 7816 40472 7817
rect 40674 7959 40844 7960
rect 40674 7925 40675 7959
rect 40675 7925 40843 7959
rect 40843 7925 40844 7959
rect 40674 7851 40844 7925
rect 40674 7817 40675 7851
rect 40675 7817 40843 7851
rect 40843 7817 40844 7851
rect 40674 7816 40844 7817
rect 41046 7959 41216 7960
rect 41046 7925 41047 7959
rect 41047 7925 41215 7959
rect 41215 7925 41216 7959
rect 41046 7851 41216 7925
rect 41046 7817 41047 7851
rect 41047 7817 41215 7851
rect 41215 7817 41216 7851
rect 41046 7816 41216 7817
rect 41418 7959 41588 7960
rect 41418 7925 41419 7959
rect 41419 7925 41587 7959
rect 41587 7925 41588 7959
rect 41418 7851 41588 7925
rect 41418 7817 41419 7851
rect 41419 7817 41587 7851
rect 41587 7817 41588 7851
rect 41418 7816 41588 7817
rect 41790 7959 41960 7960
rect 41790 7925 41791 7959
rect 41791 7925 41959 7959
rect 41959 7925 41960 7959
rect 41790 7851 41960 7925
rect 41790 7817 41791 7851
rect 41791 7817 41959 7851
rect 41959 7817 41960 7851
rect 41790 7816 41960 7817
rect 42162 7959 42332 7960
rect 42162 7925 42163 7959
rect 42163 7925 42331 7959
rect 42331 7925 42332 7959
rect 42162 7851 42332 7925
rect 42162 7817 42163 7851
rect 42163 7817 42331 7851
rect 42331 7817 42332 7851
rect 42162 7816 42332 7817
rect 42534 7959 42704 7960
rect 42534 7925 42535 7959
rect 42535 7925 42703 7959
rect 42703 7925 42704 7959
rect 42534 7851 42704 7925
rect 42534 7817 42535 7851
rect 42535 7817 42703 7851
rect 42703 7817 42704 7851
rect 42534 7816 42704 7817
rect 42906 7959 43076 7960
rect 42906 7925 42907 7959
rect 42907 7925 43075 7959
rect 43075 7925 43076 7959
rect 42906 7851 43076 7925
rect 42906 7817 42907 7851
rect 42907 7817 43075 7851
rect 43075 7817 43076 7851
rect 42906 7816 43076 7817
rect 43278 7959 43448 7960
rect 43278 7925 43279 7959
rect 43279 7925 43447 7959
rect 43447 7925 43448 7959
rect 43278 7851 43448 7925
rect 43278 7817 43279 7851
rect 43279 7817 43447 7851
rect 43447 7817 43448 7851
rect 43278 7816 43448 7817
rect 43650 7959 43820 7960
rect 43650 7925 43651 7959
rect 43651 7925 43819 7959
rect 43819 7925 43820 7959
rect 43650 7851 43820 7925
rect 43650 7817 43651 7851
rect 43651 7817 43819 7851
rect 43819 7817 43820 7851
rect 43650 7816 43820 7817
rect 38070 7323 38240 7336
rect 38070 7289 38071 7323
rect 38071 7289 38239 7323
rect 38239 7289 38240 7323
rect 38070 7276 38240 7289
rect 38442 7323 38612 7336
rect 38442 7289 38443 7323
rect 38443 7289 38611 7323
rect 38611 7289 38612 7323
rect 38442 7276 38612 7289
rect 35702 6594 36308 7216
rect 38814 7323 38984 7336
rect 38814 7289 38815 7323
rect 38815 7289 38983 7323
rect 38983 7289 38984 7323
rect 38814 7276 38984 7289
rect 39186 7323 39356 7336
rect 39186 7289 39187 7323
rect 39187 7289 39355 7323
rect 39355 7289 39356 7323
rect 39186 7276 39356 7289
rect 39558 7323 39728 7336
rect 39558 7289 39559 7323
rect 39559 7289 39727 7323
rect 39727 7289 39728 7323
rect 39558 7276 39728 7289
rect 39930 7323 40100 7336
rect 39930 7289 39931 7323
rect 39931 7289 40099 7323
rect 40099 7289 40100 7323
rect 39930 7276 40100 7289
rect 40302 7323 40472 7336
rect 40302 7289 40303 7323
rect 40303 7289 40471 7323
rect 40471 7289 40472 7323
rect 40302 7276 40472 7289
rect 40674 7323 40844 7336
rect 40674 7289 40675 7323
rect 40675 7289 40843 7323
rect 40843 7289 40844 7323
rect 40674 7276 40844 7289
rect 41046 7323 41216 7336
rect 41046 7289 41047 7323
rect 41047 7289 41215 7323
rect 41215 7289 41216 7323
rect 41046 7276 41216 7289
rect 41418 7323 41588 7336
rect 41418 7289 41419 7323
rect 41419 7289 41587 7323
rect 41587 7289 41588 7323
rect 41418 7276 41588 7289
rect 41790 7323 41960 7336
rect 41790 7289 41791 7323
rect 41791 7289 41959 7323
rect 41959 7289 41960 7323
rect 41790 7276 41960 7289
rect 42162 7323 42332 7336
rect 42162 7289 42163 7323
rect 42163 7289 42331 7323
rect 42331 7289 42332 7323
rect 42162 7276 42332 7289
rect 42534 7323 42704 7336
rect 42534 7289 42535 7323
rect 42535 7289 42703 7323
rect 42703 7289 42704 7323
rect 42534 7276 42704 7289
rect 42906 7323 43076 7336
rect 42906 7289 42907 7323
rect 42907 7289 43075 7323
rect 43075 7289 43076 7323
rect 42906 7276 43076 7289
rect 44022 9123 44192 9136
rect 44022 9089 44023 9123
rect 44023 9089 44191 9123
rect 44191 9089 44192 9123
rect 44022 9076 44192 9089
rect 44394 9123 44564 9136
rect 44394 9089 44395 9123
rect 44395 9089 44563 9123
rect 44563 9089 44564 9123
rect 44394 9076 44564 9089
rect 44766 9123 44936 9136
rect 44766 9089 44767 9123
rect 44767 9089 44935 9123
rect 44935 9089 44936 9123
rect 44766 9076 44936 9089
rect 45138 9123 45308 9136
rect 45138 9089 45139 9123
rect 45139 9089 45307 9123
rect 45307 9089 45308 9123
rect 45138 9076 45308 9089
rect 45510 9123 45680 9136
rect 45510 9089 45511 9123
rect 45511 9089 45679 9123
rect 45679 9089 45680 9123
rect 45510 9076 45680 9089
rect 45882 9123 46052 9136
rect 45882 9089 45883 9123
rect 45883 9089 46051 9123
rect 46051 9089 46052 9123
rect 45882 9076 46052 9089
rect 46254 9123 46424 9136
rect 46254 9089 46255 9123
rect 46255 9089 46423 9123
rect 46423 9089 46424 9123
rect 46254 9076 46424 9089
rect 46626 9123 46796 9136
rect 46626 9089 46627 9123
rect 46627 9089 46795 9123
rect 46795 9089 46796 9123
rect 46626 9076 46796 9089
rect 46998 9123 47168 9136
rect 46998 9089 46999 9123
rect 46999 9089 47167 9123
rect 47167 9089 47168 9123
rect 46998 9076 47168 9089
rect 47370 9123 47540 9136
rect 47370 9089 47371 9123
rect 47371 9089 47539 9123
rect 47539 9089 47540 9123
rect 47370 9076 47540 9089
rect 47742 9123 47912 9136
rect 47742 9089 47743 9123
rect 47743 9089 47911 9123
rect 47911 9089 47912 9123
rect 47742 9076 47912 9089
rect 48114 9123 48284 9136
rect 48114 9089 48115 9123
rect 48115 9089 48283 9123
rect 48283 9089 48284 9123
rect 48114 9076 48284 9089
rect 48486 9123 48656 9136
rect 48486 9089 48487 9123
rect 48487 9089 48655 9123
rect 48655 9089 48656 9123
rect 48486 9076 48656 9089
rect 48858 9123 49028 9136
rect 48858 9089 48859 9123
rect 48859 9089 49027 9123
rect 49027 9089 49028 9123
rect 48858 9076 49028 9089
rect 49230 9123 49400 9136
rect 49230 9089 49231 9123
rect 49231 9089 49399 9123
rect 49399 9089 49400 9123
rect 49230 9076 49400 9089
rect 49602 9123 49772 9136
rect 49602 9089 49603 9123
rect 49603 9089 49771 9123
rect 49771 9089 49772 9123
rect 49602 9076 49772 9089
rect 44022 8595 44192 8596
rect 44022 8561 44023 8595
rect 44023 8561 44191 8595
rect 44191 8561 44192 8595
rect 44022 8487 44192 8561
rect 44022 8453 44023 8487
rect 44023 8453 44191 8487
rect 44191 8453 44192 8487
rect 44022 8452 44192 8453
rect 44394 8595 44564 8596
rect 44394 8561 44395 8595
rect 44395 8561 44563 8595
rect 44563 8561 44564 8595
rect 44394 8487 44564 8561
rect 44394 8453 44395 8487
rect 44395 8453 44563 8487
rect 44563 8453 44564 8487
rect 44394 8452 44564 8453
rect 44766 8595 44936 8596
rect 44766 8561 44767 8595
rect 44767 8561 44935 8595
rect 44935 8561 44936 8595
rect 44766 8487 44936 8561
rect 44766 8453 44767 8487
rect 44767 8453 44935 8487
rect 44935 8453 44936 8487
rect 44766 8452 44936 8453
rect 45138 8595 45308 8596
rect 45138 8561 45139 8595
rect 45139 8561 45307 8595
rect 45307 8561 45308 8595
rect 45138 8487 45308 8561
rect 45138 8453 45139 8487
rect 45139 8453 45307 8487
rect 45307 8453 45308 8487
rect 45138 8452 45308 8453
rect 45510 8595 45680 8596
rect 45510 8561 45511 8595
rect 45511 8561 45679 8595
rect 45679 8561 45680 8595
rect 45510 8487 45680 8561
rect 45510 8453 45511 8487
rect 45511 8453 45679 8487
rect 45679 8453 45680 8487
rect 45510 8452 45680 8453
rect 45882 8595 46052 8596
rect 45882 8561 45883 8595
rect 45883 8561 46051 8595
rect 46051 8561 46052 8595
rect 45882 8487 46052 8561
rect 45882 8453 45883 8487
rect 45883 8453 46051 8487
rect 46051 8453 46052 8487
rect 45882 8452 46052 8453
rect 46254 8595 46424 8596
rect 46254 8561 46255 8595
rect 46255 8561 46423 8595
rect 46423 8561 46424 8595
rect 46254 8487 46424 8561
rect 46254 8453 46255 8487
rect 46255 8453 46423 8487
rect 46423 8453 46424 8487
rect 46254 8452 46424 8453
rect 46626 8595 46796 8596
rect 46626 8561 46627 8595
rect 46627 8561 46795 8595
rect 46795 8561 46796 8595
rect 46626 8487 46796 8561
rect 46626 8453 46627 8487
rect 46627 8453 46795 8487
rect 46795 8453 46796 8487
rect 46626 8452 46796 8453
rect 46998 8595 47168 8596
rect 46998 8561 46999 8595
rect 46999 8561 47167 8595
rect 47167 8561 47168 8595
rect 46998 8487 47168 8561
rect 46998 8453 46999 8487
rect 46999 8453 47167 8487
rect 47167 8453 47168 8487
rect 46998 8452 47168 8453
rect 47370 8595 47540 8596
rect 47370 8561 47371 8595
rect 47371 8561 47539 8595
rect 47539 8561 47540 8595
rect 47370 8487 47540 8561
rect 47370 8453 47371 8487
rect 47371 8453 47539 8487
rect 47539 8453 47540 8487
rect 47370 8452 47540 8453
rect 47742 8595 47912 8596
rect 47742 8561 47743 8595
rect 47743 8561 47911 8595
rect 47911 8561 47912 8595
rect 47742 8487 47912 8561
rect 47742 8453 47743 8487
rect 47743 8453 47911 8487
rect 47911 8453 47912 8487
rect 47742 8452 47912 8453
rect 48114 8595 48284 8596
rect 48114 8561 48115 8595
rect 48115 8561 48283 8595
rect 48283 8561 48284 8595
rect 48114 8487 48284 8561
rect 48114 8453 48115 8487
rect 48115 8453 48283 8487
rect 48283 8453 48284 8487
rect 48114 8452 48284 8453
rect 48486 8595 48656 8596
rect 48486 8561 48487 8595
rect 48487 8561 48655 8595
rect 48655 8561 48656 8595
rect 48486 8487 48656 8561
rect 48486 8453 48487 8487
rect 48487 8453 48655 8487
rect 48655 8453 48656 8487
rect 48486 8452 48656 8453
rect 48858 8595 49028 8596
rect 48858 8561 48859 8595
rect 48859 8561 49027 8595
rect 49027 8561 49028 8595
rect 48858 8487 49028 8561
rect 48858 8453 48859 8487
rect 48859 8453 49027 8487
rect 49027 8453 49028 8487
rect 48858 8452 49028 8453
rect 49230 8595 49400 8596
rect 49230 8561 49231 8595
rect 49231 8561 49399 8595
rect 49399 8561 49400 8595
rect 49230 8487 49400 8561
rect 49230 8453 49231 8487
rect 49231 8453 49399 8487
rect 49399 8453 49400 8487
rect 49230 8452 49400 8453
rect 49602 8595 49772 8596
rect 49602 8561 49603 8595
rect 49603 8561 49771 8595
rect 49771 8561 49772 8595
rect 49602 8487 49772 8561
rect 49602 8453 49603 8487
rect 49603 8453 49771 8487
rect 49771 8453 49772 8487
rect 49602 8452 49772 8453
rect 44022 7959 44192 7960
rect 44022 7925 44023 7959
rect 44023 7925 44191 7959
rect 44191 7925 44192 7959
rect 44022 7851 44192 7925
rect 44022 7817 44023 7851
rect 44023 7817 44191 7851
rect 44191 7817 44192 7851
rect 44022 7816 44192 7817
rect 44394 7959 44564 7960
rect 44394 7925 44395 7959
rect 44395 7925 44563 7959
rect 44563 7925 44564 7959
rect 44394 7851 44564 7925
rect 44394 7817 44395 7851
rect 44395 7817 44563 7851
rect 44563 7817 44564 7851
rect 44394 7816 44564 7817
rect 44766 7959 44936 7960
rect 44766 7925 44767 7959
rect 44767 7925 44935 7959
rect 44935 7925 44936 7959
rect 44766 7851 44936 7925
rect 44766 7817 44767 7851
rect 44767 7817 44935 7851
rect 44935 7817 44936 7851
rect 44766 7816 44936 7817
rect 45138 7959 45308 7960
rect 45138 7925 45139 7959
rect 45139 7925 45307 7959
rect 45307 7925 45308 7959
rect 45138 7851 45308 7925
rect 45138 7817 45139 7851
rect 45139 7817 45307 7851
rect 45307 7817 45308 7851
rect 45138 7816 45308 7817
rect 45510 7959 45680 7960
rect 45510 7925 45511 7959
rect 45511 7925 45679 7959
rect 45679 7925 45680 7959
rect 45510 7851 45680 7925
rect 45510 7817 45511 7851
rect 45511 7817 45679 7851
rect 45679 7817 45680 7851
rect 45510 7816 45680 7817
rect 45882 7959 46052 7960
rect 45882 7925 45883 7959
rect 45883 7925 46051 7959
rect 46051 7925 46052 7959
rect 45882 7851 46052 7925
rect 45882 7817 45883 7851
rect 45883 7817 46051 7851
rect 46051 7817 46052 7851
rect 45882 7816 46052 7817
rect 46254 7959 46424 7960
rect 46254 7925 46255 7959
rect 46255 7925 46423 7959
rect 46423 7925 46424 7959
rect 46254 7851 46424 7925
rect 46254 7817 46255 7851
rect 46255 7817 46423 7851
rect 46423 7817 46424 7851
rect 46254 7816 46424 7817
rect 46626 7959 46796 7960
rect 46626 7925 46627 7959
rect 46627 7925 46795 7959
rect 46795 7925 46796 7959
rect 46626 7851 46796 7925
rect 46626 7817 46627 7851
rect 46627 7817 46795 7851
rect 46795 7817 46796 7851
rect 46626 7816 46796 7817
rect 46998 7959 47168 7960
rect 46998 7925 46999 7959
rect 46999 7925 47167 7959
rect 47167 7925 47168 7959
rect 46998 7851 47168 7925
rect 46998 7817 46999 7851
rect 46999 7817 47167 7851
rect 47167 7817 47168 7851
rect 46998 7816 47168 7817
rect 47370 7959 47540 7960
rect 47370 7925 47371 7959
rect 47371 7925 47539 7959
rect 47539 7925 47540 7959
rect 47370 7851 47540 7925
rect 47370 7817 47371 7851
rect 47371 7817 47539 7851
rect 47539 7817 47540 7851
rect 47370 7816 47540 7817
rect 47742 7959 47912 7960
rect 47742 7925 47743 7959
rect 47743 7925 47911 7959
rect 47911 7925 47912 7959
rect 47742 7851 47912 7925
rect 47742 7817 47743 7851
rect 47743 7817 47911 7851
rect 47911 7817 47912 7851
rect 47742 7816 47912 7817
rect 48114 7959 48284 7960
rect 48114 7925 48115 7959
rect 48115 7925 48283 7959
rect 48283 7925 48284 7959
rect 48114 7851 48284 7925
rect 48114 7817 48115 7851
rect 48115 7817 48283 7851
rect 48283 7817 48284 7851
rect 48114 7816 48284 7817
rect 48486 7959 48656 7960
rect 48486 7925 48487 7959
rect 48487 7925 48655 7959
rect 48655 7925 48656 7959
rect 48486 7851 48656 7925
rect 48486 7817 48487 7851
rect 48487 7817 48655 7851
rect 48655 7817 48656 7851
rect 48486 7816 48656 7817
rect 48858 7959 49028 7960
rect 48858 7925 48859 7959
rect 48859 7925 49027 7959
rect 49027 7925 49028 7959
rect 48858 7851 49028 7925
rect 48858 7817 48859 7851
rect 48859 7817 49027 7851
rect 49027 7817 49028 7851
rect 48858 7816 49028 7817
rect 49230 7959 49400 7960
rect 49230 7925 49231 7959
rect 49231 7925 49399 7959
rect 49399 7925 49400 7959
rect 49230 7851 49400 7925
rect 49230 7817 49231 7851
rect 49231 7817 49399 7851
rect 49399 7817 49400 7851
rect 49230 7816 49400 7817
rect 49602 7959 49772 7960
rect 49602 7925 49603 7959
rect 49603 7925 49771 7959
rect 49771 7925 49772 7959
rect 49602 7851 49772 7925
rect 49602 7817 49603 7851
rect 49603 7817 49771 7851
rect 49771 7817 49772 7851
rect 49602 7816 49772 7817
rect 43278 7323 43448 7336
rect 43278 7289 43279 7323
rect 43279 7289 43447 7323
rect 43447 7289 43448 7323
rect 43278 7276 43448 7289
rect 43650 7323 43820 7336
rect 43650 7289 43651 7323
rect 43651 7289 43819 7323
rect 43819 7289 43820 7323
rect 43650 7276 43820 7289
rect 44022 7323 44192 7336
rect 44022 7289 44023 7323
rect 44023 7289 44191 7323
rect 44191 7289 44192 7323
rect 44022 7276 44192 7289
rect 44394 7323 44564 7336
rect 44394 7289 44395 7323
rect 44395 7289 44563 7323
rect 44563 7289 44564 7323
rect 44394 7276 44564 7289
rect 44766 7323 44936 7336
rect 44766 7289 44767 7323
rect 44767 7289 44935 7323
rect 44935 7289 44936 7323
rect 44766 7276 44936 7289
rect 45138 7323 45308 7336
rect 45138 7289 45139 7323
rect 45139 7289 45307 7323
rect 45307 7289 45308 7323
rect 45138 7276 45308 7289
rect 45510 7323 45680 7336
rect 45510 7289 45511 7323
rect 45511 7289 45679 7323
rect 45679 7289 45680 7323
rect 45510 7276 45680 7289
rect 45882 7323 46052 7336
rect 45882 7289 45883 7323
rect 45883 7289 46051 7323
rect 46051 7289 46052 7323
rect 45882 7276 46052 7289
rect 46254 7323 46424 7336
rect 46254 7289 46255 7323
rect 46255 7289 46423 7323
rect 46423 7289 46424 7323
rect 46254 7276 46424 7289
rect 46626 7323 46796 7336
rect 46626 7289 46627 7323
rect 46627 7289 46795 7323
rect 46795 7289 46796 7323
rect 46626 7276 46796 7289
rect 46998 7323 47168 7336
rect 46998 7289 46999 7323
rect 46999 7289 47167 7323
rect 47167 7289 47168 7323
rect 46998 7276 47168 7289
rect 47370 7323 47540 7336
rect 47370 7289 47371 7323
rect 47371 7289 47539 7323
rect 47539 7289 47540 7323
rect 47370 7276 47540 7289
rect 47742 7323 47912 7336
rect 47742 7289 47743 7323
rect 47743 7289 47911 7323
rect 47911 7289 47912 7323
rect 47742 7276 47912 7289
rect 48114 7323 48284 7336
rect 48114 7289 48115 7323
rect 48115 7289 48283 7323
rect 48283 7289 48284 7323
rect 48114 7276 48284 7289
rect 48486 7323 48656 7336
rect 48486 7289 48487 7323
rect 48487 7289 48655 7323
rect 48655 7289 48656 7323
rect 48486 7276 48656 7289
rect 48858 7323 49028 7336
rect 48858 7289 48859 7323
rect 48859 7289 49027 7323
rect 49027 7289 49028 7323
rect 48858 7276 49028 7289
rect 49230 7323 49400 7336
rect 49230 7289 49231 7323
rect 49231 7289 49399 7323
rect 49399 7289 49400 7323
rect 49230 7276 49400 7289
rect 49602 7323 49772 7336
rect 49602 7289 49603 7323
rect 49603 7289 49771 7323
rect 49771 7289 49772 7323
rect 49602 7276 49772 7289
rect 39558 6735 39728 6750
rect 39558 6701 39559 6735
rect 39559 6701 39727 6735
rect 39727 6701 39728 6735
rect 39558 6686 39728 6701
rect 39930 6735 40100 6750
rect 39930 6701 39931 6735
rect 39931 6701 40099 6735
rect 40099 6701 40100 6735
rect 39930 6686 40100 6701
rect 40302 6735 40472 6750
rect 40302 6701 40303 6735
rect 40303 6701 40471 6735
rect 40471 6701 40472 6735
rect 40302 6686 40472 6701
rect 40674 6735 40844 6750
rect 40674 6701 40675 6735
rect 40675 6701 40843 6735
rect 40843 6701 40844 6735
rect 40674 6686 40844 6701
rect 41046 6735 41216 6750
rect 41046 6701 41047 6735
rect 41047 6701 41215 6735
rect 41215 6701 41216 6735
rect 41046 6686 41216 6701
rect 41418 6735 41588 6750
rect 41418 6701 41419 6735
rect 41419 6701 41587 6735
rect 41587 6701 41588 6735
rect 41418 6686 41588 6701
rect 41790 6735 41960 6750
rect 41790 6701 41791 6735
rect 41791 6701 41959 6735
rect 41959 6701 41960 6735
rect 41790 6686 41960 6701
rect 42162 6735 42332 6750
rect 42162 6701 42163 6735
rect 42163 6701 42331 6735
rect 42331 6701 42332 6735
rect 42162 6686 42332 6701
rect 44154 6696 44436 6968
rect 44898 6696 45180 6968
rect 45642 6696 45924 6968
rect 46386 6696 46668 6968
rect 47130 6696 47412 6968
rect 47874 6696 48156 6968
rect 48618 6696 48900 6968
rect 49362 6696 49644 6968
rect 39558 5807 39728 5808
rect 39558 5773 39559 5807
rect 39559 5773 39727 5807
rect 39727 5773 39728 5807
rect 39558 5699 39728 5773
rect 39558 5665 39559 5699
rect 39559 5665 39727 5699
rect 39727 5665 39728 5699
rect 39558 5664 39728 5665
rect 39930 5807 40100 5808
rect 39930 5773 39931 5807
rect 39931 5773 40099 5807
rect 40099 5773 40100 5807
rect 39930 5699 40100 5773
rect 39930 5665 39931 5699
rect 39931 5665 40099 5699
rect 40099 5665 40100 5699
rect 39930 5664 40100 5665
rect 40302 5807 40472 5808
rect 40302 5773 40303 5807
rect 40303 5773 40471 5807
rect 40471 5773 40472 5807
rect 40302 5699 40472 5773
rect 40302 5665 40303 5699
rect 40303 5665 40471 5699
rect 40471 5665 40472 5699
rect 40302 5664 40472 5665
rect 40674 5807 40844 5808
rect 40674 5773 40675 5807
rect 40675 5773 40843 5807
rect 40843 5773 40844 5807
rect 40674 5699 40844 5773
rect 40674 5665 40675 5699
rect 40675 5665 40843 5699
rect 40843 5665 40844 5699
rect 40674 5664 40844 5665
rect 41046 5807 41216 5808
rect 41046 5773 41047 5807
rect 41047 5773 41215 5807
rect 41215 5773 41216 5807
rect 41046 5699 41216 5773
rect 41046 5665 41047 5699
rect 41047 5665 41215 5699
rect 41215 5665 41216 5699
rect 41046 5664 41216 5665
rect 41418 5807 41588 5808
rect 41418 5773 41419 5807
rect 41419 5773 41587 5807
rect 41587 5773 41588 5807
rect 41418 5699 41588 5773
rect 41418 5665 41419 5699
rect 41419 5665 41587 5699
rect 41587 5665 41588 5699
rect 41418 5664 41588 5665
rect 41790 5807 41960 5808
rect 41790 5773 41791 5807
rect 41791 5773 41959 5807
rect 41959 5773 41960 5807
rect 41790 5699 41960 5773
rect 41790 5665 41791 5699
rect 41791 5665 41959 5699
rect 41959 5665 41960 5699
rect 41790 5664 41960 5665
rect 42162 5807 42332 5808
rect 42162 5773 42163 5807
rect 42163 5773 42331 5807
rect 42331 5773 42332 5807
rect 42162 5699 42332 5773
rect 42162 5665 42163 5699
rect 42163 5665 42331 5699
rect 42331 5665 42332 5699
rect 42162 5664 42332 5665
rect 43036 4980 43318 5252
rect 39558 4771 39728 4772
rect 39558 4737 39559 4771
rect 39559 4737 39727 4771
rect 39727 4737 39728 4771
rect 39558 4663 39728 4737
rect 39558 4629 39559 4663
rect 39559 4629 39727 4663
rect 39727 4629 39728 4663
rect 39558 4628 39728 4629
rect 39930 4771 40100 4772
rect 39930 4737 39931 4771
rect 39931 4737 40099 4771
rect 40099 4737 40100 4771
rect 39930 4663 40100 4737
rect 39930 4629 39931 4663
rect 39931 4629 40099 4663
rect 40099 4629 40100 4663
rect 39930 4628 40100 4629
rect 40302 4771 40472 4772
rect 40302 4737 40303 4771
rect 40303 4737 40471 4771
rect 40471 4737 40472 4771
rect 40302 4663 40472 4737
rect 40302 4629 40303 4663
rect 40303 4629 40471 4663
rect 40471 4629 40472 4663
rect 40302 4628 40472 4629
rect 40674 4771 40844 4772
rect 40674 4737 40675 4771
rect 40675 4737 40843 4771
rect 40843 4737 40844 4771
rect 40674 4663 40844 4737
rect 40674 4629 40675 4663
rect 40675 4629 40843 4663
rect 40843 4629 40844 4663
rect 40674 4628 40844 4629
rect 41046 4771 41216 4772
rect 41046 4737 41047 4771
rect 41047 4737 41215 4771
rect 41215 4737 41216 4771
rect 41046 4663 41216 4737
rect 41046 4629 41047 4663
rect 41047 4629 41215 4663
rect 41215 4629 41216 4663
rect 41046 4628 41216 4629
rect 41418 4771 41588 4772
rect 41418 4737 41419 4771
rect 41419 4737 41587 4771
rect 41587 4737 41588 4771
rect 41418 4663 41588 4737
rect 41418 4629 41419 4663
rect 41419 4629 41587 4663
rect 41587 4629 41588 4663
rect 41418 4628 41588 4629
rect 41790 4771 41960 4772
rect 41790 4737 41791 4771
rect 41791 4737 41959 4771
rect 41959 4737 41960 4771
rect 41790 4663 41960 4737
rect 41790 4629 41791 4663
rect 41791 4629 41959 4663
rect 41959 4629 41960 4663
rect 41790 4628 41960 4629
rect 42162 4771 42332 4772
rect 42162 4737 42163 4771
rect 42163 4737 42331 4771
rect 42331 4737 42332 4771
rect 42162 4663 42332 4737
rect 42162 4629 42163 4663
rect 42163 4629 42331 4663
rect 42331 4629 42332 4663
rect 42162 4628 42332 4629
rect 43460 4548 43612 4712
rect 43460 4148 43612 4312
rect 39558 3735 39728 3736
rect 39558 3701 39559 3735
rect 39559 3701 39727 3735
rect 39727 3701 39728 3735
rect 39558 3627 39728 3701
rect 39558 3593 39559 3627
rect 39559 3593 39727 3627
rect 39727 3593 39728 3627
rect 39558 3592 39728 3593
rect 39930 3735 40100 3736
rect 39930 3701 39931 3735
rect 39931 3701 40099 3735
rect 40099 3701 40100 3735
rect 39930 3627 40100 3701
rect 39930 3593 39931 3627
rect 39931 3593 40099 3627
rect 40099 3593 40100 3627
rect 39930 3592 40100 3593
rect 40302 3735 40472 3736
rect 40302 3701 40303 3735
rect 40303 3701 40471 3735
rect 40471 3701 40472 3735
rect 40302 3627 40472 3701
rect 40302 3593 40303 3627
rect 40303 3593 40471 3627
rect 40471 3593 40472 3627
rect 40302 3592 40472 3593
rect 40674 3735 40844 3736
rect 40674 3701 40675 3735
rect 40675 3701 40843 3735
rect 40843 3701 40844 3735
rect 40674 3627 40844 3701
rect 40674 3593 40675 3627
rect 40675 3593 40843 3627
rect 40843 3593 40844 3627
rect 40674 3592 40844 3593
rect 41046 3735 41216 3736
rect 41046 3701 41047 3735
rect 41047 3701 41215 3735
rect 41215 3701 41216 3735
rect 41046 3627 41216 3701
rect 41046 3593 41047 3627
rect 41047 3593 41215 3627
rect 41215 3593 41216 3627
rect 41046 3592 41216 3593
rect 41418 3735 41588 3736
rect 41418 3701 41419 3735
rect 41419 3701 41587 3735
rect 41587 3701 41588 3735
rect 41418 3627 41588 3701
rect 41418 3593 41419 3627
rect 41419 3593 41587 3627
rect 41587 3593 41588 3627
rect 41418 3592 41588 3593
rect 41790 3735 41960 3736
rect 41790 3701 41791 3735
rect 41791 3701 41959 3735
rect 41959 3701 41960 3735
rect 41790 3627 41960 3701
rect 41790 3593 41791 3627
rect 41791 3593 41959 3627
rect 41959 3593 41960 3627
rect 41790 3592 41960 3593
rect 42162 3735 42332 3736
rect 42162 3701 42163 3735
rect 42163 3701 42331 3735
rect 42331 3701 42332 3735
rect 42162 3627 42332 3701
rect 42162 3593 42163 3627
rect 42163 3593 42331 3627
rect 42331 3593 42332 3627
rect 42162 3592 42332 3593
rect 43460 3748 43612 3912
rect 39558 2699 39728 2710
rect 39558 2665 39559 2699
rect 39559 2665 39727 2699
rect 39727 2665 39728 2699
rect 39558 2656 39728 2665
rect 39930 2699 40100 2710
rect 39930 2665 39931 2699
rect 39931 2665 40099 2699
rect 40099 2665 40100 2699
rect 39930 2656 40100 2665
rect 40302 2699 40472 2710
rect 40302 2665 40303 2699
rect 40303 2665 40471 2699
rect 40471 2665 40472 2699
rect 40302 2656 40472 2665
rect 40674 2699 40844 2710
rect 40674 2665 40675 2699
rect 40675 2665 40843 2699
rect 40843 2665 40844 2699
rect 40674 2656 40844 2665
rect 41046 2699 41216 2710
rect 41046 2665 41047 2699
rect 41047 2665 41215 2699
rect 41215 2665 41216 2699
rect 41046 2656 41216 2665
rect 41418 2699 41588 2710
rect 41418 2665 41419 2699
rect 41419 2665 41587 2699
rect 41587 2665 41588 2699
rect 41418 2656 41588 2665
rect 41790 2699 41960 2710
rect 41790 2665 41791 2699
rect 41791 2665 41959 2699
rect 41959 2665 41960 2699
rect 41790 2656 41960 2665
rect 40538 2190 41352 2370
rect 39558 2041 39728 2052
rect 39558 2007 39559 2041
rect 39559 2007 39727 2041
rect 39727 2007 39728 2041
rect 39558 1996 39728 2007
rect 39930 2041 40100 2052
rect 39930 2007 39931 2041
rect 39931 2007 40099 2041
rect 40099 2007 40100 2041
rect 39930 1996 40100 2007
rect 40302 2041 40472 2052
rect 40302 2007 40303 2041
rect 40303 2007 40471 2041
rect 40471 2007 40472 2041
rect 40302 1996 40472 2007
rect 40674 2041 40844 2052
rect 40674 2007 40675 2041
rect 40675 2007 40843 2041
rect 40843 2007 40844 2041
rect 40674 1996 40844 2007
rect 41046 2041 41216 2052
rect 41046 2007 41047 2041
rect 41047 2007 41215 2041
rect 41215 2007 41216 2041
rect 41046 1996 41216 2007
rect 42162 2699 42332 2710
rect 42162 2665 42163 2699
rect 42163 2665 42331 2699
rect 42331 2665 42332 2699
rect 42162 2656 42332 2665
rect 42664 2514 42946 2786
rect 41418 2041 41588 2052
rect 41418 2007 41419 2041
rect 41419 2007 41587 2041
rect 41587 2007 41588 2041
rect 41418 1996 41588 2007
rect 41790 2041 41960 2052
rect 41790 2007 41791 2041
rect 41791 2007 41959 2041
rect 41959 2007 41960 2041
rect 41790 1996 41960 2007
rect 42162 2041 42332 2052
rect 42162 2007 42163 2041
rect 42163 2007 42331 2041
rect 42331 2007 42332 2041
rect 42162 1996 42332 2007
rect 42534 2041 42704 2052
rect 42534 2007 42535 2041
rect 42535 2007 42703 2041
rect 42703 2007 42704 2041
rect 42534 1996 42704 2007
rect 43460 3348 43612 3512
rect 43408 2514 43690 2786
rect 44152 2514 44434 2786
rect 44896 2514 45178 2786
rect 45640 2514 45922 2786
rect 46384 2514 46666 2786
rect 47128 2514 47410 2786
rect 47872 2514 48154 2786
rect 43044 2190 43294 2440
rect 42906 2041 43076 2052
rect 42906 2007 42907 2041
rect 42907 2007 43075 2041
rect 43075 2007 43076 2041
rect 42906 1996 43076 2007
rect 43278 2041 43448 2052
rect 43278 2007 43279 2041
rect 43279 2007 43447 2041
rect 43447 2007 43448 2041
rect 43278 1996 43448 2007
rect 43650 2041 43820 2052
rect 43650 2007 43651 2041
rect 43651 2007 43819 2041
rect 43819 2007 43820 2041
rect 43650 1996 43820 2007
rect 44022 2041 44192 2052
rect 44022 2007 44023 2041
rect 44023 2007 44191 2041
rect 44191 2007 44192 2041
rect 44022 1996 44192 2007
rect 44394 2041 44564 2052
rect 44394 2007 44395 2041
rect 44395 2007 44563 2041
rect 44563 2007 44564 2041
rect 44394 1996 44564 2007
rect 44766 2041 44936 2052
rect 44766 2007 44767 2041
rect 44767 2007 44935 2041
rect 44935 2007 44936 2041
rect 44766 1996 44936 2007
rect 45138 2041 45308 2052
rect 45138 2007 45139 2041
rect 45139 2007 45307 2041
rect 45307 2007 45308 2041
rect 45138 1996 45308 2007
rect 45510 2041 45680 2052
rect 45510 2007 45511 2041
rect 45511 2007 45679 2041
rect 45679 2007 45680 2041
rect 45510 1996 45680 2007
rect 45882 2041 46052 2052
rect 45882 2007 45883 2041
rect 45883 2007 46051 2041
rect 46051 2007 46052 2041
rect 45882 1996 46052 2007
rect 46254 2041 46424 2052
rect 46254 2007 46255 2041
rect 46255 2007 46423 2041
rect 46423 2007 46424 2041
rect 46254 1996 46424 2007
rect 46626 2041 46796 2052
rect 46626 2007 46627 2041
rect 46627 2007 46795 2041
rect 46795 2007 46796 2041
rect 46626 1996 46796 2007
rect 46998 2041 47168 2052
rect 46998 2007 46999 2041
rect 46999 2007 47167 2041
rect 47167 2007 47168 2041
rect 46998 1996 47168 2007
rect 47370 2041 47540 2052
rect 47370 2007 47371 2041
rect 47371 2007 47539 2041
rect 47539 2007 47540 2041
rect 47370 1996 47540 2007
rect 47742 2041 47912 2052
rect 47742 2007 47743 2041
rect 47743 2007 47911 2041
rect 47911 2007 47912 2041
rect 47742 1996 47912 2007
rect 48114 2041 48284 2052
rect 48114 2007 48115 2041
rect 48115 2007 48283 2041
rect 48283 2007 48284 2041
rect 48114 1996 48284 2007
rect 39558 1731 39728 1732
rect 39558 1697 39559 1731
rect 39559 1697 39727 1731
rect 39727 1697 39728 1731
rect 39558 1623 39728 1697
rect 39558 1589 39559 1623
rect 39559 1589 39727 1623
rect 39727 1589 39728 1623
rect 39558 1588 39728 1589
rect 39930 1731 40100 1732
rect 39930 1697 39931 1731
rect 39931 1697 40099 1731
rect 40099 1697 40100 1731
rect 39930 1623 40100 1697
rect 39930 1589 39931 1623
rect 39931 1589 40099 1623
rect 40099 1589 40100 1623
rect 39930 1588 40100 1589
rect 40302 1731 40472 1732
rect 40302 1697 40303 1731
rect 40303 1697 40471 1731
rect 40471 1697 40472 1731
rect 40302 1623 40472 1697
rect 40302 1589 40303 1623
rect 40303 1589 40471 1623
rect 40471 1589 40472 1623
rect 40302 1588 40472 1589
rect 40674 1731 40844 1732
rect 40674 1697 40675 1731
rect 40675 1697 40843 1731
rect 40843 1697 40844 1731
rect 40674 1623 40844 1697
rect 40674 1589 40675 1623
rect 40675 1589 40843 1623
rect 40843 1589 40844 1623
rect 40674 1588 40844 1589
rect 41046 1731 41216 1732
rect 41046 1697 41047 1731
rect 41047 1697 41215 1731
rect 41215 1697 41216 1731
rect 41046 1623 41216 1697
rect 41046 1589 41047 1623
rect 41047 1589 41215 1623
rect 41215 1589 41216 1623
rect 41046 1588 41216 1589
rect 41418 1731 41588 1732
rect 41418 1697 41419 1731
rect 41419 1697 41587 1731
rect 41587 1697 41588 1731
rect 41418 1623 41588 1697
rect 41418 1589 41419 1623
rect 41419 1589 41587 1623
rect 41587 1589 41588 1623
rect 41418 1588 41588 1589
rect 41790 1731 41960 1732
rect 41790 1697 41791 1731
rect 41791 1697 41959 1731
rect 41959 1697 41960 1731
rect 41790 1623 41960 1697
rect 41790 1589 41791 1623
rect 41791 1589 41959 1623
rect 41959 1589 41960 1623
rect 41790 1588 41960 1589
rect 42162 1731 42332 1732
rect 42162 1697 42163 1731
rect 42163 1697 42331 1731
rect 42331 1697 42332 1731
rect 42162 1623 42332 1697
rect 42162 1589 42163 1623
rect 42163 1589 42331 1623
rect 42331 1589 42332 1623
rect 42162 1588 42332 1589
rect 42534 1731 42704 1732
rect 42534 1697 42535 1731
rect 42535 1697 42703 1731
rect 42703 1697 42704 1731
rect 42534 1623 42704 1697
rect 42534 1589 42535 1623
rect 42535 1589 42703 1623
rect 42703 1589 42704 1623
rect 42534 1588 42704 1589
rect 42906 1731 43076 1732
rect 42906 1697 42907 1731
rect 42907 1697 43075 1731
rect 43075 1697 43076 1731
rect 42906 1623 43076 1697
rect 42906 1589 42907 1623
rect 42907 1589 43075 1623
rect 43075 1589 43076 1623
rect 42906 1588 43076 1589
rect 43278 1731 43448 1732
rect 43278 1697 43279 1731
rect 43279 1697 43447 1731
rect 43447 1697 43448 1731
rect 43278 1623 43448 1697
rect 43278 1589 43279 1623
rect 43279 1589 43447 1623
rect 43447 1589 43448 1623
rect 43278 1588 43448 1589
rect 43650 1731 43820 1732
rect 43650 1697 43651 1731
rect 43651 1697 43819 1731
rect 43819 1697 43820 1731
rect 43650 1623 43820 1697
rect 43650 1589 43651 1623
rect 43651 1589 43819 1623
rect 43819 1589 43820 1623
rect 43650 1588 43820 1589
rect 44022 1731 44192 1732
rect 44022 1697 44023 1731
rect 44023 1697 44191 1731
rect 44191 1697 44192 1731
rect 44022 1623 44192 1697
rect 44022 1589 44023 1623
rect 44023 1589 44191 1623
rect 44191 1589 44192 1623
rect 44022 1588 44192 1589
rect 44394 1731 44564 1732
rect 44394 1697 44395 1731
rect 44395 1697 44563 1731
rect 44563 1697 44564 1731
rect 44394 1623 44564 1697
rect 44394 1589 44395 1623
rect 44395 1589 44563 1623
rect 44563 1589 44564 1623
rect 44394 1588 44564 1589
rect 44766 1731 44936 1732
rect 44766 1697 44767 1731
rect 44767 1697 44935 1731
rect 44935 1697 44936 1731
rect 44766 1623 44936 1697
rect 44766 1589 44767 1623
rect 44767 1589 44935 1623
rect 44935 1589 44936 1623
rect 44766 1588 44936 1589
rect 45138 1731 45308 1732
rect 45138 1697 45139 1731
rect 45139 1697 45307 1731
rect 45307 1697 45308 1731
rect 45138 1623 45308 1697
rect 45138 1589 45139 1623
rect 45139 1589 45307 1623
rect 45307 1589 45308 1623
rect 45138 1588 45308 1589
rect 45510 1731 45680 1732
rect 45510 1697 45511 1731
rect 45511 1697 45679 1731
rect 45679 1697 45680 1731
rect 45510 1623 45680 1697
rect 45510 1589 45511 1623
rect 45511 1589 45679 1623
rect 45679 1589 45680 1623
rect 45510 1588 45680 1589
rect 45882 1731 46052 1732
rect 45882 1697 45883 1731
rect 45883 1697 46051 1731
rect 46051 1697 46052 1731
rect 45882 1623 46052 1697
rect 45882 1589 45883 1623
rect 45883 1589 46051 1623
rect 46051 1589 46052 1623
rect 45882 1588 46052 1589
rect 46254 1731 46424 1732
rect 46254 1697 46255 1731
rect 46255 1697 46423 1731
rect 46423 1697 46424 1731
rect 46254 1623 46424 1697
rect 46254 1589 46255 1623
rect 46255 1589 46423 1623
rect 46423 1589 46424 1623
rect 46254 1588 46424 1589
rect 46626 1731 46796 1732
rect 46626 1697 46627 1731
rect 46627 1697 46795 1731
rect 46795 1697 46796 1731
rect 46626 1623 46796 1697
rect 46626 1589 46627 1623
rect 46627 1589 46795 1623
rect 46795 1589 46796 1623
rect 46626 1588 46796 1589
rect 46998 1731 47168 1732
rect 46998 1697 46999 1731
rect 46999 1697 47167 1731
rect 47167 1697 47168 1731
rect 46998 1623 47168 1697
rect 46998 1589 46999 1623
rect 46999 1589 47167 1623
rect 47167 1589 47168 1623
rect 46998 1588 47168 1589
rect 47370 1731 47540 1732
rect 47370 1697 47371 1731
rect 47371 1697 47539 1731
rect 47539 1697 47540 1731
rect 47370 1623 47540 1697
rect 47370 1589 47371 1623
rect 47371 1589 47539 1623
rect 47539 1589 47540 1623
rect 47370 1588 47540 1589
rect 47742 1731 47912 1732
rect 47742 1697 47743 1731
rect 47743 1697 47911 1731
rect 47911 1697 47912 1731
rect 47742 1623 47912 1697
rect 47742 1589 47743 1623
rect 47743 1589 47911 1623
rect 47911 1589 47912 1623
rect 47742 1588 47912 1589
rect 48114 1731 48284 1732
rect 48114 1697 48115 1731
rect 48115 1697 48283 1731
rect 48283 1697 48284 1731
rect 48114 1623 48284 1697
rect 48114 1589 48115 1623
rect 48115 1589 48283 1623
rect 48283 1589 48284 1623
rect 48114 1588 48284 1589
rect 39558 1313 39728 1314
rect 39558 1279 39559 1313
rect 39559 1279 39727 1313
rect 39727 1279 39728 1313
rect 39558 1205 39728 1279
rect 39558 1171 39559 1205
rect 39559 1171 39727 1205
rect 39727 1171 39728 1205
rect 39558 1170 39728 1171
rect 39930 1313 40100 1314
rect 39930 1279 39931 1313
rect 39931 1279 40099 1313
rect 40099 1279 40100 1313
rect 39930 1205 40100 1279
rect 39930 1171 39931 1205
rect 39931 1171 40099 1205
rect 40099 1171 40100 1205
rect 39930 1170 40100 1171
rect 40302 1313 40472 1314
rect 40302 1279 40303 1313
rect 40303 1279 40471 1313
rect 40471 1279 40472 1313
rect 40302 1205 40472 1279
rect 40302 1171 40303 1205
rect 40303 1171 40471 1205
rect 40471 1171 40472 1205
rect 40302 1170 40472 1171
rect 40674 1313 40844 1314
rect 40674 1279 40675 1313
rect 40675 1279 40843 1313
rect 40843 1279 40844 1313
rect 40674 1205 40844 1279
rect 40674 1171 40675 1205
rect 40675 1171 40843 1205
rect 40843 1171 40844 1205
rect 40674 1170 40844 1171
rect 41046 1313 41216 1314
rect 41046 1279 41047 1313
rect 41047 1279 41215 1313
rect 41215 1279 41216 1313
rect 41046 1205 41216 1279
rect 41046 1171 41047 1205
rect 41047 1171 41215 1205
rect 41215 1171 41216 1205
rect 41046 1170 41216 1171
rect 41418 1313 41588 1314
rect 41418 1279 41419 1313
rect 41419 1279 41587 1313
rect 41587 1279 41588 1313
rect 41418 1205 41588 1279
rect 41418 1171 41419 1205
rect 41419 1171 41587 1205
rect 41587 1171 41588 1205
rect 41418 1170 41588 1171
rect 41790 1313 41960 1314
rect 41790 1279 41791 1313
rect 41791 1279 41959 1313
rect 41959 1279 41960 1313
rect 41790 1205 41960 1279
rect 41790 1171 41791 1205
rect 41791 1171 41959 1205
rect 41959 1171 41960 1205
rect 41790 1170 41960 1171
rect 42162 1313 42332 1314
rect 42162 1279 42163 1313
rect 42163 1279 42331 1313
rect 42331 1279 42332 1313
rect 42162 1205 42332 1279
rect 42162 1171 42163 1205
rect 42163 1171 42331 1205
rect 42331 1171 42332 1205
rect 42162 1170 42332 1171
rect 42534 1313 42704 1314
rect 42534 1279 42535 1313
rect 42535 1279 42703 1313
rect 42703 1279 42704 1313
rect 42534 1205 42704 1279
rect 42534 1171 42535 1205
rect 42535 1171 42703 1205
rect 42703 1171 42704 1205
rect 42534 1170 42704 1171
rect 42906 1313 43076 1314
rect 42906 1279 42907 1313
rect 42907 1279 43075 1313
rect 43075 1279 43076 1313
rect 42906 1205 43076 1279
rect 42906 1171 42907 1205
rect 42907 1171 43075 1205
rect 43075 1171 43076 1205
rect 42906 1170 43076 1171
rect 43278 1313 43448 1314
rect 43278 1279 43279 1313
rect 43279 1279 43447 1313
rect 43447 1279 43448 1313
rect 43278 1205 43448 1279
rect 43278 1171 43279 1205
rect 43279 1171 43447 1205
rect 43447 1171 43448 1205
rect 43278 1170 43448 1171
rect 43650 1313 43820 1314
rect 43650 1279 43651 1313
rect 43651 1279 43819 1313
rect 43819 1279 43820 1313
rect 43650 1205 43820 1279
rect 43650 1171 43651 1205
rect 43651 1171 43819 1205
rect 43819 1171 43820 1205
rect 43650 1170 43820 1171
rect 44022 1313 44192 1314
rect 44022 1279 44023 1313
rect 44023 1279 44191 1313
rect 44191 1279 44192 1313
rect 44022 1205 44192 1279
rect 44022 1171 44023 1205
rect 44023 1171 44191 1205
rect 44191 1171 44192 1205
rect 44022 1170 44192 1171
rect 44394 1313 44564 1314
rect 44394 1279 44395 1313
rect 44395 1279 44563 1313
rect 44563 1279 44564 1313
rect 44394 1205 44564 1279
rect 44394 1171 44395 1205
rect 44395 1171 44563 1205
rect 44563 1171 44564 1205
rect 44394 1170 44564 1171
rect 44766 1313 44936 1314
rect 44766 1279 44767 1313
rect 44767 1279 44935 1313
rect 44935 1279 44936 1313
rect 44766 1205 44936 1279
rect 44766 1171 44767 1205
rect 44767 1171 44935 1205
rect 44935 1171 44936 1205
rect 44766 1170 44936 1171
rect 45138 1313 45308 1314
rect 45138 1279 45139 1313
rect 45139 1279 45307 1313
rect 45307 1279 45308 1313
rect 45138 1205 45308 1279
rect 45138 1171 45139 1205
rect 45139 1171 45307 1205
rect 45307 1171 45308 1205
rect 45138 1170 45308 1171
rect 45510 1313 45680 1314
rect 45510 1279 45511 1313
rect 45511 1279 45679 1313
rect 45679 1279 45680 1313
rect 45510 1205 45680 1279
rect 45510 1171 45511 1205
rect 45511 1171 45679 1205
rect 45679 1171 45680 1205
rect 45510 1170 45680 1171
rect 45882 1313 46052 1314
rect 45882 1279 45883 1313
rect 45883 1279 46051 1313
rect 46051 1279 46052 1313
rect 45882 1205 46052 1279
rect 45882 1171 45883 1205
rect 45883 1171 46051 1205
rect 46051 1171 46052 1205
rect 45882 1170 46052 1171
rect 46254 1313 46424 1314
rect 46254 1279 46255 1313
rect 46255 1279 46423 1313
rect 46423 1279 46424 1313
rect 46254 1205 46424 1279
rect 46254 1171 46255 1205
rect 46255 1171 46423 1205
rect 46423 1171 46424 1205
rect 46254 1170 46424 1171
rect 46626 1313 46796 1314
rect 46626 1279 46627 1313
rect 46627 1279 46795 1313
rect 46795 1279 46796 1313
rect 46626 1205 46796 1279
rect 46626 1171 46627 1205
rect 46627 1171 46795 1205
rect 46795 1171 46796 1205
rect 46626 1170 46796 1171
rect 46998 1313 47168 1314
rect 46998 1279 46999 1313
rect 46999 1279 47167 1313
rect 47167 1279 47168 1313
rect 46998 1205 47168 1279
rect 46998 1171 46999 1205
rect 46999 1171 47167 1205
rect 47167 1171 47168 1205
rect 46998 1170 47168 1171
rect 47370 1313 47540 1314
rect 47370 1279 47371 1313
rect 47371 1279 47539 1313
rect 47539 1279 47540 1313
rect 47370 1205 47540 1279
rect 47370 1171 47371 1205
rect 47371 1171 47539 1205
rect 47539 1171 47540 1205
rect 47370 1170 47540 1171
rect 47742 1313 47912 1314
rect 47742 1279 47743 1313
rect 47743 1279 47911 1313
rect 47911 1279 47912 1313
rect 47742 1205 47912 1279
rect 47742 1171 47743 1205
rect 47743 1171 47911 1205
rect 47911 1171 47912 1205
rect 47742 1170 47912 1171
rect 48114 1313 48284 1314
rect 48114 1279 48115 1313
rect 48115 1279 48283 1313
rect 48283 1279 48284 1313
rect 48114 1205 48284 1279
rect 48114 1171 48115 1205
rect 48115 1171 48283 1205
rect 48283 1171 48284 1205
rect 48114 1170 48284 1171
rect 39558 895 39728 896
rect 39558 861 39559 895
rect 39559 861 39727 895
rect 39727 861 39728 895
rect 39558 787 39728 861
rect 39558 753 39559 787
rect 39559 753 39727 787
rect 39727 753 39728 787
rect 39558 752 39728 753
rect 39930 895 40100 896
rect 39930 861 39931 895
rect 39931 861 40099 895
rect 40099 861 40100 895
rect 39930 787 40100 861
rect 39930 753 39931 787
rect 39931 753 40099 787
rect 40099 753 40100 787
rect 39930 752 40100 753
rect 40302 895 40472 896
rect 40302 861 40303 895
rect 40303 861 40471 895
rect 40471 861 40472 895
rect 40302 787 40472 861
rect 40302 753 40303 787
rect 40303 753 40471 787
rect 40471 753 40472 787
rect 40302 752 40472 753
rect 40674 895 40844 896
rect 40674 861 40675 895
rect 40675 861 40843 895
rect 40843 861 40844 895
rect 40674 787 40844 861
rect 40674 753 40675 787
rect 40675 753 40843 787
rect 40843 753 40844 787
rect 40674 752 40844 753
rect 41046 895 41216 896
rect 41046 861 41047 895
rect 41047 861 41215 895
rect 41215 861 41216 895
rect 41046 787 41216 861
rect 41046 753 41047 787
rect 41047 753 41215 787
rect 41215 753 41216 787
rect 41046 752 41216 753
rect 41418 895 41588 896
rect 41418 861 41419 895
rect 41419 861 41587 895
rect 41587 861 41588 895
rect 41418 787 41588 861
rect 41418 753 41419 787
rect 41419 753 41587 787
rect 41587 753 41588 787
rect 41418 752 41588 753
rect 41790 895 41960 896
rect 41790 861 41791 895
rect 41791 861 41959 895
rect 41959 861 41960 895
rect 41790 787 41960 861
rect 41790 753 41791 787
rect 41791 753 41959 787
rect 41959 753 41960 787
rect 41790 752 41960 753
rect 42162 895 42332 896
rect 42162 861 42163 895
rect 42163 861 42331 895
rect 42331 861 42332 895
rect 42162 787 42332 861
rect 42162 753 42163 787
rect 42163 753 42331 787
rect 42331 753 42332 787
rect 42162 752 42332 753
rect 42534 895 42704 896
rect 42534 861 42535 895
rect 42535 861 42703 895
rect 42703 861 42704 895
rect 42534 787 42704 861
rect 42534 753 42535 787
rect 42535 753 42703 787
rect 42703 753 42704 787
rect 42534 752 42704 753
rect 42906 895 43076 896
rect 42906 861 42907 895
rect 42907 861 43075 895
rect 43075 861 43076 895
rect 42906 787 43076 861
rect 42906 753 42907 787
rect 42907 753 43075 787
rect 43075 753 43076 787
rect 42906 752 43076 753
rect 43278 895 43448 896
rect 43278 861 43279 895
rect 43279 861 43447 895
rect 43447 861 43448 895
rect 43278 787 43448 861
rect 43278 753 43279 787
rect 43279 753 43447 787
rect 43447 753 43448 787
rect 43278 752 43448 753
rect 43650 895 43820 896
rect 43650 861 43651 895
rect 43651 861 43819 895
rect 43819 861 43820 895
rect 43650 787 43820 861
rect 43650 753 43651 787
rect 43651 753 43819 787
rect 43819 753 43820 787
rect 43650 752 43820 753
rect 44022 895 44192 896
rect 44022 861 44023 895
rect 44023 861 44191 895
rect 44191 861 44192 895
rect 44022 787 44192 861
rect 44022 753 44023 787
rect 44023 753 44191 787
rect 44191 753 44192 787
rect 44022 752 44192 753
rect 44394 895 44564 896
rect 44394 861 44395 895
rect 44395 861 44563 895
rect 44563 861 44564 895
rect 44394 787 44564 861
rect 44394 753 44395 787
rect 44395 753 44563 787
rect 44563 753 44564 787
rect 44394 752 44564 753
rect 44766 895 44936 896
rect 44766 861 44767 895
rect 44767 861 44935 895
rect 44935 861 44936 895
rect 44766 787 44936 861
rect 44766 753 44767 787
rect 44767 753 44935 787
rect 44935 753 44936 787
rect 44766 752 44936 753
rect 45138 895 45308 896
rect 45138 861 45139 895
rect 45139 861 45307 895
rect 45307 861 45308 895
rect 45138 787 45308 861
rect 45138 753 45139 787
rect 45139 753 45307 787
rect 45307 753 45308 787
rect 45138 752 45308 753
rect 45510 895 45680 896
rect 45510 861 45511 895
rect 45511 861 45679 895
rect 45679 861 45680 895
rect 45510 787 45680 861
rect 45510 753 45511 787
rect 45511 753 45679 787
rect 45679 753 45680 787
rect 45510 752 45680 753
rect 45882 895 46052 896
rect 45882 861 45883 895
rect 45883 861 46051 895
rect 46051 861 46052 895
rect 45882 787 46052 861
rect 45882 753 45883 787
rect 45883 753 46051 787
rect 46051 753 46052 787
rect 45882 752 46052 753
rect 46254 895 46424 896
rect 46254 861 46255 895
rect 46255 861 46423 895
rect 46423 861 46424 895
rect 46254 787 46424 861
rect 46254 753 46255 787
rect 46255 753 46423 787
rect 46423 753 46424 787
rect 46254 752 46424 753
rect 46626 895 46796 896
rect 46626 861 46627 895
rect 46627 861 46795 895
rect 46795 861 46796 895
rect 46626 787 46796 861
rect 46626 753 46627 787
rect 46627 753 46795 787
rect 46795 753 46796 787
rect 46626 752 46796 753
rect 46998 895 47168 896
rect 46998 861 46999 895
rect 46999 861 47167 895
rect 47167 861 47168 895
rect 46998 787 47168 861
rect 46998 753 46999 787
rect 46999 753 47167 787
rect 47167 753 47168 787
rect 46998 752 47168 753
rect 47370 895 47540 896
rect 47370 861 47371 895
rect 47371 861 47539 895
rect 47539 861 47540 895
rect 47370 787 47540 861
rect 47370 753 47371 787
rect 47371 753 47539 787
rect 47539 753 47540 787
rect 47370 752 47540 753
rect 47742 895 47912 896
rect 47742 861 47743 895
rect 47743 861 47911 895
rect 47911 861 47912 895
rect 47742 787 47912 861
rect 47742 753 47743 787
rect 47743 753 47911 787
rect 47911 753 47912 787
rect 47742 752 47912 753
rect 48114 895 48284 896
rect 48114 861 48115 895
rect 48115 861 48283 895
rect 48283 861 48284 895
rect 48114 787 48284 861
rect 48114 753 48115 787
rect 48115 753 48283 787
rect 48283 753 48284 787
rect 48114 752 48284 753
rect 39558 477 39728 488
rect 39558 443 39559 477
rect 39559 443 39727 477
rect 39727 443 39728 477
rect 39558 432 39728 443
rect 39930 477 40100 488
rect 39930 443 39931 477
rect 39931 443 40099 477
rect 40099 443 40100 477
rect 39930 432 40100 443
rect 40302 477 40472 488
rect 40302 443 40303 477
rect 40303 443 40471 477
rect 40471 443 40472 477
rect 40302 432 40472 443
rect 40674 477 40844 488
rect 40674 443 40675 477
rect 40675 443 40843 477
rect 40843 443 40844 477
rect 40674 432 40844 443
rect 41046 477 41216 488
rect 41046 443 41047 477
rect 41047 443 41215 477
rect 41215 443 41216 477
rect 41046 432 41216 443
rect 41418 477 41588 488
rect 41418 443 41419 477
rect 41419 443 41587 477
rect 41587 443 41588 477
rect 41418 432 41588 443
rect 41790 477 41960 488
rect 41790 443 41791 477
rect 41791 443 41959 477
rect 41959 443 41960 477
rect 41790 432 41960 443
rect 42162 477 42332 488
rect 42162 443 42163 477
rect 42163 443 42331 477
rect 42331 443 42332 477
rect 42162 432 42332 443
rect 42534 477 42704 488
rect 42534 443 42535 477
rect 42535 443 42703 477
rect 42703 443 42704 477
rect 42534 432 42704 443
rect 42906 477 43076 488
rect 42906 443 42907 477
rect 42907 443 43075 477
rect 43075 443 43076 477
rect 42906 432 43076 443
rect 43278 477 43448 488
rect 43278 443 43279 477
rect 43279 443 43447 477
rect 43447 443 43448 477
rect 43278 432 43448 443
rect 43650 477 43820 488
rect 43650 443 43651 477
rect 43651 443 43819 477
rect 43819 443 43820 477
rect 43650 432 43820 443
rect 44022 477 44192 488
rect 44022 443 44023 477
rect 44023 443 44191 477
rect 44191 443 44192 477
rect 44022 432 44192 443
rect 44394 477 44564 488
rect 44394 443 44395 477
rect 44395 443 44563 477
rect 44563 443 44564 477
rect 44394 432 44564 443
rect 44766 477 44936 488
rect 44766 443 44767 477
rect 44767 443 44935 477
rect 44935 443 44936 477
rect 44766 432 44936 443
rect 45138 477 45308 488
rect 45138 443 45139 477
rect 45139 443 45307 477
rect 45307 443 45308 477
rect 45138 432 45308 443
rect 45510 477 45680 488
rect 45510 443 45511 477
rect 45511 443 45679 477
rect 45679 443 45680 477
rect 45510 432 45680 443
rect 45882 477 46052 488
rect 45882 443 45883 477
rect 45883 443 46051 477
rect 46051 443 46052 477
rect 45882 432 46052 443
rect 46254 477 46424 488
rect 46254 443 46255 477
rect 46255 443 46423 477
rect 46423 443 46424 477
rect 46254 432 46424 443
rect 46626 477 46796 488
rect 46626 443 46627 477
rect 46627 443 46795 477
rect 46795 443 46796 477
rect 46626 432 46796 443
rect 46998 477 47168 488
rect 46998 443 46999 477
rect 46999 443 47167 477
rect 47167 443 47168 477
rect 46998 432 47168 443
rect 47370 477 47540 488
rect 47370 443 47371 477
rect 47371 443 47539 477
rect 47539 443 47540 477
rect 47370 432 47540 443
rect 47742 477 47912 488
rect 47742 443 47743 477
rect 47743 443 47911 477
rect 47911 443 47912 477
rect 47742 432 47912 443
rect 48114 477 48284 488
rect 48114 443 48115 477
rect 48115 443 48283 477
rect 48283 443 48284 477
rect 48114 432 48284 443
rect 39378 78 39578 278
rect 40102 78 40302 278
rect 40846 78 41046 278
rect 41590 78 41790 278
rect 42334 78 42534 278
rect 43078 78 43278 278
rect 43822 78 44022 278
rect 44566 78 44766 278
rect 45310 78 45510 278
rect 46054 78 46254 278
rect 46798 78 46998 278
rect 47542 78 47742 278
rect 48286 78 48486 278
<< metal2 >>
rect 35528 11896 36446 11906
rect 35528 10918 36446 10928
rect 38240 9524 38440 9534
rect 38240 9314 38440 9324
rect 38984 9524 39184 9534
rect 38984 9314 39184 9324
rect 39728 9524 39928 9534
rect 39728 9314 39928 9324
rect 40472 9524 40672 9534
rect 40472 9314 40672 9324
rect 41216 9524 41416 9534
rect 41216 9314 41416 9324
rect 41960 9524 42160 9534
rect 41960 9314 42160 9324
rect 42704 9524 42904 9534
rect 42704 9314 42904 9324
rect 43448 9524 43648 9534
rect 43448 9314 43648 9324
rect 43820 9524 44020 9534
rect 43820 9314 44020 9324
rect 44564 9524 44764 9534
rect 44564 9314 44764 9324
rect 45308 9524 45508 9534
rect 45308 9314 45508 9324
rect 46052 9524 46252 9534
rect 46052 9314 46252 9324
rect 46796 9524 46996 9534
rect 46796 9314 46996 9324
rect 47540 9524 47740 9534
rect 47540 9314 47740 9324
rect 48284 9524 48484 9534
rect 48284 9314 48484 9324
rect 49028 9524 49228 9534
rect 49028 9314 49228 9324
rect 49772 9524 49972 9534
rect 49772 9314 49972 9324
rect 38070 9136 49782 9146
rect 38240 9076 38442 9136
rect 38612 9076 38814 9136
rect 38984 9076 39186 9136
rect 39356 9076 39558 9136
rect 39728 9076 39930 9136
rect 40100 9076 40302 9136
rect 40472 9076 40674 9136
rect 40844 9076 41046 9136
rect 41216 9076 41418 9136
rect 41588 9076 41790 9136
rect 41960 9076 42162 9136
rect 42332 9076 42534 9136
rect 42704 9076 42906 9136
rect 43076 9076 43278 9136
rect 43448 9076 43650 9136
rect 43820 9076 44022 9136
rect 44192 9076 44394 9136
rect 44564 9076 44766 9136
rect 44936 9076 45138 9136
rect 45308 9076 45510 9136
rect 45680 9076 45882 9136
rect 46052 9076 46254 9136
rect 46424 9076 46626 9136
rect 46796 9076 46998 9136
rect 47168 9076 47370 9136
rect 47540 9076 47742 9136
rect 47912 9076 48114 9136
rect 48284 9076 48486 9136
rect 48656 9076 48858 9136
rect 49028 9076 49230 9136
rect 49400 9076 49602 9136
rect 49772 9076 49782 9136
rect 38070 9066 49782 9076
rect 38070 8596 49772 8606
rect 38240 8452 38442 8596
rect 38612 8452 38814 8596
rect 38984 8452 39186 8596
rect 39356 8452 39558 8596
rect 39728 8452 39930 8596
rect 40100 8452 40302 8596
rect 40472 8452 40674 8596
rect 40844 8452 41046 8596
rect 41216 8452 41418 8596
rect 41588 8452 41790 8596
rect 41960 8452 42162 8596
rect 42332 8452 42534 8596
rect 42704 8452 42906 8596
rect 43076 8452 43278 8596
rect 43448 8452 43650 8596
rect 43820 8452 44022 8596
rect 44192 8452 44394 8596
rect 44564 8452 44766 8596
rect 44936 8452 45138 8596
rect 45308 8452 45510 8596
rect 45680 8452 45882 8596
rect 46052 8452 46254 8596
rect 46424 8452 46626 8596
rect 46796 8452 46998 8596
rect 47168 8452 47370 8596
rect 47540 8452 47742 8596
rect 47912 8452 48114 8596
rect 48284 8452 48486 8596
rect 48656 8452 48858 8596
rect 49028 8452 49230 8596
rect 49400 8452 49602 8596
rect 38070 8442 49772 8452
rect 38070 7960 49772 7970
rect 38240 7816 38442 7960
rect 38612 7816 38814 7960
rect 38984 7816 39186 7960
rect 39356 7816 39558 7960
rect 39728 7816 39930 7960
rect 40100 7816 40302 7960
rect 40472 7816 40674 7960
rect 40844 7816 41046 7960
rect 41216 7816 41418 7960
rect 41588 7816 41790 7960
rect 41960 7816 42162 7960
rect 42332 7816 42534 7960
rect 42704 7816 42906 7960
rect 43076 7816 43278 7960
rect 43448 7816 43650 7960
rect 43820 7816 44022 7960
rect 44192 7816 44394 7960
rect 44564 7816 44766 7960
rect 44936 7816 45138 7960
rect 45308 7816 45510 7960
rect 45680 7816 45882 7960
rect 46052 7816 46254 7960
rect 46424 7816 46626 7960
rect 46796 7816 46998 7960
rect 47168 7816 47370 7960
rect 47540 7816 47742 7960
rect 47912 7816 48114 7960
rect 48284 7816 48486 7960
rect 48656 7816 48858 7960
rect 49028 7816 49230 7960
rect 49400 7816 49602 7960
rect 38070 7806 49772 7816
rect 38070 7336 49772 7346
rect 38240 7276 38442 7336
rect 38612 7276 38814 7336
rect 38984 7276 39186 7336
rect 39356 7276 39558 7336
rect 39728 7276 39930 7336
rect 40100 7276 40302 7336
rect 40472 7276 40674 7336
rect 40844 7276 41046 7336
rect 41216 7276 41418 7336
rect 41588 7276 41790 7336
rect 41960 7276 42162 7336
rect 42332 7276 42534 7336
rect 42704 7276 42906 7336
rect 43076 7276 43278 7336
rect 43448 7276 43650 7336
rect 43820 7276 44022 7336
rect 44192 7276 44394 7336
rect 44564 7276 44766 7336
rect 44936 7276 45138 7336
rect 45308 7276 45510 7336
rect 45680 7276 45882 7336
rect 46052 7276 46254 7336
rect 46424 7276 46626 7336
rect 46796 7276 46998 7336
rect 47168 7276 47370 7336
rect 47540 7276 47742 7336
rect 47912 7276 48114 7336
rect 48284 7276 48486 7336
rect 48656 7276 48858 7336
rect 49028 7276 49230 7336
rect 49400 7276 49602 7336
rect 38070 7266 49772 7276
rect 35702 7216 36308 7226
rect 44154 6968 49644 6978
rect 36308 6850 42146 6948
rect 39744 6760 39914 6850
rect 41976 6760 42146 6850
rect 39558 6750 40100 6760
rect 39728 6686 39930 6750
rect 39558 6676 40100 6686
rect 40302 6750 41588 6760
rect 40472 6686 40674 6750
rect 40844 6686 41046 6750
rect 41216 6686 41418 6750
rect 40302 6676 41588 6686
rect 41790 6750 42332 6760
rect 41960 6686 42162 6750
rect 44436 6696 44898 6968
rect 45180 6696 45642 6968
rect 45924 6696 46386 6968
rect 46668 6696 47130 6968
rect 47412 6696 47874 6968
rect 48156 6696 48618 6968
rect 48900 6696 49362 6968
rect 44154 6686 49644 6696
rect 41790 6676 42332 6686
rect 35702 6584 36308 6594
rect 39802 5818 39856 6676
rect 40546 5818 40600 6676
rect 41290 5818 41344 6676
rect 42034 5818 42088 6676
rect 39558 5808 40100 5818
rect 39728 5664 39930 5808
rect 39558 5654 40100 5664
rect 40302 5808 41588 5818
rect 40472 5664 40674 5808
rect 40844 5664 41046 5808
rect 41216 5664 41418 5808
rect 40302 5654 41588 5664
rect 41790 5808 42332 5818
rect 41960 5664 42162 5808
rect 41790 5654 42332 5664
rect 39802 4782 39856 5654
rect 40546 4782 40600 5654
rect 41290 4782 41344 5654
rect 42034 4782 42088 5654
rect 43036 5252 43318 5262
rect 43036 4970 43318 4980
rect 39558 4772 40100 4782
rect 39728 4628 39930 4772
rect 39558 4618 40100 4628
rect 40302 4772 41588 4782
rect 40472 4628 40674 4772
rect 40844 4628 41046 4772
rect 41216 4628 41418 4772
rect 40302 4618 41588 4628
rect 41790 4772 42332 4782
rect 41960 4628 42162 4772
rect 41790 4618 42332 4628
rect 43460 4712 43612 4722
rect 39802 3746 39856 4618
rect 40546 3746 40600 4618
rect 41290 3746 41344 4618
rect 42034 3746 42088 4618
rect 43460 4538 43612 4548
rect 43460 4312 43612 4322
rect 43460 4138 43612 4148
rect 43460 3912 43612 3922
rect 39558 3736 40100 3746
rect 39728 3592 39930 3736
rect 39558 3582 40100 3592
rect 40302 3736 41588 3746
rect 40472 3592 40674 3736
rect 40844 3592 41046 3736
rect 41216 3592 41418 3736
rect 40302 3582 41588 3592
rect 41790 3736 42332 3746
rect 43460 3738 43612 3748
rect 41960 3592 42162 3736
rect 41790 3582 42332 3592
rect 39802 2720 39856 3582
rect 40546 2720 40600 3582
rect 41290 2720 41344 3582
rect 42034 2720 42088 3582
rect 43460 3512 43612 3522
rect 43460 3338 43612 3348
rect 42664 2786 48164 2796
rect 39558 2710 40100 2720
rect 39728 2656 39930 2710
rect 39558 2646 40100 2656
rect 40302 2710 41588 2720
rect 40472 2656 40674 2710
rect 40844 2656 41046 2710
rect 41216 2656 41418 2710
rect 40302 2646 41588 2656
rect 41790 2710 42332 2720
rect 41960 2656 42162 2710
rect 41790 2646 42332 2656
rect 40488 2546 40658 2646
rect 41232 2546 41402 2646
rect 38802 2448 41402 2546
rect 42946 2622 43408 2786
rect 42664 2504 42946 2514
rect 43690 2622 44152 2786
rect 43408 2504 43690 2514
rect 44434 2622 44896 2786
rect 44152 2504 44434 2514
rect 45178 2622 45640 2786
rect 44896 2504 45178 2514
rect 45922 2622 46384 2786
rect 45640 2504 45922 2514
rect 46666 2622 47128 2786
rect 46384 2504 46666 2514
rect 47410 2622 47872 2786
rect 47128 2504 47410 2514
rect 48154 2622 48164 2786
rect 47872 2504 48154 2514
rect 43044 2440 43294 2450
rect 40538 2370 43044 2380
rect 41352 2236 43044 2370
rect 41352 2190 42518 2236
rect 40538 2180 42518 2190
rect 43044 2180 43294 2190
rect 42392 2062 42518 2180
rect 39558 2052 42344 2062
rect 39728 1996 39930 2052
rect 40100 1996 40302 2052
rect 40472 1996 40674 2052
rect 40844 1996 41046 2052
rect 41216 1996 41418 2052
rect 41588 1996 41790 2052
rect 41960 1996 42162 2052
rect 42332 1996 42344 2052
rect 39558 1986 42344 1996
rect 42392 2052 48284 2062
rect 42392 1996 42534 2052
rect 42704 1996 42906 2052
rect 43076 1996 43278 2052
rect 43448 1996 43650 2052
rect 43820 1996 44022 2052
rect 44192 1996 44394 2052
rect 44564 1996 44766 2052
rect 44936 1996 45138 2052
rect 45308 1996 45510 2052
rect 45680 1996 45882 2052
rect 46052 1996 46254 2052
rect 46424 1996 46626 2052
rect 46796 1996 46998 2052
rect 47168 1996 47370 2052
rect 47540 1996 47742 2052
rect 47912 1996 48114 2052
rect 42392 1986 48284 1996
rect 42392 1742 42518 1986
rect 39558 1732 42344 1742
rect 39728 1588 39930 1732
rect 40100 1588 40302 1732
rect 40472 1588 40674 1732
rect 40844 1588 41046 1732
rect 41216 1588 41418 1732
rect 41588 1588 41790 1732
rect 41960 1588 42162 1732
rect 42332 1588 42344 1732
rect 39558 1578 42344 1588
rect 42392 1732 48284 1742
rect 42392 1588 42534 1732
rect 42704 1588 42906 1732
rect 43076 1588 43278 1732
rect 43448 1588 43650 1732
rect 43820 1588 44022 1732
rect 44192 1588 44394 1732
rect 44564 1588 44766 1732
rect 44936 1588 45138 1732
rect 45308 1588 45510 1732
rect 45680 1588 45882 1732
rect 46052 1588 46254 1732
rect 46424 1588 46626 1732
rect 46796 1588 46998 1732
rect 47168 1588 47370 1732
rect 47540 1588 47742 1732
rect 47912 1588 48114 1732
rect 42392 1578 48284 1588
rect 42392 1324 42518 1578
rect 39558 1314 42344 1324
rect 39728 1170 39930 1314
rect 40100 1170 40302 1314
rect 40472 1170 40674 1314
rect 40844 1170 41046 1314
rect 41216 1170 41418 1314
rect 41588 1170 41790 1314
rect 41960 1170 42162 1314
rect 42332 1170 42344 1314
rect 39558 1160 42344 1170
rect 42392 1314 48284 1324
rect 42392 1170 42534 1314
rect 42704 1170 42906 1314
rect 43076 1170 43278 1314
rect 43448 1170 43650 1314
rect 43820 1170 44022 1314
rect 44192 1170 44394 1314
rect 44564 1170 44766 1314
rect 44936 1170 45138 1314
rect 45308 1170 45510 1314
rect 45680 1170 45882 1314
rect 46052 1170 46254 1314
rect 46424 1170 46626 1314
rect 46796 1170 46998 1314
rect 47168 1170 47370 1314
rect 47540 1170 47742 1314
rect 47912 1170 48114 1314
rect 42392 1160 48284 1170
rect 42392 906 42518 1160
rect 39558 896 42344 906
rect 39728 752 39930 896
rect 40100 752 40302 896
rect 40472 752 40674 896
rect 40844 752 41046 896
rect 41216 752 41418 896
rect 41588 752 41790 896
rect 41960 752 42162 896
rect 42332 752 42344 896
rect 39558 742 42344 752
rect 42392 896 48284 906
rect 42392 752 42534 896
rect 42704 752 42906 896
rect 43076 752 43278 896
rect 43448 752 43650 896
rect 43820 752 44022 896
rect 44192 752 44394 896
rect 44564 752 44766 896
rect 44936 752 45138 896
rect 45308 752 45510 896
rect 45680 752 45882 896
rect 46052 752 46254 896
rect 46424 752 46626 896
rect 46796 752 46998 896
rect 47168 752 47370 896
rect 47540 752 47742 896
rect 47912 752 48114 896
rect 42392 742 48284 752
rect 42392 498 42518 742
rect 39558 488 42344 498
rect 39728 432 39930 488
rect 40100 432 40302 488
rect 40472 432 40674 488
rect 40844 432 41046 488
rect 41216 432 41418 488
rect 41588 432 41790 488
rect 41960 432 42162 488
rect 42332 432 42344 488
rect 39558 422 42344 432
rect 42392 488 48284 498
rect 42392 432 42534 488
rect 42704 432 42906 488
rect 43076 432 43278 488
rect 43448 432 43650 488
rect 43820 432 44022 488
rect 44192 432 44394 488
rect 44564 432 44766 488
rect 44936 432 45138 488
rect 45308 432 45510 488
rect 45680 432 45882 488
rect 46052 432 46254 488
rect 46424 432 46626 488
rect 46796 432 46998 488
rect 47168 432 47370 488
rect 47540 432 47742 488
rect 47912 432 48114 488
rect 42392 422 48284 432
rect 39378 278 39578 288
rect 39378 68 39578 78
rect 40102 278 40302 288
rect 40102 68 40302 78
rect 40846 278 41046 288
rect 40846 68 41046 78
rect 41590 278 41790 288
rect 41590 68 41790 78
rect 42334 278 42534 288
rect 42334 68 42534 78
rect 43078 278 43278 288
rect 43078 68 43278 78
rect 43822 278 44022 288
rect 43822 68 44022 78
rect 44566 278 44766 288
rect 44566 68 44766 78
rect 45310 278 45510 288
rect 45310 68 45510 78
rect 46054 278 46254 288
rect 46054 68 46254 78
rect 46798 278 46998 288
rect 46798 68 46998 78
rect 47542 278 47742 288
rect 47542 68 47742 78
rect 48286 278 48486 288
rect 48286 68 48486 78
<< via2 >>
rect 35528 10928 36446 11896
rect 38240 9324 38440 9524
rect 38984 9324 39184 9524
rect 39728 9324 39928 9524
rect 40472 9324 40672 9524
rect 41216 9324 41416 9524
rect 41960 9324 42160 9524
rect 42704 9324 42904 9524
rect 43448 9324 43648 9524
rect 43820 9324 44020 9524
rect 44564 9324 44764 9524
rect 45308 9324 45508 9524
rect 46052 9324 46252 9524
rect 46796 9324 46996 9524
rect 47540 9324 47740 9524
rect 48284 9324 48484 9524
rect 49028 9324 49228 9524
rect 49772 9324 49972 9524
rect 45642 6696 45924 6968
rect 46386 6696 46668 6968
rect 47130 6696 47412 6968
rect 47874 6696 48156 6968
rect 43036 4980 43318 5252
rect 43460 4548 43612 4712
rect 43460 4148 43612 4312
rect 43460 3748 43612 3912
rect 43460 3348 43612 3512
rect 45640 2514 45922 2786
rect 46384 2514 46666 2786
rect 47128 2514 47410 2786
rect 47872 2514 48154 2786
rect 39378 78 39578 278
rect 40102 78 40302 278
rect 40846 78 41046 278
rect 41590 78 41790 278
rect 42334 78 42534 278
rect 43078 78 43278 278
rect 43822 78 44022 278
rect 44566 78 44766 278
rect 45310 78 45510 278
rect 46054 78 46254 278
rect 46798 78 46998 278
rect 47542 78 47742 278
rect 48286 78 48486 278
<< metal3 >>
rect 35518 11896 36456 11901
rect 35518 10928 35528 11896
rect 36446 10928 36456 11896
rect 35518 10923 36456 10928
rect 36804 10882 51914 25982
rect 38230 9524 38450 9529
rect 38230 9324 38240 9524
rect 38440 9324 38450 9524
rect 38230 9319 38450 9324
rect 38974 9524 39194 9529
rect 38974 9324 38984 9524
rect 39184 9324 39194 9524
rect 38974 9319 39194 9324
rect 39718 9524 39938 9529
rect 39718 9324 39728 9524
rect 39928 9324 39938 9524
rect 39718 9319 39938 9324
rect 40462 9524 40682 9529
rect 40462 9324 40472 9524
rect 40672 9324 40682 9524
rect 40462 9319 40682 9324
rect 41206 9524 41426 9529
rect 41206 9324 41216 9524
rect 41416 9324 41426 9524
rect 41206 9319 41426 9324
rect 41950 9524 42170 9529
rect 41950 9324 41960 9524
rect 42160 9324 42170 9524
rect 41950 9319 42170 9324
rect 42694 9524 42914 9529
rect 42694 9324 42704 9524
rect 42904 9324 42914 9524
rect 42694 9319 42914 9324
rect 43438 9524 43658 9529
rect 43438 9324 43448 9524
rect 43648 9324 43658 9524
rect 43438 9319 43658 9324
rect 43810 9524 44030 9529
rect 43810 9324 43820 9524
rect 44020 9324 44030 9524
rect 43810 9319 44030 9324
rect 44554 9524 44774 9529
rect 44554 9324 44564 9524
rect 44764 9324 44774 9524
rect 44554 9319 44774 9324
rect 45298 9524 45518 9529
rect 45298 9324 45308 9524
rect 45508 9324 45518 9524
rect 45298 9319 45518 9324
rect 46042 9524 46262 9529
rect 46042 9324 46052 9524
rect 46252 9324 46262 9524
rect 46042 9319 46262 9324
rect 46786 9524 47006 9529
rect 46786 9324 46796 9524
rect 46996 9324 47006 9524
rect 46786 9319 47006 9324
rect 47530 9524 47750 9529
rect 47530 9324 47540 9524
rect 47740 9324 47750 9524
rect 47530 9319 47750 9324
rect 48274 9524 48494 9529
rect 48274 9324 48284 9524
rect 48484 9324 48494 9524
rect 48274 9319 48494 9324
rect 49018 9524 49238 9529
rect 49018 9324 49028 9524
rect 49228 9324 49238 9524
rect 49018 9319 49238 9324
rect 49762 9524 49982 9529
rect 49762 9324 49772 9524
rect 49972 9324 49982 9524
rect 49762 9319 49982 9324
rect 50586 7002 50942 10882
rect 45632 6968 45934 6973
rect 45632 6696 45642 6968
rect 45924 6696 45934 6968
rect 45632 6490 45934 6696
rect 46376 6968 46678 6973
rect 46376 6696 46386 6968
rect 46668 6696 46678 6968
rect 46376 6490 46678 6696
rect 47120 6968 47422 6973
rect 47120 6696 47130 6968
rect 47412 6696 47422 6968
rect 47120 6490 47422 6696
rect 47864 6968 48166 6973
rect 47864 6696 47874 6968
rect 48156 6696 48166 6968
rect 47864 6490 48166 6696
rect 50032 6490 53008 7002
rect 43026 5252 43328 5257
rect 43026 4980 43036 5252
rect 43318 4980 43328 5252
rect 43026 4975 43328 4980
rect 43450 4712 43622 4717
rect 43450 4548 43460 4712
rect 43612 4548 43622 4712
rect 43450 4543 43622 4548
rect 43802 4514 53008 6490
rect 43450 4312 43622 4317
rect 43450 4148 43460 4312
rect 43612 4148 43622 4312
rect 43450 4143 43622 4148
rect 43802 4028 53482 4514
rect 43450 3912 43622 3917
rect 43450 3748 43460 3912
rect 43612 3748 43622 3912
rect 43450 3743 43622 3748
rect 43450 3512 43622 3517
rect 43450 3348 43460 3512
rect 43612 3348 43622 3512
rect 43802 3490 53008 4028
rect 43450 3343 43622 3348
rect 45630 2786 45932 3490
rect 45630 2514 45640 2786
rect 45922 2514 45932 2786
rect 45630 2509 45932 2514
rect 46374 2786 46676 3490
rect 46374 2514 46384 2786
rect 46666 2514 46676 2786
rect 46374 2509 46676 2514
rect 47118 2786 47420 3490
rect 47118 2514 47128 2786
rect 47410 2514 47420 2786
rect 47118 2509 47420 2514
rect 47862 2786 48164 3490
rect 47862 2514 47872 2786
rect 48154 2514 48164 2786
rect 47862 2509 48164 2514
rect 50032 802 53008 3490
rect 39368 278 39588 283
rect 39368 78 39378 278
rect 39578 78 39588 278
rect 39368 73 39588 78
rect 40092 278 40312 283
rect 40092 78 40102 278
rect 40302 78 40312 278
rect 40092 73 40312 78
rect 40836 278 41056 283
rect 40836 78 40846 278
rect 41046 78 41056 278
rect 40836 73 41056 78
rect 41580 278 41800 283
rect 41580 78 41590 278
rect 41790 78 41800 278
rect 41580 73 41800 78
rect 42324 278 42544 283
rect 42324 78 42334 278
rect 42534 78 42544 278
rect 42324 73 42544 78
rect 43068 278 43288 283
rect 43068 78 43078 278
rect 43278 78 43288 278
rect 43068 73 43288 78
rect 43812 278 44032 283
rect 43812 78 43822 278
rect 44022 78 44032 278
rect 43812 73 44032 78
rect 44556 278 44776 283
rect 44556 78 44566 278
rect 44766 78 44776 278
rect 44556 73 44776 78
rect 45300 278 45520 283
rect 45300 78 45310 278
rect 45510 78 45520 278
rect 45300 73 45520 78
rect 46044 278 46264 283
rect 46044 78 46054 278
rect 46254 78 46264 278
rect 46044 73 46264 78
rect 46788 278 47008 283
rect 46788 78 46798 278
rect 46998 78 47008 278
rect 46788 73 47008 78
rect 47532 278 47752 283
rect 47532 78 47542 278
rect 47742 78 47752 278
rect 47532 73 47752 78
rect 48276 278 48496 283
rect 48276 78 48286 278
rect 48486 78 48496 278
rect 48276 73 48496 78
<< via3 >>
rect 35528 10928 36446 11896
rect 38240 9324 38440 9524
rect 38984 9324 39184 9524
rect 39728 9324 39928 9524
rect 40472 9324 40672 9524
rect 41216 9324 41416 9524
rect 41960 9324 42160 9524
rect 42704 9324 42904 9524
rect 43448 9324 43648 9524
rect 43820 9324 44020 9524
rect 44564 9324 44764 9524
rect 45308 9324 45508 9524
rect 46052 9324 46252 9524
rect 46796 9324 46996 9524
rect 47540 9324 47740 9524
rect 48284 9324 48484 9524
rect 49028 9324 49228 9524
rect 49772 9324 49972 9524
rect 43036 4980 43318 5252
rect 43460 4548 43612 4712
rect 43460 4148 43612 4312
rect 43460 3748 43612 3912
rect 43460 3348 43612 3512
rect 39378 78 39578 278
rect 40102 78 40302 278
rect 40846 78 41046 278
rect 41590 78 41790 278
rect 42334 78 42534 278
rect 43078 78 43278 278
rect 43822 78 44022 278
rect 44566 78 44766 278
rect 45310 78 45510 278
rect 46054 78 46254 278
rect 46798 78 46998 278
rect 47542 78 47742 278
rect 48286 78 48486 278
<< mimcap >>
rect 36905 25842 40405 25882
rect 36905 22422 36945 25842
rect 40365 22422 40405 25842
rect 36905 22382 40405 22422
rect 40724 25842 44224 25882
rect 40724 22422 40764 25842
rect 44184 22422 44224 25842
rect 40724 22382 44224 22422
rect 44543 25842 48043 25882
rect 44543 22422 44583 25842
rect 48003 22422 48043 25842
rect 44543 22382 48043 22422
rect 48362 25842 51862 25882
rect 48362 22422 48402 25842
rect 51822 22422 51862 25842
rect 48362 22382 51862 22422
rect 36905 22042 40405 22082
rect 36905 18622 36945 22042
rect 40365 18622 40405 22042
rect 36905 18582 40405 18622
rect 40724 22042 44224 22082
rect 40724 18622 40764 22042
rect 44184 18622 44224 22042
rect 40724 18582 44224 18622
rect 44543 22042 48043 22082
rect 44543 18622 44583 22042
rect 48003 18622 48043 22042
rect 44543 18582 48043 18622
rect 48362 22042 51862 22082
rect 48362 18622 48402 22042
rect 51822 18622 51862 22042
rect 48362 18582 51862 18622
rect 36905 18242 40405 18282
rect 36905 14822 36945 18242
rect 40365 14822 40405 18242
rect 36905 14782 40405 14822
rect 40724 18242 44224 18282
rect 40724 14822 40764 18242
rect 44184 14822 44224 18242
rect 40724 14782 44224 14822
rect 44543 18242 48043 18282
rect 44543 14822 44583 18242
rect 48003 14822 48043 18242
rect 44543 14782 48043 14822
rect 48362 18242 51862 18282
rect 48362 14822 48402 18242
rect 51822 14822 51862 18242
rect 48362 14782 51862 14822
rect 36905 14442 40405 14482
rect 36905 11022 36945 14442
rect 40365 11022 40405 14442
rect 36905 10982 40405 11022
rect 40724 14442 44224 14482
rect 40724 11022 40764 14442
rect 44184 11022 44224 14442
rect 40724 10982 44224 11022
rect 44543 14442 48043 14482
rect 44543 11022 44583 14442
rect 48003 11022 48043 14442
rect 44543 10982 48043 11022
rect 48362 14442 51862 14482
rect 48362 11022 48402 14442
rect 51822 11022 51862 14442
rect 48362 10982 51862 11022
rect 50132 6862 52932 6902
rect 43902 6350 49902 6390
rect 43902 3630 43942 6350
rect 49862 3630 49902 6350
rect 43902 3590 49902 3630
rect 50132 942 50172 6862
rect 52892 942 52932 6862
rect 50132 902 52932 942
<< mimcapcontact >>
rect 36945 22422 40365 25842
rect 40764 22422 44184 25842
rect 44583 22422 48003 25842
rect 48402 22422 51822 25842
rect 36945 18622 40365 22042
rect 40764 18622 44184 22042
rect 44583 18622 48003 22042
rect 48402 18622 51822 22042
rect 36945 14822 40365 18242
rect 40764 14822 44184 18242
rect 44583 14822 48003 18242
rect 48402 14822 51822 18242
rect 36945 11022 40365 14442
rect 40764 11022 44184 14442
rect 44583 11022 48003 14442
rect 48402 11022 51822 14442
rect 43942 3630 49862 6350
rect 50172 942 52892 6862
<< metal4 >>
rect 38603 25982 38707 26032
rect 42422 25982 42526 26032
rect 46241 25982 46345 26032
rect 50060 25982 50164 26032
rect 36804 25842 51914 25982
rect 36804 22422 36945 25842
rect 40365 22422 40764 25842
rect 44184 22422 44583 25842
rect 48003 22422 48402 25842
rect 51822 22422 51914 25842
rect 36804 22042 51914 22422
rect 36804 18622 36945 22042
rect 40365 18622 40764 22042
rect 44184 18622 44583 22042
rect 48003 18622 48402 22042
rect 51822 18622 51914 22042
rect 36804 18242 51914 18622
rect 36804 14822 36945 18242
rect 40365 14822 40764 18242
rect 44184 14822 44583 18242
rect 48003 14822 48402 18242
rect 51822 14822 51914 18242
rect 36804 14442 51914 14822
rect 35527 11896 36447 11897
rect 35527 10928 35528 11896
rect 36446 11726 36447 11896
rect 36804 11726 36945 14442
rect 36446 11150 36945 11726
rect 36446 10928 36447 11150
rect 35527 10927 36447 10928
rect 36804 11022 36945 11150
rect 40365 11022 40764 14442
rect 44184 11022 44583 14442
rect 48003 11022 48402 14442
rect 51822 11022 51914 14442
rect 36804 10882 51914 11022
rect 38603 10832 38707 10882
rect 42422 10832 42526 10882
rect 46241 10832 46345 10882
rect 50060 10832 50164 10882
rect 37634 9524 50158 10302
rect 37634 9324 38240 9524
rect 38440 9324 38984 9524
rect 39184 9324 39728 9524
rect 39928 9324 40472 9524
rect 40672 9324 41216 9524
rect 41416 9324 41960 9524
rect 42160 9324 42704 9524
rect 42904 9324 43448 9524
rect 43648 9324 43820 9524
rect 44020 9324 44564 9524
rect 44764 9324 45308 9524
rect 45508 9324 46052 9524
rect 46252 9324 46796 9524
rect 46996 9324 47540 9524
rect 47740 9324 48284 9524
rect 48484 9324 49028 9524
rect 49228 9324 49772 9524
rect 49972 9324 50158 9524
rect 37634 9298 50158 9324
rect 50171 6862 52893 6863
rect 50171 6352 50172 6862
rect 49816 6351 50172 6352
rect 43941 6350 50172 6351
rect 43035 5252 43319 5253
rect 43035 4980 43036 5252
rect 43318 5224 43319 5252
rect 43941 5224 43942 6350
rect 43318 5006 43942 5224
rect 43318 4980 43319 5006
rect 43035 4979 43319 4980
rect 43426 4712 43636 4810
rect 43426 4548 43460 4712
rect 43612 4548 43636 4712
rect 43426 4312 43636 4548
rect 43426 4148 43460 4312
rect 43612 4148 43636 4312
rect 43426 3912 43636 4148
rect 43426 3748 43460 3912
rect 43612 3748 43636 3912
rect 43426 3512 43636 3748
rect 43941 3630 43942 5006
rect 49862 3630 50172 6350
rect 43941 3629 50172 3630
rect 49816 3628 50172 3629
rect 43426 3348 43460 3512
rect 43612 3348 43636 3512
rect 43426 302 43636 3348
rect 50171 942 50172 3628
rect 52892 942 52893 6862
rect 50171 941 52893 942
rect 37634 278 50158 302
rect 37634 78 39378 278
rect 39578 78 40102 278
rect 40302 78 40846 278
rect 41046 78 41590 278
rect 41790 78 42334 278
rect 42534 78 43078 278
rect 43278 78 43822 278
rect 44022 78 44566 278
rect 44766 78 45310 278
rect 45510 78 46054 278
rect 46254 78 46798 278
rect 46998 78 47542 278
rect 47742 78 48286 278
rect 48486 78 50158 278
rect 37634 -702 50158 78
<< labels >>
flabel metal4 39558 9792 39558 9792 0 FreeSans 1600 0 0 0 vdd
port 0 nsew
flabel metal4 38326 -452 38326 -452 0 FreeSans 1600 0 0 0 vss
port 4 nsew
flabel metal2 36670 6904 36670 6904 0 FreeSans 1600 0 0 0 vi
port 1 nsew
flabel metal1 38030 7876 38030 7876 0 FreeSans 1600 0 0 0 vbias
port 2 nsew
flabel metal3 53248 4194 53248 4194 0 FreeSans 1600 0 0 0 vout
port 5 nsew
flabel metal2 38884 2478 38884 2478 0 FreeSans 1600 0 0 0 vref
port 3 nsew
<< end >>
