magic
tech sky130A
timestamp 1632370638
<< nwell >>
rect 48349 -3336 63487 11802
rect 48349 -21336 63487 -6198
rect 48349 -39336 63487 -24198
rect 48349 -57341 63487 -42203
<< pwell >>
rect 48280 11802 63556 11871
rect 48280 -3336 48349 11802
rect 63487 -3336 63556 11802
rect 48280 -3405 63556 -3336
rect 48280 -6198 63556 -6129
rect 48280 -21336 48349 -6198
rect 63487 -21336 63556 -6198
rect 48280 -21405 63556 -21336
rect 48280 -24198 63556 -24129
rect 48280 -39336 48349 -24198
rect 63487 -39336 63556 -24198
rect 48280 -39405 63556 -39336
rect 48280 -42203 63556 -42134
rect 48280 -57341 48349 -42203
rect 63487 -57341 63556 -42203
rect 48280 -57410 63556 -57341
<< psubdiff >>
rect 48298 11836 48346 11853
rect 63490 11836 63538 11853
rect 48298 11805 48315 11836
rect 63521 11805 63538 11836
rect 48298 -3370 48315 -3339
rect 63521 -3370 63538 -3339
rect 48298 -3387 48346 -3370
rect 63490 -3387 63538 -3370
rect 48298 -6164 48346 -6147
rect 63490 -6164 63538 -6147
rect 48298 -6195 48315 -6164
rect 63521 -6195 63538 -6164
rect 48298 -21370 48315 -21339
rect 63521 -21370 63538 -21339
rect 48298 -21387 48346 -21370
rect 63490 -21387 63538 -21370
rect 48298 -24164 48346 -24147
rect 63490 -24164 63538 -24147
rect 48298 -24195 48315 -24164
rect 63521 -24195 63538 -24164
rect 48298 -39370 48315 -39339
rect 63521 -39370 63538 -39339
rect 48298 -39387 48346 -39370
rect 63490 -39387 63538 -39370
rect 48298 -42169 48346 -42152
rect 63490 -42169 63538 -42152
rect 48298 -42200 48315 -42169
rect 63521 -42200 63538 -42169
rect 48298 -57375 48315 -57344
rect 63521 -57375 63538 -57344
rect 48298 -57392 48346 -57375
rect 63490 -57392 63538 -57375
<< nsubdiff >>
rect 48367 11767 48415 11784
rect 63421 11767 63469 11784
rect 48367 11736 48384 11767
rect 63452 11736 63469 11767
rect 48367 -3301 48384 -3270
rect 63452 -3301 63469 -3270
rect 48367 -3318 48415 -3301
rect 63421 -3318 63469 -3301
rect 48367 -6233 48415 -6216
rect 63421 -6233 63469 -6216
rect 48367 -6264 48384 -6233
rect 63452 -6264 63469 -6233
rect 48367 -21301 48384 -21270
rect 63452 -21301 63469 -21270
rect 48367 -21318 48415 -21301
rect 63421 -21318 63469 -21301
rect 48367 -24233 48415 -24216
rect 63421 -24233 63469 -24216
rect 48367 -24264 48384 -24233
rect 63452 -24264 63469 -24233
rect 48367 -39301 48384 -39270
rect 63452 -39301 63469 -39270
rect 48367 -39318 48415 -39301
rect 63421 -39318 63469 -39301
rect 48367 -42238 48415 -42221
rect 63421 -42238 63469 -42221
rect 48367 -42269 48384 -42238
rect 63452 -42269 63469 -42238
rect 48367 -57306 48384 -57275
rect 63452 -57306 63469 -57275
rect 48367 -57323 48415 -57306
rect 63421 -57323 63469 -57306
<< psubdiffcont >>
rect 48346 11836 63490 11853
rect 48298 -3339 48315 11805
rect 63521 -3339 63538 11805
rect 48346 -3387 63490 -3370
rect 48346 -6164 63490 -6147
rect 48298 -21339 48315 -6195
rect 63521 -21339 63538 -6195
rect 48346 -21387 63490 -21370
rect 48346 -24164 63490 -24147
rect 48298 -39339 48315 -24195
rect 63521 -39339 63538 -24195
rect 48346 -39387 63490 -39370
rect 48346 -42169 63490 -42152
rect 48298 -57344 48315 -42200
rect 63521 -57344 63538 -42200
rect 48346 -57392 63490 -57375
<< nsubdiffcont >>
rect 48415 11767 63421 11784
rect 48367 -3270 48384 11736
rect 63452 -3270 63469 11736
rect 48415 -3318 63421 -3301
rect 48415 -6233 63421 -6216
rect 48367 -21270 48384 -6264
rect 63452 -21270 63469 -6264
rect 48415 -21318 63421 -21301
rect 48415 -24233 63421 -24216
rect 48367 -39270 48384 -24264
rect 63452 -39270 63469 -24264
rect 48415 -39318 63421 -39301
rect 48415 -42238 63421 -42221
rect 48367 -57275 48384 -42269
rect 63452 -57275 63469 -42269
rect 48415 -57323 63421 -57306
<< pdiode >>
rect 48418 11727 63418 11733
rect 48418 -3261 48424 11727
rect 63412 -3261 63418 11727
rect 48418 -3267 63418 -3261
rect 48418 -6273 63418 -6267
rect 48418 -21261 48424 -6273
rect 63412 -21261 63418 -6273
rect 48418 -21267 63418 -21261
rect 48418 -24273 63418 -24267
rect 48418 -39261 48424 -24273
rect 63412 -39261 63418 -24273
rect 48418 -39267 63418 -39261
rect 48418 -42278 63418 -42272
rect 48418 -57266 48424 -42278
rect 63412 -57266 63418 -42278
rect 48418 -57272 63418 -57266
<< pdiodec >>
rect 48424 -3261 63412 11727
rect 48424 -21261 63412 -6273
rect 48424 -39261 63412 -24273
rect 48424 -57266 63412 -42278
<< locali >>
rect 48298 11836 48346 11853
rect 63490 11836 63538 11853
rect 48298 11805 48315 11836
rect 63521 11805 63538 11836
rect 48367 11767 48415 11784
rect 63421 11767 63469 11784
rect 48367 11736 48384 11767
rect 63452 11736 63469 11767
rect 48416 -3261 48424 11727
rect 63412 -3261 63420 11727
rect 48367 -3301 48384 -3270
rect 63452 -3301 63469 -3270
rect 48367 -3318 48410 -3301
rect 63425 -3318 63469 -3301
rect 48298 -3370 48315 -3339
rect 63521 -3370 63538 -3339
rect 48298 -3387 48346 -3370
rect 63490 -3387 63538 -3370
rect 48298 -6164 48346 -6147
rect 63490 -6164 63538 -6147
rect 48298 -6195 48315 -6164
rect 63521 -6195 63538 -6164
rect 48367 -6233 48415 -6216
rect 63421 -6233 63469 -6216
rect 48367 -6264 48384 -6233
rect 63452 -6264 63469 -6233
rect 48416 -21261 48424 -6273
rect 63412 -21261 63420 -6273
rect 48367 -21301 48384 -21270
rect 63452 -21301 63469 -21270
rect 48367 -21318 48415 -21301
rect 63430 -21318 63469 -21301
rect 48298 -21370 48315 -21339
rect 63521 -21370 63538 -21339
rect 48298 -21387 48346 -21370
rect 63490 -21387 63538 -21370
rect 48298 -24164 48346 -24147
rect 63490 -24164 63538 -24147
rect 48298 -24195 48315 -24164
rect 63521 -24195 63538 -24164
rect 48367 -24233 48415 -24216
rect 63421 -24233 63469 -24216
rect 48367 -24264 48384 -24233
rect 63452 -24264 63469 -24233
rect 48416 -39261 48424 -24273
rect 63412 -39261 63420 -24273
rect 48367 -39301 48384 -39270
rect 63452 -39301 63469 -39270
rect 48367 -39318 48415 -39301
rect 63425 -39318 63469 -39301
rect 48298 -39370 48315 -39339
rect 63521 -39370 63538 -39339
rect 48298 -39387 48346 -39370
rect 63490 -39387 63538 -39370
rect 48298 -42169 48346 -42152
rect 63490 -42169 63538 -42152
rect 48298 -42200 48315 -42169
rect 63521 -42200 63538 -42169
rect 48367 -42238 48415 -42221
rect 63421 -42238 63469 -42221
rect 48367 -42269 48384 -42238
rect 63452 -42269 63469 -42238
rect 48416 -57266 48424 -42278
rect 63412 -57266 63420 -42278
rect 48367 -57306 48384 -57275
rect 63452 -57305 63469 -57275
rect 48367 -57323 48410 -57306
rect 48298 -57375 48315 -57344
rect 63521 -57375 63538 -57344
rect 48298 -57392 48346 -57375
rect 63490 -57392 63538 -57375
<< viali >>
rect 48424 -3261 63412 11727
rect 48410 -3301 63425 -3295
rect 48410 -3318 48415 -3301
rect 48415 -3318 63421 -3301
rect 63421 -3318 63425 -3301
rect 48410 -3350 63425 -3318
rect 48424 -21261 63412 -6273
rect 48415 -21301 63430 -21295
rect 48415 -21318 63421 -21301
rect 63421 -21318 63430 -21301
rect 48415 -21350 63430 -21318
rect 48424 -39261 63412 -24273
rect 48415 -39301 63425 -39295
rect 48415 -39318 63421 -39301
rect 63421 -39318 63425 -39301
rect 48415 -39345 63425 -39318
rect 48424 -57266 63412 -42278
rect 48410 -57306 63490 -57305
rect 48410 -57323 48415 -57306
rect 48415 -57323 63421 -57306
rect 63421 -57323 63490 -57306
rect 48410 -57375 63490 -57323
rect 48410 -57392 63490 -57375
rect 48410 -57410 63490 -57392
<< metal1 >>
rect 48418 11727 63418 11730
rect 48418 -3261 48424 11727
rect 63412 -3261 63418 11727
rect 48418 -3264 63418 -3261
rect 48404 -3295 63431 -3292
rect 48404 -3350 48410 -3295
rect 63425 -3350 63431 -3295
rect 48404 -3353 63431 -3350
rect 48415 -6273 63425 -3353
rect 48415 -6275 48424 -6273
rect 48418 -21261 48424 -6275
rect 63412 -6275 63425 -6273
rect 63412 -21261 63418 -6275
rect 48418 -21264 63418 -21261
rect 48409 -21295 63436 -21292
rect 48409 -21350 48415 -21295
rect 63430 -21350 63436 -21295
rect 48409 -21353 63436 -21350
rect 48415 -24273 63430 -21353
rect 48415 -24275 48424 -24273
rect 48418 -39261 48424 -24275
rect 63412 -24275 63430 -24273
rect 63412 -39261 63418 -24275
rect 48418 -39264 63418 -39261
rect 48409 -39295 63431 -39292
rect 48409 -39345 48415 -39295
rect 63425 -39345 63431 -39295
rect 48409 -39348 63431 -39345
rect 48415 -42278 63425 -39348
rect 48415 -42280 48424 -42278
rect 48418 -57266 48424 -42280
rect 63412 -42280 63425 -42278
rect 63412 -57266 63418 -42280
rect 48418 -57269 63418 -57266
rect 48404 -57305 63496 -57302
rect 48404 -57410 48410 -57305
rect 63490 -57410 63496 -57305
rect 48404 -57413 63496 -57410
<< labels >>
flabel viali 56875 10630 56875 10630 0 FreeSans 16000 0 0 0 vdd
flabel viali 48595 -57365 48595 -57365 0 FreeSans 16000 0 0 0 vss
<< end >>
