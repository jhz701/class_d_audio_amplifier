magic
tech sky130A
magscale 1 2
timestamp 1625589597
<< nwell >>
rect -46 198 4911 1336
rect -46 174 4767 198
rect -46 165 530 174
<< nmos >>
rect 219 -510 249 -10
rect 315 -510 345 -10
rect 525 -510 555 -10
rect 621 -510 651 -10
rect 717 -510 747 -10
rect 813 -510 843 -10
rect 909 -510 939 -10
rect 1005 -510 1035 -10
rect 1101 -510 1131 -10
rect 1197 -510 1227 -10
rect 1423 -510 1453 -10
rect 1519 -510 1549 -10
rect 1615 -510 1645 -10
rect 1711 -510 1741 -10
rect 1807 -510 1837 -10
rect 1903 -510 1933 -10
rect 1999 -510 2029 -10
rect 2095 -510 2125 -10
rect 2191 -510 2221 -10
rect 2287 -510 2317 -10
rect 2383 -510 2413 -10
rect 2479 -510 2509 -10
rect 2575 -510 2605 -10
rect 2671 -510 2701 -10
rect 2767 -510 2797 -10
rect 2863 -510 2893 -10
rect 2959 -510 2989 -10
rect 3055 -510 3085 -10
rect 3151 -510 3181 -10
rect 3247 -510 3277 -10
rect 3343 -510 3373 -10
rect 3439 -510 3469 -10
rect 3535 -510 3565 -10
rect 3631 -510 3661 -10
rect 3727 -510 3757 -10
rect 3823 -510 3853 -10
rect 3919 -510 3949 -10
rect 4015 -510 4045 -10
rect 4111 -510 4141 -10
rect 4207 -510 4237 -10
rect 4303 -510 4333 -10
rect 4399 -510 4429 -10
rect 4495 -510 4525 -10
rect 4591 -510 4621 -10
rect 4687 -510 4717 -10
rect 4783 -510 4813 -10
<< pmos >>
rect 219 234 249 1234
rect 315 234 345 1234
rect 525 236 555 1236
rect 621 236 651 1236
rect 717 236 747 1236
rect 813 236 843 1236
rect 909 236 939 1236
rect 1005 236 1035 1236
rect 1101 236 1131 1236
rect 1197 236 1227 1236
rect 1423 236 1453 1236
rect 1519 236 1549 1236
rect 1615 236 1645 1236
rect 1711 236 1741 1236
rect 1807 236 1837 1236
rect 1903 236 1933 1236
rect 1999 236 2029 1236
rect 2095 236 2125 1236
rect 2191 236 2221 1236
rect 2287 236 2317 1236
rect 2383 236 2413 1236
rect 2479 236 2509 1236
rect 2575 236 2605 1236
rect 2671 236 2701 1236
rect 2767 236 2797 1236
rect 2863 236 2893 1236
rect 2959 236 2989 1236
rect 3055 236 3085 1236
rect 3151 236 3181 1236
rect 3247 236 3277 1236
rect 3343 236 3373 1236
rect 3439 236 3469 1236
rect 3535 236 3565 1236
rect 3631 236 3661 1236
rect 3727 236 3757 1236
rect 3823 236 3853 1236
rect 3919 236 3949 1236
rect 4015 236 4045 1236
rect 4111 236 4141 1236
rect 4207 236 4237 1236
rect 4303 236 4333 1236
rect 4399 236 4429 1236
rect 4495 236 4525 1236
rect 4591 236 4621 1236
rect 4687 236 4717 1236
rect 4783 236 4813 1236
<< ndiff >>
rect 157 -22 219 -10
rect 157 -498 169 -22
rect 203 -498 219 -22
rect 157 -510 219 -498
rect 249 -22 315 -10
rect 249 -498 265 -22
rect 299 -498 315 -22
rect 249 -510 315 -498
rect 345 -22 407 -10
rect 345 -498 361 -22
rect 395 -498 407 -22
rect 345 -510 407 -498
rect 463 -22 525 -10
rect 463 -498 475 -22
rect 509 -498 525 -22
rect 463 -510 525 -498
rect 555 -22 621 -10
rect 555 -498 571 -22
rect 605 -498 621 -22
rect 555 -510 621 -498
rect 651 -22 717 -10
rect 651 -498 667 -22
rect 701 -498 717 -22
rect 651 -510 717 -498
rect 747 -22 813 -10
rect 747 -498 763 -22
rect 797 -498 813 -22
rect 747 -510 813 -498
rect 843 -22 909 -10
rect 843 -498 859 -22
rect 893 -498 909 -22
rect 843 -510 909 -498
rect 939 -22 1005 -10
rect 939 -498 955 -22
rect 989 -498 1005 -22
rect 939 -510 1005 -498
rect 1035 -22 1101 -10
rect 1035 -498 1051 -22
rect 1085 -498 1101 -22
rect 1035 -510 1101 -498
rect 1131 -22 1197 -10
rect 1131 -498 1147 -22
rect 1181 -498 1197 -22
rect 1131 -510 1197 -498
rect 1227 -22 1289 -10
rect 1227 -498 1243 -22
rect 1277 -498 1289 -22
rect 1227 -510 1289 -498
rect 1361 -22 1423 -10
rect 1361 -498 1373 -22
rect 1407 -498 1423 -22
rect 1361 -510 1423 -498
rect 1453 -22 1519 -10
rect 1453 -498 1469 -22
rect 1503 -498 1519 -22
rect 1453 -510 1519 -498
rect 1549 -22 1615 -10
rect 1549 -498 1565 -22
rect 1599 -498 1615 -22
rect 1549 -510 1615 -498
rect 1645 -22 1711 -10
rect 1645 -498 1661 -22
rect 1695 -498 1711 -22
rect 1645 -510 1711 -498
rect 1741 -22 1807 -10
rect 1741 -498 1757 -22
rect 1791 -498 1807 -22
rect 1741 -510 1807 -498
rect 1837 -22 1903 -10
rect 1837 -498 1853 -22
rect 1887 -498 1903 -22
rect 1837 -510 1903 -498
rect 1933 -22 1999 -10
rect 1933 -498 1949 -22
rect 1983 -498 1999 -22
rect 1933 -510 1999 -498
rect 2029 -22 2095 -10
rect 2029 -498 2045 -22
rect 2079 -498 2095 -22
rect 2029 -510 2095 -498
rect 2125 -22 2191 -10
rect 2125 -498 2141 -22
rect 2175 -498 2191 -22
rect 2125 -510 2191 -498
rect 2221 -22 2287 -10
rect 2221 -498 2237 -22
rect 2271 -498 2287 -22
rect 2221 -510 2287 -498
rect 2317 -22 2383 -10
rect 2317 -498 2333 -22
rect 2367 -498 2383 -22
rect 2317 -510 2383 -498
rect 2413 -22 2479 -10
rect 2413 -498 2429 -22
rect 2463 -498 2479 -22
rect 2413 -510 2479 -498
rect 2509 -22 2575 -10
rect 2509 -498 2525 -22
rect 2559 -498 2575 -22
rect 2509 -510 2575 -498
rect 2605 -22 2671 -10
rect 2605 -498 2621 -22
rect 2655 -498 2671 -22
rect 2605 -510 2671 -498
rect 2701 -22 2767 -10
rect 2701 -498 2717 -22
rect 2751 -498 2767 -22
rect 2701 -510 2767 -498
rect 2797 -22 2863 -10
rect 2797 -498 2813 -22
rect 2847 -498 2863 -22
rect 2797 -510 2863 -498
rect 2893 -22 2959 -10
rect 2893 -498 2909 -22
rect 2943 -498 2959 -22
rect 2893 -510 2959 -498
rect 2989 -22 3055 -10
rect 2989 -498 3005 -22
rect 3039 -498 3055 -22
rect 2989 -510 3055 -498
rect 3085 -22 3151 -10
rect 3085 -498 3101 -22
rect 3135 -498 3151 -22
rect 3085 -510 3151 -498
rect 3181 -22 3247 -10
rect 3181 -498 3197 -22
rect 3231 -498 3247 -22
rect 3181 -510 3247 -498
rect 3277 -22 3343 -10
rect 3277 -498 3293 -22
rect 3327 -498 3343 -22
rect 3277 -510 3343 -498
rect 3373 -22 3439 -10
rect 3373 -498 3389 -22
rect 3423 -498 3439 -22
rect 3373 -510 3439 -498
rect 3469 -22 3535 -10
rect 3469 -498 3485 -22
rect 3519 -498 3535 -22
rect 3469 -510 3535 -498
rect 3565 -22 3631 -10
rect 3565 -498 3581 -22
rect 3615 -498 3631 -22
rect 3565 -510 3631 -498
rect 3661 -22 3727 -10
rect 3661 -498 3677 -22
rect 3711 -498 3727 -22
rect 3661 -510 3727 -498
rect 3757 -22 3823 -10
rect 3757 -498 3773 -22
rect 3807 -498 3823 -22
rect 3757 -510 3823 -498
rect 3853 -22 3919 -10
rect 3853 -498 3869 -22
rect 3903 -498 3919 -22
rect 3853 -510 3919 -498
rect 3949 -22 4015 -10
rect 3949 -498 3965 -22
rect 3999 -498 4015 -22
rect 3949 -510 4015 -498
rect 4045 -22 4111 -10
rect 4045 -498 4061 -22
rect 4095 -498 4111 -22
rect 4045 -510 4111 -498
rect 4141 -22 4207 -10
rect 4141 -498 4157 -22
rect 4191 -498 4207 -22
rect 4141 -510 4207 -498
rect 4237 -22 4303 -10
rect 4237 -498 4253 -22
rect 4287 -498 4303 -22
rect 4237 -510 4303 -498
rect 4333 -22 4399 -10
rect 4333 -498 4349 -22
rect 4383 -498 4399 -22
rect 4333 -510 4399 -498
rect 4429 -22 4495 -10
rect 4429 -498 4445 -22
rect 4479 -498 4495 -22
rect 4429 -510 4495 -498
rect 4525 -22 4591 -10
rect 4525 -498 4541 -22
rect 4575 -498 4591 -22
rect 4525 -510 4591 -498
rect 4621 -22 4687 -10
rect 4621 -498 4637 -22
rect 4671 -498 4687 -22
rect 4621 -510 4687 -498
rect 4717 -22 4783 -10
rect 4717 -498 4733 -22
rect 4767 -498 4783 -22
rect 4717 -510 4783 -498
rect 4813 -22 4875 -10
rect 4813 -498 4829 -22
rect 4863 -498 4875 -22
rect 4813 -510 4875 -498
<< pdiff >>
rect 157 1222 219 1234
rect 157 246 169 1222
rect 203 246 219 1222
rect 157 234 219 246
rect 249 1222 315 1234
rect 249 246 265 1222
rect 299 246 315 1222
rect 249 234 315 246
rect 345 1222 407 1234
rect 345 246 361 1222
rect 395 246 407 1222
rect 345 234 407 246
rect 463 1224 525 1236
rect 463 248 475 1224
rect 509 248 525 1224
rect 463 236 525 248
rect 555 1224 621 1236
rect 555 248 571 1224
rect 605 248 621 1224
rect 555 236 621 248
rect 651 1224 717 1236
rect 651 248 667 1224
rect 701 248 717 1224
rect 651 236 717 248
rect 747 1224 813 1236
rect 747 248 763 1224
rect 797 248 813 1224
rect 747 236 813 248
rect 843 1224 909 1236
rect 843 248 859 1224
rect 893 248 909 1224
rect 843 236 909 248
rect 939 1224 1005 1236
rect 939 248 955 1224
rect 989 248 1005 1224
rect 939 236 1005 248
rect 1035 1224 1101 1236
rect 1035 248 1051 1224
rect 1085 248 1101 1224
rect 1035 236 1101 248
rect 1131 1224 1197 1236
rect 1131 248 1147 1224
rect 1181 248 1197 1224
rect 1131 236 1197 248
rect 1227 1224 1289 1236
rect 1227 248 1243 1224
rect 1277 248 1289 1224
rect 1227 236 1289 248
rect 1361 1224 1423 1236
rect 1361 248 1373 1224
rect 1407 248 1423 1224
rect 1361 236 1423 248
rect 1453 1224 1519 1236
rect 1453 248 1469 1224
rect 1503 248 1519 1224
rect 1453 236 1519 248
rect 1549 1224 1615 1236
rect 1549 248 1565 1224
rect 1599 248 1615 1224
rect 1549 236 1615 248
rect 1645 1224 1711 1236
rect 1645 248 1661 1224
rect 1695 248 1711 1224
rect 1645 236 1711 248
rect 1741 1224 1807 1236
rect 1741 248 1757 1224
rect 1791 248 1807 1224
rect 1741 236 1807 248
rect 1837 1224 1903 1236
rect 1837 248 1853 1224
rect 1887 248 1903 1224
rect 1837 236 1903 248
rect 1933 1224 1999 1236
rect 1933 248 1949 1224
rect 1983 248 1999 1224
rect 1933 236 1999 248
rect 2029 1224 2095 1236
rect 2029 248 2045 1224
rect 2079 248 2095 1224
rect 2029 236 2095 248
rect 2125 1224 2191 1236
rect 2125 248 2141 1224
rect 2175 248 2191 1224
rect 2125 236 2191 248
rect 2221 1224 2287 1236
rect 2221 248 2237 1224
rect 2271 248 2287 1224
rect 2221 236 2287 248
rect 2317 1224 2383 1236
rect 2317 248 2333 1224
rect 2367 248 2383 1224
rect 2317 236 2383 248
rect 2413 1224 2479 1236
rect 2413 248 2429 1224
rect 2463 248 2479 1224
rect 2413 236 2479 248
rect 2509 1224 2575 1236
rect 2509 248 2525 1224
rect 2559 248 2575 1224
rect 2509 236 2575 248
rect 2605 1224 2671 1236
rect 2605 248 2621 1224
rect 2655 248 2671 1224
rect 2605 236 2671 248
rect 2701 1224 2767 1236
rect 2701 248 2717 1224
rect 2751 248 2767 1224
rect 2701 236 2767 248
rect 2797 1224 2863 1236
rect 2797 248 2813 1224
rect 2847 248 2863 1224
rect 2797 236 2863 248
rect 2893 1224 2959 1236
rect 2893 248 2909 1224
rect 2943 248 2959 1224
rect 2893 236 2959 248
rect 2989 1224 3055 1236
rect 2989 248 3005 1224
rect 3039 248 3055 1224
rect 2989 236 3055 248
rect 3085 1224 3151 1236
rect 3085 248 3101 1224
rect 3135 248 3151 1224
rect 3085 236 3151 248
rect 3181 1224 3247 1236
rect 3181 248 3197 1224
rect 3231 248 3247 1224
rect 3181 236 3247 248
rect 3277 1224 3343 1236
rect 3277 248 3293 1224
rect 3327 248 3343 1224
rect 3277 236 3343 248
rect 3373 1224 3439 1236
rect 3373 248 3389 1224
rect 3423 248 3439 1224
rect 3373 236 3439 248
rect 3469 1224 3535 1236
rect 3469 248 3485 1224
rect 3519 248 3535 1224
rect 3469 236 3535 248
rect 3565 1224 3631 1236
rect 3565 248 3581 1224
rect 3615 248 3631 1224
rect 3565 236 3631 248
rect 3661 1224 3727 1236
rect 3661 248 3677 1224
rect 3711 248 3727 1224
rect 3661 236 3727 248
rect 3757 1224 3823 1236
rect 3757 248 3773 1224
rect 3807 248 3823 1224
rect 3757 236 3823 248
rect 3853 1224 3919 1236
rect 3853 248 3869 1224
rect 3903 248 3919 1224
rect 3853 236 3919 248
rect 3949 1224 4015 1236
rect 3949 248 3965 1224
rect 3999 248 4015 1224
rect 3949 236 4015 248
rect 4045 1224 4111 1236
rect 4045 248 4061 1224
rect 4095 248 4111 1224
rect 4045 236 4111 248
rect 4141 1224 4207 1236
rect 4141 248 4157 1224
rect 4191 248 4207 1224
rect 4141 236 4207 248
rect 4237 1224 4303 1236
rect 4237 248 4253 1224
rect 4287 248 4303 1224
rect 4237 236 4303 248
rect 4333 1224 4399 1236
rect 4333 248 4349 1224
rect 4383 248 4399 1224
rect 4333 236 4399 248
rect 4429 1224 4495 1236
rect 4429 248 4445 1224
rect 4479 248 4495 1224
rect 4429 236 4495 248
rect 4525 1224 4591 1236
rect 4525 248 4541 1224
rect 4575 248 4591 1224
rect 4525 236 4591 248
rect 4621 1224 4687 1236
rect 4621 248 4637 1224
rect 4671 248 4687 1224
rect 4621 236 4687 248
rect 4717 1224 4783 1236
rect 4717 248 4733 1224
rect 4767 248 4783 1224
rect 4717 236 4783 248
rect 4813 1224 4875 1236
rect 4813 248 4829 1224
rect 4863 248 4875 1224
rect 4813 236 4875 248
<< ndiffc >>
rect 169 -498 203 -22
rect 265 -498 299 -22
rect 361 -498 395 -22
rect 475 -498 509 -22
rect 571 -498 605 -22
rect 667 -498 701 -22
rect 763 -498 797 -22
rect 859 -498 893 -22
rect 955 -498 989 -22
rect 1051 -498 1085 -22
rect 1147 -498 1181 -22
rect 1243 -498 1277 -22
rect 1373 -498 1407 -22
rect 1469 -498 1503 -22
rect 1565 -498 1599 -22
rect 1661 -498 1695 -22
rect 1757 -498 1791 -22
rect 1853 -498 1887 -22
rect 1949 -498 1983 -22
rect 2045 -498 2079 -22
rect 2141 -498 2175 -22
rect 2237 -498 2271 -22
rect 2333 -498 2367 -22
rect 2429 -498 2463 -22
rect 2525 -498 2559 -22
rect 2621 -498 2655 -22
rect 2717 -498 2751 -22
rect 2813 -498 2847 -22
rect 2909 -498 2943 -22
rect 3005 -498 3039 -22
rect 3101 -498 3135 -22
rect 3197 -498 3231 -22
rect 3293 -498 3327 -22
rect 3389 -498 3423 -22
rect 3485 -498 3519 -22
rect 3581 -498 3615 -22
rect 3677 -498 3711 -22
rect 3773 -498 3807 -22
rect 3869 -498 3903 -22
rect 3965 -498 3999 -22
rect 4061 -498 4095 -22
rect 4157 -498 4191 -22
rect 4253 -498 4287 -22
rect 4349 -498 4383 -22
rect 4445 -498 4479 -22
rect 4541 -498 4575 -22
rect 4637 -498 4671 -22
rect 4733 -498 4767 -22
rect 4829 -498 4863 -22
<< pdiffc >>
rect 169 246 203 1222
rect 265 246 299 1222
rect 361 246 395 1222
rect 475 248 509 1224
rect 571 248 605 1224
rect 667 248 701 1224
rect 763 248 797 1224
rect 859 248 893 1224
rect 955 248 989 1224
rect 1051 248 1085 1224
rect 1147 248 1181 1224
rect 1243 248 1277 1224
rect 1373 248 1407 1224
rect 1469 248 1503 1224
rect 1565 248 1599 1224
rect 1661 248 1695 1224
rect 1757 248 1791 1224
rect 1853 248 1887 1224
rect 1949 248 1983 1224
rect 2045 248 2079 1224
rect 2141 248 2175 1224
rect 2237 248 2271 1224
rect 2333 248 2367 1224
rect 2429 248 2463 1224
rect 2525 248 2559 1224
rect 2621 248 2655 1224
rect 2717 248 2751 1224
rect 2813 248 2847 1224
rect 2909 248 2943 1224
rect 3005 248 3039 1224
rect 3101 248 3135 1224
rect 3197 248 3231 1224
rect 3293 248 3327 1224
rect 3389 248 3423 1224
rect 3485 248 3519 1224
rect 3581 248 3615 1224
rect 3677 248 3711 1224
rect 3773 248 3807 1224
rect 3869 248 3903 1224
rect 3965 248 3999 1224
rect 4061 248 4095 1224
rect 4157 248 4191 1224
rect 4253 248 4287 1224
rect 4349 248 4383 1224
rect 4445 248 4479 1224
rect 4541 248 4575 1224
rect 4637 248 4671 1224
rect 4733 248 4767 1224
rect 4829 248 4863 1224
<< poly >>
rect 219 1234 249 1260
rect 315 1234 345 1260
rect 525 1236 555 1262
rect 621 1236 651 1262
rect 717 1236 747 1262
rect 813 1236 843 1262
rect 909 1236 939 1262
rect 1005 1236 1035 1262
rect 1101 1236 1131 1262
rect 1197 1236 1227 1262
rect 1423 1236 1453 1262
rect 1519 1236 1549 1262
rect 1615 1236 1645 1262
rect 1711 1236 1741 1262
rect 1807 1236 1837 1262
rect 1903 1236 1933 1262
rect 1999 1236 2029 1262
rect 2095 1236 2125 1262
rect 2191 1236 2221 1262
rect 2287 1236 2317 1262
rect 2383 1236 2413 1262
rect 2479 1236 2509 1262
rect 2575 1236 2605 1262
rect 2671 1236 2701 1262
rect 2767 1236 2797 1262
rect 2863 1236 2893 1262
rect 2959 1236 2989 1262
rect 3055 1236 3085 1262
rect 3151 1236 3181 1262
rect 3247 1236 3277 1262
rect 3343 1236 3373 1262
rect 3439 1236 3469 1262
rect 3535 1236 3565 1262
rect 3631 1236 3661 1262
rect 3727 1236 3757 1262
rect 3823 1236 3853 1262
rect 3919 1236 3949 1262
rect 4015 1236 4045 1262
rect 4111 1236 4141 1262
rect 4207 1236 4237 1262
rect 4303 1236 4333 1262
rect 4399 1236 4429 1262
rect 4495 1236 4525 1262
rect 4591 1236 4621 1262
rect 4687 1236 4717 1262
rect 4783 1236 4813 1262
rect 219 143 249 234
rect 315 143 345 234
rect 157 121 345 143
rect 157 99 182 121
rect 203 99 345 121
rect 157 77 345 99
rect 219 -10 249 77
rect 315 -10 345 77
rect 525 163 555 236
rect 621 163 651 236
rect 717 163 747 236
rect 813 163 843 236
rect 909 163 939 236
rect 1005 163 1035 236
rect 1101 163 1131 236
rect 1197 163 1227 236
rect 525 124 1227 163
rect 525 102 583 124
rect 1170 102 1227 124
rect 525 48 1227 102
rect 525 -10 555 48
rect 621 -10 651 48
rect 717 -10 747 48
rect 813 -10 843 48
rect 909 -10 939 48
rect 1005 -10 1035 48
rect 1101 -10 1131 48
rect 1197 -10 1227 48
rect 1423 210 1453 236
rect 1519 210 1549 236
rect 1615 210 1645 236
rect 1711 210 1741 236
rect 1807 210 1837 236
rect 1903 210 1933 236
rect 1999 210 2029 236
rect 2095 210 2125 236
rect 2191 210 2221 236
rect 2287 210 2317 236
rect 2383 210 2413 236
rect 2479 210 2509 236
rect 2575 210 2605 236
rect 2671 210 2701 236
rect 2767 210 2797 236
rect 2863 210 2893 236
rect 2959 210 2989 236
rect 3055 210 3085 236
rect 3151 210 3181 236
rect 3247 210 3277 236
rect 3343 210 3373 236
rect 3439 210 3469 236
rect 3535 210 3565 236
rect 3631 210 3661 236
rect 3727 210 3757 236
rect 3823 210 3853 236
rect 3919 210 3949 236
rect 4015 210 4045 236
rect 4111 210 4141 236
rect 4207 210 4237 236
rect 4303 210 4333 236
rect 4399 210 4429 236
rect 4495 210 4525 236
rect 4591 210 4621 236
rect 4687 210 4717 236
rect 4783 210 4813 236
rect 1423 124 4813 210
rect 1423 102 1581 124
rect 1423 101 4581 102
rect 4716 101 4813 124
rect 1423 16 4813 101
rect 1423 -10 1453 16
rect 1519 -10 1549 16
rect 1615 -10 1645 16
rect 1711 -10 1741 16
rect 1807 -10 1837 16
rect 1903 -10 1933 16
rect 1999 -10 2029 16
rect 2095 -10 2125 16
rect 2191 -10 2221 16
rect 2287 -10 2317 16
rect 2383 -10 2413 16
rect 2479 -10 2509 16
rect 2575 -10 2605 16
rect 2671 -10 2701 16
rect 2767 -10 2797 16
rect 2863 -10 2893 16
rect 2959 -10 2989 16
rect 3055 -10 3085 16
rect 3151 -10 3181 16
rect 3247 -10 3277 16
rect 3343 -10 3373 16
rect 3439 -10 3469 16
rect 3535 -10 3565 16
rect 3631 -10 3661 16
rect 3727 -10 3757 16
rect 3823 -10 3853 16
rect 3919 -10 3949 16
rect 4015 -10 4045 16
rect 4111 -10 4141 16
rect 4207 -10 4237 16
rect 4303 -10 4333 16
rect 4399 -10 4429 16
rect 4495 -10 4525 16
rect 4591 -10 4621 16
rect 4687 -10 4717 16
rect 4783 -10 4813 16
rect 219 -536 249 -510
rect 315 -536 345 -510
rect 525 -536 555 -510
rect 621 -536 651 -510
rect 717 -536 747 -510
rect 813 -536 843 -510
rect 909 -536 939 -510
rect 1005 -536 1035 -510
rect 1101 -536 1131 -510
rect 1197 -536 1227 -510
rect 1423 -536 1453 -510
rect 1519 -536 1549 -510
rect 1615 -536 1645 -510
rect 1711 -536 1741 -510
rect 1807 -536 1837 -510
rect 1903 -536 1933 -510
rect 1999 -536 2029 -510
rect 2095 -536 2125 -510
rect 2191 -536 2221 -510
rect 2287 -536 2317 -510
rect 2383 -536 2413 -510
rect 2479 -536 2509 -510
rect 2575 -536 2605 -510
rect 2671 -536 2701 -510
rect 2767 -536 2797 -510
rect 2863 -536 2893 -510
rect 2959 -536 2989 -510
rect 3055 -536 3085 -510
rect 3151 -536 3181 -510
rect 3247 -536 3277 -510
rect 3343 -536 3373 -510
rect 3439 -536 3469 -510
rect 3535 -536 3565 -510
rect 3631 -536 3661 -510
rect 3727 -536 3757 -510
rect 3823 -536 3853 -510
rect 3919 -536 3949 -510
rect 4015 -536 4045 -510
rect 4111 -536 4141 -510
rect 4207 -536 4237 -510
rect 4303 -536 4333 -510
rect 4399 -536 4429 -510
rect 4495 -536 4525 -510
rect 4591 -536 4621 -510
rect 4687 -536 4717 -510
rect 4783 -536 4813 -510
<< polycont >>
rect 182 99 203 121
rect 583 102 1170 124
rect 1581 102 4716 124
rect 4581 101 4716 102
<< locali >>
rect 169 1276 395 1310
rect 169 1222 203 1276
rect 169 230 203 246
rect 265 1222 299 1238
rect 167 121 219 137
rect 167 99 182 121
rect 203 99 219 121
rect 167 83 219 99
rect 265 130 299 246
rect 361 1222 395 1276
rect 361 230 395 246
rect 475 1276 1277 1310
rect 475 1224 509 1276
rect 475 232 509 248
rect 571 1224 605 1240
rect 571 198 605 248
rect 667 1224 701 1276
rect 667 232 701 248
rect 763 1224 797 1240
rect 763 198 797 248
rect 859 1224 893 1276
rect 859 232 893 248
rect 955 1224 989 1240
rect 955 198 989 248
rect 1051 1224 1085 1276
rect 1051 232 1085 248
rect 1147 1224 1181 1240
rect 1147 198 1181 248
rect 1243 1224 1277 1276
rect 1243 232 1277 248
rect 1373 1276 4863 1310
rect 1373 1224 1407 1276
rect 1373 232 1407 248
rect 1469 1224 1503 1240
rect 1469 198 1503 248
rect 1565 1224 1599 1276
rect 1565 232 1599 248
rect 1661 1224 1695 1240
rect 1661 198 1695 248
rect 1757 1224 1791 1276
rect 1757 232 1791 248
rect 1853 1224 1887 1240
rect 1853 198 1887 248
rect 1949 1224 1983 1276
rect 1949 232 1983 248
rect 2045 1224 2079 1240
rect 2045 198 2079 248
rect 2141 1224 2175 1276
rect 2141 232 2175 248
rect 2237 1224 2271 1240
rect 2237 198 2271 248
rect 2333 1224 2367 1276
rect 2333 232 2367 248
rect 2429 1224 2463 1240
rect 2429 198 2463 248
rect 2525 1224 2559 1276
rect 2525 232 2559 248
rect 2621 1224 2655 1240
rect 2621 198 2655 248
rect 2717 1224 2751 1276
rect 2717 232 2751 248
rect 2813 1224 2847 1240
rect 2813 198 2847 248
rect 2909 1224 2943 1276
rect 2909 232 2943 248
rect 3005 1224 3039 1240
rect 3005 198 3039 248
rect 3101 1224 3135 1276
rect 3101 232 3135 248
rect 3197 1224 3231 1240
rect 3197 198 3231 248
rect 3293 1224 3327 1276
rect 3293 232 3327 248
rect 3389 1224 3423 1240
rect 3389 198 3423 248
rect 3485 1224 3519 1276
rect 3485 232 3519 248
rect 3581 1224 3615 1240
rect 3581 198 3615 248
rect 3677 1224 3711 1276
rect 3677 232 3711 248
rect 3773 1224 3807 1240
rect 3773 198 3807 248
rect 3869 1224 3903 1276
rect 3869 232 3903 248
rect 3965 1224 3999 1240
rect 3965 198 3999 248
rect 4061 1224 4095 1276
rect 4061 232 4095 248
rect 4157 1224 4191 1240
rect 4157 198 4191 248
rect 4253 1224 4287 1276
rect 4253 232 4287 248
rect 4349 1224 4383 1240
rect 4349 198 4383 248
rect 4445 1224 4479 1276
rect 4445 232 4479 248
rect 4541 1224 4575 1240
rect 4541 198 4575 248
rect 4637 1224 4671 1276
rect 4637 232 4671 248
rect 4733 1224 4767 1240
rect 4733 198 4767 248
rect 4829 1224 4863 1276
rect 4829 232 4863 248
rect 571 164 1270 198
rect 1469 164 4841 198
rect 1236 130 1270 164
rect 265 124 1186 130
rect 265 102 583 124
rect 1170 102 1186 124
rect 265 96 1186 102
rect 1236 124 4747 130
rect 1236 102 1581 124
rect 1236 101 4581 102
rect 4716 101 4747 124
rect 1236 96 4747 101
rect 169 -22 203 -6
rect 169 -548 203 -498
rect 265 -22 299 96
rect 1236 62 1270 96
rect 4804 62 4841 164
rect 571 28 1270 62
rect 1469 28 4841 62
rect 265 -514 299 -498
rect 361 -22 395 -6
rect 361 -548 395 -498
rect 169 -582 395 -548
rect 475 -22 509 -6
rect 475 -548 509 -498
rect 571 -22 605 28
rect 571 -514 605 -498
rect 667 -22 701 -6
rect 667 -548 701 -498
rect 763 -22 797 28
rect 763 -514 797 -498
rect 859 -22 893 -6
rect 859 -548 893 -498
rect 955 -22 989 28
rect 955 -514 989 -498
rect 1051 -22 1085 -6
rect 1051 -548 1085 -498
rect 1147 -22 1181 28
rect 1147 -514 1181 -498
rect 1243 -22 1277 -6
rect 1243 -548 1277 -498
rect 475 -582 1277 -548
rect 1373 -22 1407 -6
rect 1373 -550 1407 -498
rect 1469 -22 1503 28
rect 1469 -514 1503 -498
rect 1565 -22 1599 -6
rect 1565 -550 1599 -498
rect 1661 -22 1695 28
rect 1661 -514 1695 -498
rect 1757 -22 1791 -6
rect 1757 -550 1791 -498
rect 1853 -22 1887 28
rect 1853 -514 1887 -498
rect 1949 -22 1983 -6
rect 1949 -550 1983 -498
rect 2045 -22 2079 28
rect 2045 -514 2079 -498
rect 2141 -22 2175 -6
rect 2141 -550 2175 -498
rect 2237 -22 2271 28
rect 2237 -514 2271 -498
rect 2333 -22 2367 -6
rect 2333 -550 2367 -498
rect 2429 -22 2463 28
rect 2429 -514 2463 -498
rect 2525 -22 2559 -6
rect 2525 -550 2559 -498
rect 2621 -22 2655 28
rect 2621 -514 2655 -498
rect 2717 -22 2751 -6
rect 2717 -550 2751 -498
rect 2813 -22 2847 28
rect 2813 -514 2847 -498
rect 2909 -22 2943 -6
rect 2909 -550 2943 -498
rect 3005 -22 3039 28
rect 3005 -514 3039 -498
rect 3101 -22 3135 -6
rect 3101 -550 3135 -498
rect 3197 -22 3231 28
rect 3197 -514 3231 -498
rect 3293 -22 3327 -6
rect 3293 -550 3327 -498
rect 3389 -22 3423 28
rect 3389 -514 3423 -498
rect 3485 -22 3519 -6
rect 3485 -550 3519 -498
rect 3581 -22 3615 28
rect 3581 -514 3615 -498
rect 3677 -22 3711 -6
rect 3677 -550 3711 -498
rect 3773 -22 3807 28
rect 3773 -514 3807 -498
rect 3869 -22 3903 -6
rect 3869 -550 3903 -498
rect 3965 -22 3999 28
rect 3965 -514 3999 -498
rect 4061 -22 4095 -6
rect 4061 -550 4095 -498
rect 4157 -22 4191 28
rect 4157 -514 4191 -498
rect 4253 -22 4287 -6
rect 4253 -550 4287 -498
rect 4349 -22 4383 28
rect 4349 -514 4383 -498
rect 4445 -22 4479 -6
rect 4445 -550 4479 -498
rect 4541 -22 4575 28
rect 4541 -514 4575 -498
rect 4637 -22 4671 -6
rect 4637 -550 4671 -498
rect 4733 -22 4767 28
rect 4733 -514 4767 -498
rect 4829 -22 4863 -6
rect 4829 -550 4863 -498
rect 1373 -584 4863 -550
<< viali >>
rect 169 246 203 1222
rect 265 246 299 1222
rect 361 246 395 1222
rect 475 248 509 1224
rect 571 248 605 1224
rect 667 248 701 1224
rect 763 248 797 1224
rect 859 248 893 1224
rect 955 248 989 1224
rect 1051 248 1085 1224
rect 1147 248 1181 1224
rect 1243 248 1277 1224
rect 1373 248 1407 1224
rect 1469 248 1503 1224
rect 1565 248 1599 1224
rect 1661 248 1695 1224
rect 1757 248 1791 1224
rect 1853 248 1887 1224
rect 1949 248 1983 1224
rect 2045 248 2079 1224
rect 2141 248 2175 1224
rect 2237 248 2271 1224
rect 2333 248 2367 1224
rect 2429 248 2463 1224
rect 2525 248 2559 1224
rect 2621 248 2655 1224
rect 2717 248 2751 1224
rect 2813 248 2847 1224
rect 2909 248 2943 1224
rect 3005 248 3039 1224
rect 3101 248 3135 1224
rect 3197 248 3231 1224
rect 3293 248 3327 1224
rect 3389 248 3423 1224
rect 3485 248 3519 1224
rect 3581 248 3615 1224
rect 3677 248 3711 1224
rect 3773 248 3807 1224
rect 3869 248 3903 1224
rect 3965 248 3999 1224
rect 4061 248 4095 1224
rect 4157 248 4191 1224
rect 4253 248 4287 1224
rect 4349 248 4383 1224
rect 4445 248 4479 1224
rect 4541 248 4575 1224
rect 4637 248 4671 1224
rect 4733 248 4767 1224
rect 4829 248 4863 1224
rect 169 -498 203 -22
rect 265 -498 299 -22
rect 361 -498 395 -22
rect 475 -498 509 -22
rect 571 -498 605 -22
rect 667 -498 701 -22
rect 763 -498 797 -22
rect 859 -498 893 -22
rect 955 -498 989 -22
rect 1051 -498 1085 -22
rect 1147 -498 1181 -22
rect 1243 -498 1277 -22
rect 1373 -498 1407 -22
rect 1469 -498 1503 -22
rect 1565 -498 1599 -22
rect 1661 -498 1695 -22
rect 1757 -498 1791 -22
rect 1853 -498 1887 -22
rect 1949 -498 1983 -22
rect 2045 -498 2079 -22
rect 2141 -498 2175 -22
rect 2237 -498 2271 -22
rect 2333 -498 2367 -22
rect 2429 -498 2463 -22
rect 2525 -498 2559 -22
rect 2621 -498 2655 -22
rect 2717 -498 2751 -22
rect 2813 -498 2847 -22
rect 2909 -498 2943 -22
rect 3005 -498 3039 -22
rect 3101 -498 3135 -22
rect 3197 -498 3231 -22
rect 3293 -498 3327 -22
rect 3389 -498 3423 -22
rect 3485 -498 3519 -22
rect 3581 -498 3615 -22
rect 3677 -498 3711 -22
rect 3773 -498 3807 -22
rect 3869 -498 3903 -22
rect 3965 -498 3999 -22
rect 4061 -498 4095 -22
rect 4157 -498 4191 -22
rect 4253 -498 4287 -22
rect 4349 -498 4383 -22
rect 4445 -498 4479 -22
rect 4541 -498 4575 -22
rect 4637 -498 4671 -22
rect 4733 -498 4767 -22
rect 4829 -498 4863 -22
<< metal1 >>
rect 163 1222 209 1234
rect 163 246 169 1222
rect 203 246 209 1222
rect 163 234 209 246
rect 259 1222 305 1234
rect 259 246 265 1222
rect 299 246 305 1222
rect 259 234 305 246
rect 355 1222 401 1234
rect 355 246 361 1222
rect 395 246 401 1222
rect 355 234 401 246
rect 469 1224 515 1236
rect 469 248 475 1224
rect 509 248 515 1224
rect 469 236 515 248
rect 565 1224 611 1236
rect 565 248 571 1224
rect 605 248 611 1224
rect 565 236 611 248
rect 661 1224 707 1236
rect 661 248 667 1224
rect 701 248 707 1224
rect 661 236 707 248
rect 757 1224 803 1236
rect 757 248 763 1224
rect 797 248 803 1224
rect 757 236 803 248
rect 853 1224 899 1236
rect 853 248 859 1224
rect 893 248 899 1224
rect 853 236 899 248
rect 949 1224 995 1236
rect 949 248 955 1224
rect 989 248 995 1224
rect 949 236 995 248
rect 1045 1224 1091 1236
rect 1045 248 1051 1224
rect 1085 248 1091 1224
rect 1045 236 1091 248
rect 1141 1224 1187 1236
rect 1141 248 1147 1224
rect 1181 248 1187 1224
rect 1141 236 1187 248
rect 1237 1224 1283 1236
rect 1237 248 1243 1224
rect 1277 248 1283 1224
rect 1237 236 1283 248
rect 1367 1224 1413 1236
rect 1367 248 1373 1224
rect 1407 248 1413 1224
rect 1367 236 1413 248
rect 1463 1224 1509 1236
rect 1463 248 1469 1224
rect 1503 248 1509 1224
rect 1463 236 1509 248
rect 1559 1224 1605 1236
rect 1559 248 1565 1224
rect 1599 248 1605 1224
rect 1559 236 1605 248
rect 1655 1224 1701 1236
rect 1655 248 1661 1224
rect 1695 248 1701 1224
rect 1655 236 1701 248
rect 1751 1224 1797 1236
rect 1751 248 1757 1224
rect 1791 248 1797 1224
rect 1751 236 1797 248
rect 1847 1224 1893 1236
rect 1847 248 1853 1224
rect 1887 248 1893 1224
rect 1847 236 1893 248
rect 1943 1224 1989 1236
rect 1943 248 1949 1224
rect 1983 248 1989 1224
rect 1943 236 1989 248
rect 2039 1224 2085 1236
rect 2039 248 2045 1224
rect 2079 248 2085 1224
rect 2039 236 2085 248
rect 2135 1224 2181 1236
rect 2135 248 2141 1224
rect 2175 248 2181 1224
rect 2135 236 2181 248
rect 2231 1224 2277 1236
rect 2231 248 2237 1224
rect 2271 248 2277 1224
rect 2231 236 2277 248
rect 2327 1224 2373 1236
rect 2327 248 2333 1224
rect 2367 248 2373 1224
rect 2327 236 2373 248
rect 2423 1224 2469 1236
rect 2423 248 2429 1224
rect 2463 248 2469 1224
rect 2423 236 2469 248
rect 2519 1224 2565 1236
rect 2519 248 2525 1224
rect 2559 248 2565 1224
rect 2519 236 2565 248
rect 2615 1224 2661 1236
rect 2615 248 2621 1224
rect 2655 248 2661 1224
rect 2615 236 2661 248
rect 2711 1224 2757 1236
rect 2711 248 2717 1224
rect 2751 248 2757 1224
rect 2711 236 2757 248
rect 2807 1224 2853 1236
rect 2807 248 2813 1224
rect 2847 248 2853 1224
rect 2807 236 2853 248
rect 2903 1224 2949 1236
rect 2903 248 2909 1224
rect 2943 248 2949 1224
rect 2903 236 2949 248
rect 2999 1224 3045 1236
rect 2999 248 3005 1224
rect 3039 248 3045 1224
rect 2999 236 3045 248
rect 3095 1224 3141 1236
rect 3095 248 3101 1224
rect 3135 248 3141 1224
rect 3095 236 3141 248
rect 3191 1224 3237 1236
rect 3191 248 3197 1224
rect 3231 248 3237 1224
rect 3191 236 3237 248
rect 3287 1224 3333 1236
rect 3287 248 3293 1224
rect 3327 248 3333 1224
rect 3287 236 3333 248
rect 3383 1224 3429 1236
rect 3383 248 3389 1224
rect 3423 248 3429 1224
rect 3383 236 3429 248
rect 3479 1224 3525 1236
rect 3479 248 3485 1224
rect 3519 248 3525 1224
rect 3479 236 3525 248
rect 3575 1224 3621 1236
rect 3575 248 3581 1224
rect 3615 248 3621 1224
rect 3575 236 3621 248
rect 3671 1224 3717 1236
rect 3671 248 3677 1224
rect 3711 248 3717 1224
rect 3671 236 3717 248
rect 3767 1224 3813 1236
rect 3767 248 3773 1224
rect 3807 248 3813 1224
rect 3767 236 3813 248
rect 3863 1224 3909 1236
rect 3863 248 3869 1224
rect 3903 248 3909 1224
rect 3863 236 3909 248
rect 3959 1224 4005 1236
rect 3959 248 3965 1224
rect 3999 248 4005 1224
rect 3959 236 4005 248
rect 4055 1224 4101 1236
rect 4055 248 4061 1224
rect 4095 248 4101 1224
rect 4055 236 4101 248
rect 4151 1224 4197 1236
rect 4151 248 4157 1224
rect 4191 248 4197 1224
rect 4151 236 4197 248
rect 4247 1224 4293 1236
rect 4247 248 4253 1224
rect 4287 248 4293 1224
rect 4247 236 4293 248
rect 4343 1224 4389 1236
rect 4343 248 4349 1224
rect 4383 248 4389 1224
rect 4343 236 4389 248
rect 4439 1224 4485 1236
rect 4439 248 4445 1224
rect 4479 248 4485 1224
rect 4439 236 4485 248
rect 4535 1224 4581 1236
rect 4535 248 4541 1224
rect 4575 248 4581 1224
rect 4535 236 4581 248
rect 4631 1224 4677 1236
rect 4631 248 4637 1224
rect 4671 248 4677 1224
rect 4631 236 4677 248
rect 4727 1224 4773 1236
rect 4727 248 4733 1224
rect 4767 248 4773 1224
rect 4727 236 4773 248
rect 4823 1224 4869 1236
rect 4823 248 4829 1224
rect 4863 248 4869 1224
rect 4823 236 4869 248
rect 163 -22 209 -10
rect 163 -498 169 -22
rect 203 -498 209 -22
rect 163 -510 209 -498
rect 259 -22 305 -10
rect 259 -498 265 -22
rect 299 -498 305 -22
rect 259 -510 305 -498
rect 355 -22 401 -10
rect 355 -498 361 -22
rect 395 -498 401 -22
rect 355 -510 401 -498
rect 469 -22 515 -10
rect 469 -498 475 -22
rect 509 -498 515 -22
rect 469 -510 515 -498
rect 565 -22 611 -10
rect 565 -498 571 -22
rect 605 -498 611 -22
rect 565 -510 611 -498
rect 661 -22 707 -10
rect 661 -498 667 -22
rect 701 -498 707 -22
rect 661 -510 707 -498
rect 757 -22 803 -10
rect 757 -498 763 -22
rect 797 -498 803 -22
rect 757 -510 803 -498
rect 853 -22 899 -10
rect 853 -498 859 -22
rect 893 -498 899 -22
rect 853 -510 899 -498
rect 949 -22 995 -10
rect 949 -498 955 -22
rect 989 -498 995 -22
rect 949 -510 995 -498
rect 1045 -22 1091 -10
rect 1045 -498 1051 -22
rect 1085 -498 1091 -22
rect 1045 -510 1091 -498
rect 1141 -22 1187 -10
rect 1141 -498 1147 -22
rect 1181 -498 1187 -22
rect 1141 -510 1187 -498
rect 1237 -22 1283 -10
rect 1237 -498 1243 -22
rect 1277 -498 1283 -22
rect 1237 -510 1283 -498
rect 1367 -22 1413 -10
rect 1367 -498 1373 -22
rect 1407 -498 1413 -22
rect 1367 -510 1413 -498
rect 1463 -22 1509 -10
rect 1463 -498 1469 -22
rect 1503 -498 1509 -22
rect 1463 -510 1509 -498
rect 1559 -22 1605 -10
rect 1559 -498 1565 -22
rect 1599 -498 1605 -22
rect 1559 -510 1605 -498
rect 1655 -22 1701 -10
rect 1655 -498 1661 -22
rect 1695 -498 1701 -22
rect 1655 -510 1701 -498
rect 1751 -22 1797 -10
rect 1751 -498 1757 -22
rect 1791 -498 1797 -22
rect 1751 -510 1797 -498
rect 1847 -22 1893 -10
rect 1847 -498 1853 -22
rect 1887 -498 1893 -22
rect 1847 -510 1893 -498
rect 1943 -22 1989 -10
rect 1943 -498 1949 -22
rect 1983 -498 1989 -22
rect 1943 -510 1989 -498
rect 2039 -22 2085 -10
rect 2039 -498 2045 -22
rect 2079 -498 2085 -22
rect 2039 -510 2085 -498
rect 2135 -22 2181 -10
rect 2135 -498 2141 -22
rect 2175 -498 2181 -22
rect 2135 -510 2181 -498
rect 2231 -22 2277 -10
rect 2231 -498 2237 -22
rect 2271 -498 2277 -22
rect 2231 -510 2277 -498
rect 2327 -22 2373 -10
rect 2327 -498 2333 -22
rect 2367 -498 2373 -22
rect 2327 -510 2373 -498
rect 2423 -22 2469 -10
rect 2423 -498 2429 -22
rect 2463 -498 2469 -22
rect 2423 -510 2469 -498
rect 2519 -22 2565 -10
rect 2519 -498 2525 -22
rect 2559 -498 2565 -22
rect 2519 -510 2565 -498
rect 2615 -22 2661 -10
rect 2615 -498 2621 -22
rect 2655 -498 2661 -22
rect 2615 -510 2661 -498
rect 2711 -22 2757 -10
rect 2711 -498 2717 -22
rect 2751 -498 2757 -22
rect 2711 -510 2757 -498
rect 2807 -22 2853 -10
rect 2807 -498 2813 -22
rect 2847 -498 2853 -22
rect 2807 -510 2853 -498
rect 2903 -22 2949 -10
rect 2903 -498 2909 -22
rect 2943 -498 2949 -22
rect 2903 -510 2949 -498
rect 2999 -22 3045 -10
rect 2999 -498 3005 -22
rect 3039 -498 3045 -22
rect 2999 -510 3045 -498
rect 3095 -22 3141 -10
rect 3095 -498 3101 -22
rect 3135 -498 3141 -22
rect 3095 -510 3141 -498
rect 3191 -22 3237 -10
rect 3191 -498 3197 -22
rect 3231 -498 3237 -22
rect 3191 -510 3237 -498
rect 3287 -22 3333 -10
rect 3287 -498 3293 -22
rect 3327 -498 3333 -22
rect 3287 -510 3333 -498
rect 3383 -22 3429 -10
rect 3383 -498 3389 -22
rect 3423 -498 3429 -22
rect 3383 -510 3429 -498
rect 3479 -22 3525 -10
rect 3479 -498 3485 -22
rect 3519 -498 3525 -22
rect 3479 -510 3525 -498
rect 3575 -22 3621 -10
rect 3575 -498 3581 -22
rect 3615 -498 3621 -22
rect 3575 -510 3621 -498
rect 3671 -22 3717 -10
rect 3671 -498 3677 -22
rect 3711 -498 3717 -22
rect 3671 -510 3717 -498
rect 3767 -22 3813 -10
rect 3767 -498 3773 -22
rect 3807 -498 3813 -22
rect 3767 -510 3813 -498
rect 3863 -22 3909 -10
rect 3863 -498 3869 -22
rect 3903 -498 3909 -22
rect 3863 -510 3909 -498
rect 3959 -22 4005 -10
rect 3959 -498 3965 -22
rect 3999 -498 4005 -22
rect 3959 -510 4005 -498
rect 4055 -22 4101 -10
rect 4055 -498 4061 -22
rect 4095 -498 4101 -22
rect 4055 -510 4101 -498
rect 4151 -22 4197 -10
rect 4151 -498 4157 -22
rect 4191 -498 4197 -22
rect 4151 -510 4197 -498
rect 4247 -22 4293 -10
rect 4247 -498 4253 -22
rect 4287 -498 4293 -22
rect 4247 -510 4293 -498
rect 4343 -22 4389 -10
rect 4343 -498 4349 -22
rect 4383 -498 4389 -22
rect 4343 -510 4389 -498
rect 4439 -22 4485 -10
rect 4439 -498 4445 -22
rect 4479 -498 4485 -22
rect 4439 -510 4485 -498
rect 4535 -22 4581 -10
rect 4535 -498 4541 -22
rect 4575 -498 4581 -22
rect 4535 -510 4581 -498
rect 4631 -22 4677 -10
rect 4631 -498 4637 -22
rect 4671 -498 4677 -22
rect 4631 -510 4677 -498
rect 4727 -22 4773 -10
rect 4727 -498 4733 -22
rect 4767 -498 4773 -22
rect 4727 -510 4773 -498
rect 4823 -22 4869 -10
rect 4823 -498 4829 -22
rect 4863 -498 4869 -22
rect 4823 -510 4869 -498
<< end >>
