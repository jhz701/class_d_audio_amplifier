* NGSPICE file created from /home/eda/magic/class_d_audio_amplifier/user_project_wrapper/user_analog_project_wrapper_empty_lvs.ext - technology: sky130A


* Top level circuit /home/eda/magic/class_d_audio_amplifier/user_project_wrapper/user_analog_project_wrapper_empty_lvs

X0 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5 a_3420293_704737# a_3424227_705357# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=2.8e+06u
X6 a_3361095_699281# a_3379272_706425# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X7 a_3369760_754598# a_3366260_744206# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X11 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X12 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X13 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X14 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X15 a_3400801_701658# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X16 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X17 a_3439418_744112# a_3442918_747574# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X18 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X19 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X20 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X21 w_3185490_798160# a_3381660_718033# a_3381660_718777# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X22 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X23 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X24 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X25 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X26 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X27 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X28 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X29 a_3407435_674425# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X30 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X31 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X32 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X33 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X34 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X35 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X36 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X37 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X38 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X39 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X40 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X41 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X42 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X43 w_3185490_798160# a_3403286_703346# a_3403286_703346# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X44 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X45 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X46 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X47 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X48 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X49 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X50 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X51 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X52 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X53 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X54 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X55 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X56 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X57 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X58 w_3185490_798160# a_3399027_674337# a_3401256_686207# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X59 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X60 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X61 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X62 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X63 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X64 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X65 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X66 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X67 w_3263498_541854# a_3379175_700273# w_3381441_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X68 a_3407542_688639# a_3381563_702505# w_3407323_687499# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X69 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X70 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X71 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X72 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X73 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X74 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X75 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X76 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X77 w_3185490_798160# a_3399027_674337# a_3399027_674337# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X78 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X79 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X80 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X81 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X82 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X83 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X84 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X85 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X86 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X87 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X88 a_3394410_690671# a_3263636_541992# w_3396510_687499# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X89 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X90 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X91 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X92 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X93 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X94 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X95 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X96 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X97 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X98 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X99 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X100 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X101 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X102 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X103 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X104 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X105 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X106 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X107 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X108 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X109 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X110 a_3335479_772599# a_3359810_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X111 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X112 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X113 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X114 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X115 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X116 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X117 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X118 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X119 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X120 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X121 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X122 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X123 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X124 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X125 w_3403067_702950# a_3381563_702505# a_3403286_704090# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X126 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X127 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X128 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X129 w_3381441_717637# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X130 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X131 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X132 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X133 a_3403001_699542# a_3403319_700774# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X134 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X135 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X136 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X137 w_3381441_717637# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X138 a_3403286_717614# a_3403286_716870# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X139 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X140 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X141 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X142 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X143 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X144 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X145 w_3263498_541854# a_3400801_701658# a_3400801_701658# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X146 a_3420294_717833# a_3420294_717833# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X147 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X148 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X149 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X150 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X151 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X152 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X153 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X154 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X155 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X156 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X157 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X158 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X159 a_3394410_690671# a_3394410_687695# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X160 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X161 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X162 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X163 a_3420293_701761# a_3422243_697443# w_3422393_701565# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X164 v2 a_3359810_749958# a_3335479_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X165 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X166 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X167 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X168 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X169 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X170 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X171 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X172 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X173 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X174 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X175 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X176 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X177 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X178 w_3263498_541854# a_3405057_686207# a_3405057_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X179 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X180 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X181 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X182 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X183 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X184 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
R0 a_3427310_772647# m3_3560250_970224# sky130_fd_pr__res_generic_m3 w=2.505e+07u l=3.7e+06u
X185 w_3381441_701565# a_3381563_702505# a_3381660_702705# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X186 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X187 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X188 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X189 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X190 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X191 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X192 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X193 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X194 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X195 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X196 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X197 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X198 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X199 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X200 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X201 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X202 a_3408579_674425# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X203 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
R1 a_3285528_930602# m3_3267050_970234# sky130_fd_pr__res_generic_m3 w=2.505e+07u l=7.55e+06u
X204 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X205 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X206 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X207 w_3185490_798160# a_3366260_744206# a_3369760_754598# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X208 w_3185490_798160# a_3359810_749958# a_3335479_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X209 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X210 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X211 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X212 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X213 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X214 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X215 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X216 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X217 w_3263498_541854# a_3408579_674425# w_3422394_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X218 a_3394410_687695# a_3394410_687695# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X219 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X220 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X221 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X222 w_3185490_798160# a_3407542_687895# a_3407542_688639# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X223 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X224 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X225 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X226 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X227 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X228 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X229 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X230 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X231 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X232 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X233 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X234 w_3263498_541854# a_3408579_674425# a_3408579_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X235 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X236 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X237 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X238 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X239 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X240 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X241 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X242 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X243 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X244 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X245 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X246 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X247 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X248 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X249 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X250 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X251 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X252 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X253 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X254 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X255 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X256 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X257 v2 a_3366260_744206# a_3369760_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X258 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X259 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X260 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X261 w_3381441_717637# a_3379272_706425# a_3381660_718777# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X262 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X263 a_3263636_541992# w_3263498_541854# sky130_fd_pr__diode_pd2nw_05v5 area=2.25e+16p
X264 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X265 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X266 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X267 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X268 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X269 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X270 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X271 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X272 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X273 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X274 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X275 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X276 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X277 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X278 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X279 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X280 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X281 w_3263498_541854# a_3401256_686207# w_3396510_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X282 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X283 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X284 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X285 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X286 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X287 a_3407542_688639# a_3381563_702505# w_3407323_687499# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X288 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X289 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X290 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X291 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X292 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X293 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X294 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X295 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X296 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X297 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X298 a_3394410_690671# a_3263636_541992# w_3396510_687499# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X299 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X300 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X301 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X302 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X303 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X304 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X305 a_3443016_749796# a_3439418_744112# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X306 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X307 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X308 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X309 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X310 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X311 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X312 a_3381563_702505# w_3474538_503344# sky130_fd_pr__diode_pd2nw_05v5 area=2.25e+16p
X313 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X314 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X315 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X316 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X317 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X318 a_3361095_699281# a_3379272_706425# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X319 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X320 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X321 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X322 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X323 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X324 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X325 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X326 a_3420294_717833# a_3381563_717833# w_3422394_717637# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X327 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X328 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X329 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X330 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X331 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X332 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X333 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X334 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X335 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X336 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X337 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X338 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X339 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X340 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X341 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X342 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X343 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X344 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X345 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X346 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X347 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X348 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X349 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X350 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X351 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X352 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X353 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X354 a_3381660_718033# a_3381660_718033# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X355 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X356 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X357 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X358 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X359 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X360 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X361 a_3386185_697443# a_3385867_698875# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X362 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X363 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X364 a_3420293_701761# a_3422243_697443# w_3422393_701565# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X365 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X366 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X367 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X368 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X369 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X370 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X371 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X372 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X373 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X374 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X375 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X376 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X377 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X378 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X379 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X380 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X381 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X382 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X383 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X384 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X385 w_3185490_798160# a_3420294_717833# a_3420294_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X386 w_3185490_798160# a_3435992_747994# a_3434368_749958# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X387 w_3185490_798160# a_3403286_716870# a_3403286_717614# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X388 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X389 w_3422394_717637# a_3420381_704937# a_3420294_720809# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X390 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X391 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X392 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X393 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X394 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X395 w_3263498_541854# a_3400801_701658# w_3403067_702950# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X396 a_3420294_720809# a_3420294_717833# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X397 w_3381441_717637# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X398 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X399 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X400 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X401 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X402 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X403 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X404 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X405 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X406 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X407 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X408 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X409 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X410 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X411 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X412 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X413 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X414 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X415 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X416 a_3428294_754598# a_3434368_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X417 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X418 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X419 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X420 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X421 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X422 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X423 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X424 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X425 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X426 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X427 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X428 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X429 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X430 w_3381441_701565# a_3361095_699281# a_3381660_701961# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X431 a_3420293_704737# a_3420293_701761# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X432 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X433 a_3381660_702705# a_3381660_701961# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X434 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X435 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X436 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X437 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X438 v2 a_3439418_744112# a_3443016_749796# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X439 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X440 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X441 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X442 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X443 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X444 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X445 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X446 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X447 w_3185490_798160# a_3394410_687695# a_3394410_687695# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X448 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X449 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X450 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X451 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X452 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X453 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X454 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X455 w_3381441_717637# a_3379272_706425# a_3381660_718777# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X456 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X457 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X458 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X459 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X460 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X461 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X462 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X463 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X464 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X465 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X466 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X467 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X468 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X469 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X470 a_3403286_716870# a_3403286_716870# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X471 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X472 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X473 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X474 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X475 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X476 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X477 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X478 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X479 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X480 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X481 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X482 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X483 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X484 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X485 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X486 a_3381660_701961# a_3381660_701961# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X487 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X488 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X489 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X490 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X491 w_3185628_870308# w_3185628_834308# sky130_fd_pr__diode_pd2nw_05v5 area=2.25e+16p
X492 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X493 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X494 w_3263498_541854# a_3405057_686207# a_3405057_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X495 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X496 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X497 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X498 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X499 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X500 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X501 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X502 a_3285528_930602# a_3361095_700871# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X503 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X504 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X505 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X506 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X507 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X508 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X509 a_3420294_717833# a_3381563_717833# w_3422394_717637# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X510 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X511 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X512 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X513 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X514 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X515 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X516 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X517 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X518 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X519 a_3383521_705357# a_3381660_702705# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=2.8e+06u
X520 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X521 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X522 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X523 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X524 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X525 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X526 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X527 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X528 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X529 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X530 a_3403286_704090# a_3403286_703346# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X531 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X532 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X533 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X534 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X535 w_3422394_717637# a_3381563_717833# a_3420294_717833# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X536 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X537 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X538 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X539 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X540 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X541 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X542 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X543 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X544 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X545 a_3443016_749796# a_3439418_744112# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X546 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X547 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X548 a_3420294_720809# a_3420381_704937# w_3422394_717637# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X549 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X550 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X551 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X552 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X553 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X554 a_3420294_717833# a_3420294_717833# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X555 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X556 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X557 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X558 w_3403067_716474# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X559 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X560 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X561 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X562 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X563 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X564 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X565 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X566 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X567 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X568 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X569 w_3185490_798160# a_3381660_718033# a_3381660_718033# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X570 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X571 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X572 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X573 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X574 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X575 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X576 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X577 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X578 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X579 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X580 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X581 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X582 a_3381660_718777# a_3381660_718033# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X583 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X584 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X585 w_3381441_717637# a_3381563_717833# a_3381660_718033# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X586 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X587 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X588 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X589 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X590 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X591 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X592 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X593 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X594 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X595 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X596 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X597 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X598 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X599 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X600 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X601 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X602 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X603 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X604 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X605 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X606 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X607 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X608 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X609 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X610 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X611 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X612 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X613 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X614 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X615 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X616 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X617 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X618 w_3185490_798160# a_3403286_716870# a_3403286_716870# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X619 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X620 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X621 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X622 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X623 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X624 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X625 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X626 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X627 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X628 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X629 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X630 w_3263498_541854# a_3407435_674425# w_3422393_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X631 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X632 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X633 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X634 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X635 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X636 w_3185490_798160# a_3434368_749958# a_3428294_754598# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X637 a_3394410_690671# a_3394410_687695# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X638 a_3407542_687895# a_3407282_686697# w_3407323_687499# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X639 a_3369760_754598# a_3366260_744206# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X640 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X641 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X642 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X643 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X644 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X645 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X646 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X647 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X648 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X649 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X650 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X651 w_3185490_798160# a_3403286_703346# a_3403286_704090# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X652 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X653 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X654 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X655 a_3367712_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X656 a_3420293_704737# a_3420293_701761# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X657 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X658 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X659 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X660 a_3381660_702705# a_3381660_701961# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X661 w_3185490_798160# a_3434368_749958# a_3428294_754598# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X662 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X663 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X664 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X665 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X666 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X667 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X668 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X669 w_3263498_541854# a_3379175_716345# a_3379175_716345# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X670 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X671 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X672 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X673 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X674 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X675 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X676 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X677 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X678 a_3379175_716345# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X679 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X680 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X681 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X682 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X683 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X684 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X685 w_3185490_798160# a_3439418_744112# a_3443016_749796# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X686 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X687 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X688 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X689 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X690 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X691 w_3263498_541854# a_3401256_686207# a_3401256_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X692 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X693 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X694 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X695 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X696 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X697 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X698 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X699 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X700 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X701 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X702 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X703 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X704 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X705 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X706 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X707 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X708 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X709 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X710 w_3263498_541854# a_3400801_701658# a_3400801_701658# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X711 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X712 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X713 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X714 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X715 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X716 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X717 w_3263498_541854# a_3400801_701658# a_3400801_701658# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X718 v2 a_3435992_747994# a_3434368_749958# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X719 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X720 a_3394410_687695# a_3394410_687695# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X721 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X722 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X723 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X724 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X725 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X726 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X727 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X728 w_3185490_798160# a_3399027_674337# a_3379175_716345# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X729 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X730 w_3422394_717637# a_3381563_717833# a_3420294_717833# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X731 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X732 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X733 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X734 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X735 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X736 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X737 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X738 a_3436064_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X739 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X740 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X741 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X742 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X743 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X744 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X745 a_3420294_720809# a_3420381_704937# w_3422394_717637# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X746 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X747 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X748 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X749 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X750 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X751 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X752 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X753 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X754 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X755 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X756 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X757 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X758 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X759 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X760 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X761 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X762 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X763 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X764 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X765 a_3408579_674425# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X766 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X767 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X768 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X769 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X770 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X771 a_3436064_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X772 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X773 a_3359810_749958# a_3362834_747994# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X774 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X775 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X776 a_3403286_703346# a_3403286_703346# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X777 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X778 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X779 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X780 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X781 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X782 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X783 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X784 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X785 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X786 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X787 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X788 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X789 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X790 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X791 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X792 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X793 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X794 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X795 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X796 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X797 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X798 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X799 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X800 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X801 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X802 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X803 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X804 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X805 a_3400801_715182# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X806 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X807 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X808 a_3403286_717614# a_3403189_717414# w_3403067_716474# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X809 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X810 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X811 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X812 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X813 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X814 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X815 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X816 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X817 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X818 a_3420293_701761# a_3420293_701761# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X819 v2 a_3439418_744112# a_3443016_749796# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X820 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X821 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X822 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X823 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X824 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X825 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X826 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X827 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X828 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X829 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X830 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X831 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X832 a_3440844_744112# a_3420382_721009# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X833 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X834 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X835 a_3428294_754598# a_3434368_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X836 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X837 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X838 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X839 w_3263498_541854# a_3401256_686207# w_3396510_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X840 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X841 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X842 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X843 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X844 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X845 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X846 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X847 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X848 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X849 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X850 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X851 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X852 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X853 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X854 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X855 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X856 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X857 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X858 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X859 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X860 a_3428294_754598# a_3434368_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X861 a_3366260_744206# a_3369760_747574# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X862 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X863 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X864 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X865 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X866 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X867 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X868 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X869 a_3367712_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X870 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X871 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X872 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X873 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X874 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X875 w_3263498_541854# a_3407435_674425# w_3422393_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X876 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X877 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X878 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X879 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X880 v2 a_3366260_744206# a_3369760_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X881 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X882 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X883 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X884 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X885 a_3403001_700774# a_3381563_717833# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X886 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X887 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X888 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X889 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X890 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X891 a_3381660_701961# a_3361095_699281# w_3381441_701565# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X892 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X893 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X894 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X895 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X896 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X897 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X898 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X899 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X900 a_3359663_699281# a_3361095_699599# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X901 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X902 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X903 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X904 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X905 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X906 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X907 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X908 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X909 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X910 w_3263498_541854# a_3379175_716345# a_3379175_716345# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X911 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X912 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X913 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X914 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X915 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X916 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X917 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X918 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X919 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X920 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X921 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X922 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X923 a_3379175_716345# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X924 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X925 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X926 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X927 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X928 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X929 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X930 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X931 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X932 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X933 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X934 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X935 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X936 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X937 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X938 w_3185490_798160# a_3399027_674337# a_3400801_701658# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X939 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X940 w_3263498_541854# a_3400801_701658# w_3403067_702950# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X941 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X942 w_3403067_702950# a_3403001_700774# a_3403286_703346# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X943 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X944 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X945 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X946 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X947 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X948 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X949 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X950 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X951 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X952 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X953 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
R2 v1 v2 sky130_fd_pr__res_generic_m5 w=7.42e+07u l=1.885e+07u
X954 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X955 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X956 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X957 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X958 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X959 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X960 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X961 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X962 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X963 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X964 a_3420293_701761# a_3422243_697443# w_3422393_701565# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X965 a_3440870_744142# a_3440844_744112# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X966 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X967 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X968 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X969 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X970 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X971 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X972 v2 a_3359810_749958# a_3335479_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X973 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X974 a_3400801_715182# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X975 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X976 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X977 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X978 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X979 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X980 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X981 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X982 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X983 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X984 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X985 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X986 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X987 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X988 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X989 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X990 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X991 a_3435992_747994# a_3436064_746854# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X992 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X993 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X994 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X995 a_3422243_697443# a_3420381_704937# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X996 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X997 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X998 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X999 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1000 w_3263498_541854# a_3401256_686207# a_3401256_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1001 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1002 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1003 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1004 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1005 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1006 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1007 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1008 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1009 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1010 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1011 w_3381441_717637# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1012 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1013 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1014 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1015 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1016 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1017 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1018 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1019 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1020 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1021 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1022 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1023 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1024 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1025 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1026 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1027 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1028 a_3403286_717614# a_3403189_717414# w_3403067_716474# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1029 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1030 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1031 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1032 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1033 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1034 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1035 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1036 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1037 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1038 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1039 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1040 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1041 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1042 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1043 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1044 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1045 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1046 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1047 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1048 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1049 a_3362906_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X1050 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1051 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1052 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1053 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1054 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1055 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1056 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1057 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1058 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1059 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1060 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1061 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1062 a_3421607_697443# a_3421289_698875# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X1063 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1064 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1065 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1066 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1067 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1068 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1069 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1070 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1071 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1072 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1073 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1074 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1075 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1076 a_3361095_699281# a_3379272_706425# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X1077 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1078 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1079 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1080 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1081 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1082 a_3420293_704737# a_3381563_702505# w_3422393_701565# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1083 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1084 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1085 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1086 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1087 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1088 w_3263498_541854# a_3408579_674425# a_3408579_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1089 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1090 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1091 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1092 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1093 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1094 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1095 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1096 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1097 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1098 w_3407323_687499# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1099 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1100 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1101 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1102 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1103 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1104 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1105 w_3185490_798160# a_3420294_717833# a_3420294_720809# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1106 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1107 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1108 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1109 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1110 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1111 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1112 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1113 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1114 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1115 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1116 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1117 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1118 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1119 a_3403286_716870# a_3381563_702505# w_3403067_716474# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1120 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1121 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1122 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1123 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1124 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1125 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1126 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1127 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1128 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1129 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1130 a_3420293_701761# a_3422243_697443# w_3422393_701565# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1131 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1132 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1133 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1134 v2 a_3439418_744112# a_3443016_749796# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1135 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1136 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1137 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1138 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1139 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1140 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1141 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1142 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1143 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1144 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1145 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1146 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1147 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1148 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1149 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1150 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1151 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1152 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1153 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1154 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1155 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1156 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1157 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1158 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1159 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1160 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1161 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1162 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1163 w_3185490_798160# a_3403286_703346# a_3403286_704090# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1164 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1165 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1166 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1167 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1168 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1169 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1170 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1171 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1172 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1173 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1174 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1175 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1176 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1177 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1178 a_3394410_687695# a_3394410_687695# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1179 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1180 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1181 w_3263498_541854# a_3379175_700273# w_3381441_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1182 a_3408579_674425# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1183 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1184 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1185 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1186 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1187 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1188 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1189 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1190 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1191 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1192 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1193 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1194 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1195 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1196 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1197 a_3359810_749958# a_3362834_747994# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1198 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1199 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1200 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1201 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1202 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1203 a_3434368_749958# a_3435992_747994# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1204 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1205 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1206 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1207 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1208 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1209 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1210 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1211 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1212 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1213 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1214 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1215 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1216 w_3381441_717637# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1217 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1218 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1219 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1220 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1221 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1222 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1223 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1224 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1225 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1226 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1227 w_3685938_653428# w_3685938_617428# sky130_fd_pr__diode_pd2nw_05v5 area=2.25e+16p
X1228 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1229 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1230 w_3403067_716474# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1231 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1232 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1233 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1234 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1235 v2 a_3434368_749958# a_3428294_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1236 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1237 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1238 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1239 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1240 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1241 a_3420294_720809# a_3420294_717833# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1242 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1243 a_3407542_688639# a_3381563_702505# w_3407323_687499# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1244 a_3381660_701961# a_3381660_701961# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1245 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1246 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1247 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1248 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1249 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X1250 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1251 w_3263498_541854# a_3405057_686207# w_3407323_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1252 w_3185490_798160# a_3407542_687895# a_3407542_687895# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1253 a_3422243_697443# a_3420381_704937# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X1254 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1255 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1256 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1257 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1258 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1259 a_3403001_699542# a_3403001_700774# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X1260 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1261 a_3443016_749796# a_3439418_744112# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1262 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1263 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1264 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1265 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1266 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1267 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1268 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1269 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1270 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1271 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1272 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1273 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1274 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1275 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1276 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1277 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1278 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1279 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1280 a_3369760_754598# a_3366260_744206# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1281 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1282 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1283 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1284 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1285 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1286 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X1287 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1288 a_3335479_772599# a_3359810_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1289 a_3361095_699281# a_3379272_706425# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X1290 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1291 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1292 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1293 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1294 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1295 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1296 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1297 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1298 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1299 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1300 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1301 a_3420293_704737# a_3381563_702505# w_3422393_701565# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1302 a_3403286_716870# a_3381563_702505# w_3403067_716474# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1303 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1304 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1305 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1306 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1307 a_3367712_744142# a_3359810_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1308 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1309 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1310 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1311 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1312 a_3394410_690671# a_3394410_687695# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1313 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1314 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1315 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1316 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1317 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1318 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1319 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1320 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1321 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1322 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1323 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1324 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1325 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1326 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1327 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1328 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1329 a_3403286_716870# a_3381563_702505# w_3403067_716474# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1330 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1331 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1332 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1333 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1334 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1335 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1336 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1337 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1338 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1339 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1340 a_3335479_772599# a_3359810_749958# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1341 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1342 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1343 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1344 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1345 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1346 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1347 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1348 a_3407542_688639# a_3407542_687895# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1349 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1350 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1351 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1352 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1353 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1354 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1355 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1356 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1357 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1358 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1359 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1360 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1361 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1362 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1363 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1364 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1365 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1366 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1367 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1368 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1369 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1370 a_3369760_754598# a_3366260_744206# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1371 a_3335479_772599# a_3359810_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1372 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1373 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1374 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1375 a_3428294_754598# a_3434368_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1376 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1377 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1378 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1379 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1380 w_3185490_798160# a_3439418_744112# a_3443016_749796# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1381 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1382 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1383 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1384 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1385 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1386 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1387 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1388 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1389 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1390 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1391 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1392 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1393 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1394 w_3263498_541854# a_3400801_701658# a_3400801_701658# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1395 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1396 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X1397 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1398 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1399 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1400 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1401 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1402 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1403 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1404 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1405 w_3263498_541854# a_3408579_674425# w_3422394_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1406 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1407 a_3440870_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X1408 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1409 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1410 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1411 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1412 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1413 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1414 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1415 a_3420294_720809# a_3420381_704937# w_3422394_717637# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1416 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1417 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1418 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1419 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1420 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1421 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1422 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1423 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1424 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1425 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1426 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1427 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1428 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1429 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1430 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1431 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1432 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1433 a_3440870_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X1434 v2 a_3442918_747574# a_3439418_744112# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1435 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1436 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1437 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1438 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1439 a_3381660_718777# a_3381660_718033# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1440 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1441 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1442 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1443 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1444 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1445 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1446 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1447 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1448 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1449 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1450 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1451 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1452 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1453 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1454 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1455 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1456 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1457 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1458 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1459 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1460 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1461 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1462 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1463 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1464 w_3185490_798160# a_3366260_744206# a_3369760_754598# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1465 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1466 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1467 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1468 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1469 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1470 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1471 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1472 a_3400801_715182# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1473 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1474 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1475 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1476 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1477 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1478 w_3263498_541854# a_3400801_701658# w_3403067_702950# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1479 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1480 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1481 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1482 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1483 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1484 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1485 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1486 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1487 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1488 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1489 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1490 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X1491 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1492 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1493 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1494 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1495 a_3428294_754598# a_3434368_749958# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1496 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1497 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1498 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1499 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1500 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1501 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1502 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1503 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1504 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1505 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1506 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1507 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1508 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1509 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1510 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1511 a_3443016_749796# a_3439418_744112# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1512 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1513 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1514 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1515 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1516 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1517 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1518 a_3367712_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X1519 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1520 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1521 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1522 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1523 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1524 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1525 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1526 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1527 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1528 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1529 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1530 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1531 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1532 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1533 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1534 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1535 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1536 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1537 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1538 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1539 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1540 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1541 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1542 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1543 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1544 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1545 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1546 a_3367712_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X1547 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1548 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1549 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1550 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1551 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1552 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1553 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1554 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1555 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1556 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1557 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1558 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1559 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1560 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1561 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1562 w_3185490_798160# a_3407542_687895# a_3407542_688639# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1563 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1564 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1565 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1566 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1567 w_3263498_541854# a_3379175_716345# a_3379175_716345# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1568 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1569 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1570 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1571 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1572 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1573 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1574 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1575 v2 a_3362834_747994# a_3359810_749958# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1576 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1577 a_3420294_720809# a_3420381_704937# w_3422394_717637# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1578 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1579 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1580 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1581 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1582 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1583 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1584 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1585 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1586 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1587 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1588 w_3263498_541854# a_3401256_686207# w_3396510_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1589 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1590 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1591 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1592 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1593 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1594 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1595 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1596 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1597 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1598 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1599 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1600 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1601 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1602 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1603 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1604 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1605 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1606 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1607 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1608 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1609 v2 a_3436064_746854# a_3435992_747994# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1610 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1611 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1612 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1613 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1614 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1615 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1616 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1617 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1618 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1619 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1620 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1621 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1622 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1623 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1624 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1625 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1626 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1627 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1628 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1629 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1630 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1631 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1632 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X1633 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1634 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1635 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1636 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1637 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1638 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1639 v2 a_3434368_749958# a_3428294_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1640 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1641 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1642 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1643 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1644 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1645 w_3263498_541854# a_3379175_700273# w_3381441_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1646 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1647 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1648 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1649 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1650 a_3381660_701961# a_3361095_699281# w_3381441_701565# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1651 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1652 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1653 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1654 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1655 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1656 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1657 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1658 a_3404273_699542# a_3403955_700774# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X1659 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1660 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1661 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1662 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1663 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1664 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1665 a_3420294_717833# a_3420294_717833# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1666 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1667 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1668 v2 a_3434368_749958# a_3428294_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1669 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1670 v2 a_3369760_747574# a_3366260_744206# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1671 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X1672 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1673 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1674 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1675 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1676 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1677 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1678 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1679 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1680 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1681 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1682 w_3396510_687499# a_3387775_698875# a_3394410_687695# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1683 a_3409645_692829# a_3405154_692359# sky130_fd_pr__cap_mim_m3_1 l=1.4e+07u w=1.4e+07u
X1684 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1685 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1686 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1687 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1688 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1689 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1690 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1691 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1692 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1693 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1694 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1695 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1696 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1697 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1698 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1699 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1700 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1701 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1702 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1703 w_3263498_541854# a_3407435_674425# w_3422393_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1704 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1705 a_3381660_718033# a_3381660_718033# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1706 a_3386185_697443# a_3386503_698875# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X1707 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1708 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1709 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1710 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1711 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1712 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1713 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1714 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1715 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1716 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1717 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1718 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1719 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1720 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1721 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1722 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1723 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1724 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1725 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1726 a_3399027_674337# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X1727 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1728 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1729 a_3394410_690671# a_3394410_687695# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1730 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1731 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1732 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1733 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1734 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1735 w_3263498_541854# a_3401256_686207# w_3396510_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1736 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1737 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1738 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1739 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1740 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1741 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1742 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1743 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1744 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1745 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1746 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1747 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1748 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1749 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1750 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1751 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1752 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1753 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1754 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1755 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1756 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1757 w_3185490_798160# a_3381660_701961# a_3381660_702705# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1758 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1759 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1760 w_3185490_798160# a_3399027_674337# a_3379175_700273# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X1761 a_3381660_702705# a_3381563_702505# w_3381441_701565# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1762 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1763 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1764 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1765 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1766 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1767 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1768 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1769 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1770 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1771 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1772 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X1773 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1774 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1775 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1776 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1777 w_3185490_798160# a_3399027_674337# a_3400801_715182# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X1778 w_3263498_541854# a_3400801_701658# a_3400801_701658# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1779 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1780 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1781 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1782 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1783 a_3407542_687895# a_3407282_686697# w_3407323_687499# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1784 a_3420293_704737# a_3420293_701761# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1785 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1786 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1787 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1788 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1789 w_3263498_541854# a_3405057_686207# w_3407323_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1790 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1791 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1792 w_3185490_798160# a_3407542_687895# a_3407542_688639# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1793 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1794 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1795 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1796 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1797 a_3381660_718033# a_3381563_717833# w_3381441_717637# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1798 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1799 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1800 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1801 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1802 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1803 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1804 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1805 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1806 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1807 a_3403286_716870# a_3403286_716870# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1808 w_3263498_541854# a_3379175_716345# w_3381441_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1809 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1810 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1811 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1812 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1813 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1814 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1815 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1816 a_3403286_704090# a_3403286_703346# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1817 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1818 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1819 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1820 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1821 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1822 a_3379175_700273# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X1823 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1824 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1825 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1826 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1827 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1828 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1829 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1830 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1831 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1832 w_3263498_541854# a_3401256_686207# a_3401256_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1833 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1834 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1835 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1836 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1837 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1838 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1839 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1840 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1841 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1842 w_3263498_541854# a_3400801_715182# w_3403067_716474# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1843 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1844 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1845 v2 a_3442918_747574# a_3439418_744112# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1846 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1847 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1848 a_3381660_718033# a_3381660_718033# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1849 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1850 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1851 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1852 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1853 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1854 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1855 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1856 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1857 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1858 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1859 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1860 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1861 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1862 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1863 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1864 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1865 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1866 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1867 w_3407323_687499# a_3407282_686697# a_3407542_687895# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1868 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1869 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1870 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1871 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1872 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1873 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1874 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1875 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1876 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1877 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1878 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1879 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1880 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1881 a_3407542_687895# a_3407542_687895# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1882 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1883 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1884 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1885 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1886 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1887 w_3263498_541854# a_3379175_700273# w_3381441_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1888 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1889 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1890 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1891 a_3420335_697443# a_3405154_692359# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X1892 a_3420294_717833# a_3381563_717833# w_3422394_717637# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1893 a_3404909_699542# a_3404591_700774# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X1894 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1895 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1896 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1897 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1898 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1899 w_3185490_798160# a_3420293_701761# a_3420293_704737# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1900 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1901 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1902 a_3443016_749796# a_3439418_744112# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1903 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1904 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1905 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1906 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1907 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1908 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1909 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1910 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1911 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1912 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1913 w_3422393_701565# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1914 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1915 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1916 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1917 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1918 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1919 w_3185490_798160# a_3381660_718033# a_3381660_718033# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1920 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1921 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1922 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1923 w_3407323_687499# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1924 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1925 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1926 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1927 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1928 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1929 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1930 w_3263498_541854# a_3408579_674425# w_3422394_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1931 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1932 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1933 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1934 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1935 a_3381660_718777# a_3381660_718033# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1936 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1937 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1938 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1939 w_3422394_717637# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1940 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1941 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1942 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1943 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1944 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1945 a_3405057_686207# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1946 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1947 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1948 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1949 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1950 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1951 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1952 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1953 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1954 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1955 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1956 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1957 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1958 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X1959 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1960 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1961 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1962 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1963 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1964 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1965 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1966 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1967 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1968 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1969 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1970 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1971 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1972 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1973 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1974 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1975 a_3361095_699281# a_3379272_706425# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X1976 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1977 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1978 v2 w_3185628_906308# sky130_fd_pr__diode_pd2nw_05v5 area=2.25e+16p
X1979 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1980 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1981 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1982 w_3396510_687499# a_3263636_541992# a_3394410_690671# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1983 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1984 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1985 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1986 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1987 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1988 a_3381660_702705# a_3381563_702505# w_3381441_701565# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1989 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1990 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1991 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1992 a_3400801_715182# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1993 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1994 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1995 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1996 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1997 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1998 a_3422243_697443# a_3420381_704937# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X1999 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2000 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2001 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2002 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2003 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2004 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2005 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2006 a_3420293_704737# a_3420293_701761# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2007 w_3403067_702950# a_3381563_702505# a_3403286_704090# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2008 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2009 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2010 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2011 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2012 w_3263498_541854# a_3400801_701658# w_3403067_702950# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2013 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2014 w_3381441_717637# a_3381563_717833# a_3381660_718033# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2015 a_3442918_747574# a_3440870_744142# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2016 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2017 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2018 w_3185490_798160# a_3399027_674337# a_3408579_674425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X2019 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2020 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2021 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2022 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2023 a_3440870_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X2024 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2025 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2026 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2027 a_3381660_718777# a_3379272_706425# w_3381441_717637# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2028 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2029 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2030 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2031 a_3367712_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X2032 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2033 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2034 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2035 w_3185490_798160# a_3420294_717833# a_3420294_720809# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2036 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2037 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2038 w_3185490_798160# a_3435992_747994# a_3434368_749958# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2039 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2040 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2041 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2042 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2043 a_3401256_686207# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2044 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2045 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2046 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2047 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2048 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2049 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2050 a_3361095_699281# a_3379272_706425# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X2051 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2052 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2053 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2054 a_3440870_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X2055 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2056 a_3405057_686207# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X2057 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2058 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2059 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2060 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2061 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2062 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2063 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2064 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2065 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2066 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2067 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2068 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2069 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2070 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2071 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2072 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2073 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2074 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2075 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2076 a_3434368_749958# a_3435992_747994# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2077 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2078 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2079 w_3263498_541854# a_3400801_715182# w_3403067_716474# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2080 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2081 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2082 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2083 w_3185490_798160# a_3381660_701961# a_3381660_701961# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2084 w_3263498_541854# a_3407435_674425# w_3422393_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2085 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2086 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2087 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2088 v2 a_3439418_744112# a_3443016_749796# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2089 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2090 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2091 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2092 a_3387457_697443# a_3387775_698875# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X2093 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2094 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2095 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2096 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2097 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2098 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2099 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2100 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2101 v2 a_3366260_744206# a_3369760_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2102 a_3400898_721334# a_3403189_717414# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=9e+06u
X2103 w_3263498_541854# a_3379175_716345# a_3379175_716345# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2104 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2105 v2 a_3359810_749958# a_3335479_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2106 a_3408579_674425# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X2107 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2108 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2109 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2110 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2111 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2112 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2113 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2114 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2115 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2116 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2117 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2118 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2119 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2120 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2121 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2122 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2123 w_3381441_717637# a_3379272_706425# a_3381660_718777# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2124 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2125 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2126 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2127 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2128 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2129 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2130 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2131 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2132 a_3367712_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X2133 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2134 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2135 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2136 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2137 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2138 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2139 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2140 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2141 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2142 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2143 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2144 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2145 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2146 w_3185490_798160# a_3359810_749958# a_3335479_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2147 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2148 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2149 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2150 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2151 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2152 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2153 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2154 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2155 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2156 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2157 w_3407323_687499# a_3381563_702505# a_3407542_688639# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2158 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2159 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2160 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2161 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2162 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2163 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2164 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2165 w_3407323_687499# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2166 a_3367712_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X2167 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2168 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2169 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2170 w_3263498_541854# a_3379175_700273# w_3381441_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2171 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2172 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2173 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2174 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2175 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2176 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2177 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2178 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2179 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2180 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2181 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2182 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2183 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2184 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2185 v2 a_3366260_744206# a_3369760_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2186 v2 a_3359810_749958# a_3335479_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2187 v2 a_3434368_749958# a_3428294_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2188 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2189 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2190 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2191 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2192 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2193 w_3185490_798160# a_3420294_717833# a_3420294_720809# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2194 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2195 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2196 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2197 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2198 w_3185490_798160# a_3420293_701761# a_3420293_701761# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2199 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2200 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2201 w_3396510_687499# a_3263636_541992# a_3394410_690671# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2202 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2203 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2204 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2205 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2206 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2207 a_3440870_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X2208 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2209 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2210 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2211 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2212 w_3381441_701565# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2213 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2214 w_3403067_716474# a_3403189_717414# a_3403286_717614# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2215 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2216 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2217 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2218 a_3422243_697443# a_3420381_704937# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X2219 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2220 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2221 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2222 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2223 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2224 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2225 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2226 w_3263498_541854# a_3400801_701658# w_3403067_702950# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2227 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2228 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2229 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2230 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2231 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2232 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2233 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2234 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2235 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2236 a_3335479_772599# a_3359810_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2237 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2238 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2239 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2240 a_3439418_744112# a_3442918_747574# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2241 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2242 a_3440870_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X2243 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2244 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2245 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2246 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2247 a_3369760_754598# a_3366260_744206# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2248 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2249 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2250 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2251 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2252 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2253 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2254 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2255 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2256 a_3394410_687695# a_3394410_687695# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2257 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2258 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2259 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2260 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2261 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2262 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2263 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2264 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2265 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2266 w_3263498_541854# a_3401256_686207# w_3396510_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2267 a_3335479_772599# a_3359810_749958# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2268 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2269 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2270 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2271 a_3369760_754598# a_3366260_744206# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2272 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2273 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X2274 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2275 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2276 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2277 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2278 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2279 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2280 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2281 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2282 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2283 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2284 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2285 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2286 a_3407282_686697# a_3408714_686379# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X2287 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2288 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2289 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2290 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2291 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2292 a_3403286_716870# a_3403286_716870# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2293 a_3362906_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X2294 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2295 w_3403067_716474# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2296 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2297 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2298 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2299 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2300 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2301 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2302 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2303 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2304 a_3369760_754598# a_3366260_744206# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2305 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2306 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2307 a_3379175_716345# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2308 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2309 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2310 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2311 w_3185490_798160# a_3439418_744112# a_3443016_749796# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2312 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2313 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2314 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2315 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2316 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2317 w_3263498_541854# a_3379175_716345# w_3381441_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2318 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2319 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2320 a_3367712_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X2321 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2322 w_3403067_702950# a_3381563_702505# a_3403286_704090# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2323 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2324 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2325 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2326 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2327 w_3185490_798160# a_3420294_717833# a_3420294_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2328 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2329 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2330 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2331 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2332 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2333 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2334 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2335 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2336 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2337 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2338 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2339 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2340 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2341 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2342 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2343 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2344 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2345 a_3367712_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X2346 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2347 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2348 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2349 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2350 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2351 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2352 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2353 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2354 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2355 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2356 a_3394410_690671# a_3263636_541992# w_3396510_687499# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2357 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2358 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2359 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2360 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2361 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2362 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2363 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2364 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2365 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X2366 w_3185490_798160# a_3381660_718033# a_3381660_718777# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2367 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2368 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2369 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2370 w_3407323_687499# a_3381563_702505# a_3407542_688639# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2371 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2372 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2373 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2374 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2375 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2376 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2377 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2378 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2379 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2380 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2381 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2382 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2383 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2384 w_3263498_541854# a_3379175_700273# a_3379175_700273# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2385 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2386 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2387 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2388 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2389 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2390 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2391 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2392 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2393 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2394 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2395 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2396 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2397 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2398 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2399 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2400 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2401 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2402 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2403 w_3263498_541854# a_3379175_700273# w_3381441_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2404 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2405 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2406 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2407 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2408 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2409 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2410 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2411 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2412 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2413 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2414 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2415 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2416 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2417 a_3405389_721804# a_3400898_721334# sky130_fd_pr__cap_mim_m3_1 l=1.4e+07u w=1.4e+07u
X2418 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2419 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2420 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2421 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2422 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2423 w_3422394_717637# a_3420381_704937# a_3420294_720809# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2424 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2425 w_3263498_541854# a_3401256_686207# w_3396510_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2426 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2427 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2428 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2429 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2430 w_3381441_717637# a_3381563_717833# a_3381660_718033# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2431 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2432 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2433 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2434 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2435 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2436 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2437 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2438 w_3422393_701565# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2439 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2440 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2441 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2442 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2443 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2444 w_3263498_541854# a_3400801_701658# a_3400801_701658# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2445 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2446 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2447 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2448 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2449 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2450 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2451 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2452 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2453 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X2454 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2455 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2456 a_3407542_687895# a_3407282_686697# w_3407323_687499# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2457 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2458 a_3405057_686207# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2459 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2460 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2461 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2462 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2463 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2464 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2465 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2466 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2467 a_3436064_746854# a_3420382_721009# a_3439444_744142# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2468 v2 a_3362906_746854# a_3362834_747994# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2469 a_3428294_754598# a_3434368_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2470 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2471 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2472 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2473 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2474 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2475 a_3443016_749796# a_3439418_744112# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2476 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2477 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2478 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2479 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2480 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2481 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2482 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2483 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2484 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2485 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2486 a_3403001_700774# a_3381563_717833# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X2487 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2488 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2489 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2490 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2491 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2492 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2493 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2494 a_3424227_705357# a_3420381_704937# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=1.4e+07u
X2495 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2496 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2497 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2498 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2499 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2500 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2501 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2502 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2503 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2504 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2505 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2506 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2507 w_3403067_702950# a_3381563_702505# a_3403286_704090# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2508 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2509 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2510 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2511 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2512 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2513 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2514 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2515 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2516 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2517 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2518 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2519 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2520 w_3403067_716474# a_3381563_702505# a_3403286_716870# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2521 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2522 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2523 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2524 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2525 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2526 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2527 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2528 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2529 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2530 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2531 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2532 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2533 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2534 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2535 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2536 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2537 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2538 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2539 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2540 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2541 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2542 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2543 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2544 a_3394410_687695# a_3394410_687695# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2545 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2546 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2547 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2548 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2549 w_3185490_798160# a_3362834_747994# a_3359810_749958# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2550 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2551 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2552 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2553 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2554 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X2555 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2556 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2557 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2558 v2 a_3367712_744142# a_3369760_747574# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2559 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2560 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2561 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2562 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2563 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2564 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2565 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2566 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2567 a_3401256_686207# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2568 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2569 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2570 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2571 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2572 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2573 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2574 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2575 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2576 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2577 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2578 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2579 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2580 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2581 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2582 w_3422394_717637# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2583 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2584 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2585 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2586 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2587 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2588 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2589 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2590 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2591 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2592 a_3428294_754598# a_3434368_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2593 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2594 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2595 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2596 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2597 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2598 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2599 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2600 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2601 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2602 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2603 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2604 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2605 w_3185490_798160# a_3381660_701961# a_3381660_702705# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2606 w_3263498_541854# a_3407435_674425# w_3422393_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2607 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2608 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2609 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2610 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2611 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2612 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2613 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2614 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2615 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2616 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2617 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2618 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2619 a_3401256_686207# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X2620 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2621 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2622 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2623 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2624 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2625 w_3263498_541854# a_3379175_700273# a_3379175_700273# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2626 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2627 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2628 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2629 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2630 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2631 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2632 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2633 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2634 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2635 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2636 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2637 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2638 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2639 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2640 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2641 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2642 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2643 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2644 w_3263498_541854# a_3401256_686207# a_3401256_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2645 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2646 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2647 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2648 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2649 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2650 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2651 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2652 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2653 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2654 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2655 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2656 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2657 a_3407435_674425# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2658 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2659 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2660 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2661 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2662 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2663 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2664 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2665 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2666 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2667 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2668 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2669 a_3403286_703346# a_3403001_700774# w_3403067_702950# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2670 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2671 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2672 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2673 w_3263498_541854# a_3405057_686207# w_3407323_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2674 w_3407323_687499# a_3407282_686697# a_3407542_687895# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2675 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2676 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2677 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2678 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2679 a_3403001_700774# a_3381563_717833# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X2680 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2681 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2682 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2683 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2684 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2685 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2686 w_3407323_687499# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2687 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2688 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2689 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2690 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2691 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2692 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2693 a_3403286_717614# a_3403286_716870# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2694 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2695 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2696 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2697 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2698 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2699 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2700 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2701 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2702 v2 a_3439418_744112# a_3443016_749796# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2703 a_3428294_754598# a_3434368_749958# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2704 a_3403637_699542# a_3403319_700774# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X2705 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2706 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2707 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2708 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2709 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2710 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2711 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2712 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2713 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2714 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2715 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2716 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2717 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2718 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2719 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2720 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2721 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2722 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2723 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2724 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2725 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2726 a_3443016_749796# a_3439418_744112# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2727 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2728 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2729 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2730 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2731 w_3185490_798160# a_3420293_701761# a_3420293_704737# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2732 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2733 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2734 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2735 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2736 w_3422393_701565# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2737 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2738 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2739 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2740 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2741 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2742 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2743 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2744 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2745 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2746 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2747 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2748 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2749 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2750 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2751 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2752 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2753 w_3381441_701565# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2754 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2755 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2756 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2757 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2758 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2759 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2760 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2761 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2762 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2763 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2764 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2765 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2766 w_3185490_798160# a_3394410_687695# a_3394410_687695# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2767 a_3405057_686207# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2768 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2769 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2770 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2771 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2772 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2773 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2774 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2775 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2776 a_3381660_718777# a_3381660_718033# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2777 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2778 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2779 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2780 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2781 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2782 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2783 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2784 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2785 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2786 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2787 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2788 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2789 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2790 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2791 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2792 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2793 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2794 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2795 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2796 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2797 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2798 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2799 a_3420293_701761# a_3420293_701761# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2800 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2801 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2802 a_3381660_701961# a_3381660_701961# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2803 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2804 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2805 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2806 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2807 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2808 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2809 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2810 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2811 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2812 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2813 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2814 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2815 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2816 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2817 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2818 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2819 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2820 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2821 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2822 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2823 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2824 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2825 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2826 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2827 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2828 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2829 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2830 w_3422394_717637# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2831 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2832 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2833 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2834 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2835 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2836 w_3185490_798160# a_3381660_701961# a_3381660_701961# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2837 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2838 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2839 w_3263498_541854# a_3407435_674425# a_3407435_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2840 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2841 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2842 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2843 w_3403067_716474# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2844 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2845 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2846 a_3443016_749796# a_3439418_744112# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2847 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2848 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2849 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2850 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2851 w_3185490_798160# a_3434368_749958# a_3428294_754598# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2852 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2853 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2854 w_3185490_798160# a_3403286_703346# a_3403286_703346# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2855 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2856 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2857 a_3379175_716345# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2858 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2859 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2860 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2861 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2862 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2863 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2864 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2865 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2866 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2867 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2868 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2869 a_3381660_718777# a_3379272_706425# w_3381441_717637# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2870 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2871 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2872 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2873 a_3440870_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X2874 w_3403067_702950# a_3403001_700774# a_3403286_703346# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2875 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2876 a_3401256_686207# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2877 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2878 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2879 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2880 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2881 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2882 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2883 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2884 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2885 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2886 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2887 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2888 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2889 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2890 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2891 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2892 a_3407542_688639# a_3407542_687895# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2893 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X2894 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2895 w_3396510_687499# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2896 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2897 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2898 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2899 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2900 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2901 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2902 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2903 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2904 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2905 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2906 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2907 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2908 a_3369760_754598# a_3366260_744206# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2909 w_3263498_541854# a_3400801_715182# w_3403067_716474# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2910 w_3263498_541854# a_3401256_686207# a_3401256_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2911 a_3440870_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X2912 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2913 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2914 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2915 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2916 a_3403286_704090# a_3403286_703346# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2917 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2918 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2919 a_3394410_687695# a_3387775_698875# w_3396510_687499# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2920 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2921 w_3263498_541854# a_3400801_715182# w_3403067_716474# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2922 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2923 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2924 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2925 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2926 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2927 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2928 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2929 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2930 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2931 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2932 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2933 w_3185490_798160# a_3399027_674337# a_3405057_686207# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X2934 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2935 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2936 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2937 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2938 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2939 a_3369760_754598# a_3366260_744206# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2940 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2941 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2942 a_3403286_717614# a_3403286_716870# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2943 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2944 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2945 w_3263498_541854# a_3379175_700273# a_3379175_700273# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2946 a_3362906_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X2947 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2948 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2949 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2950 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2951 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2952 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2953 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2954 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X2955 a_3359810_749958# a_3362834_747994# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2956 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2957 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2958 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2959 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2960 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2961 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2962 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2963 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2964 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2965 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2966 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2967 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2968 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2969 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2970 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2971 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2972 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2973 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2974 w_3185490_798160# a_3420293_701761# a_3420293_701761# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2975 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2976 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2977 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2978 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2979 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2980 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2981 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2982 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2983 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2984 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2985 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2986 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2987 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2988 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2989 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2990 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2991 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2992 a_3422243_697443# a_3420381_704937# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X2993 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2994 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2995 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2996 a_3379175_700273# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2997 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2998 a_3335479_772599# a_3359810_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2999 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3000 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3001 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3002 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3003 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3004 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3005 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3006 w_3263498_541854# a_3400801_701658# a_3400801_701658# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3007 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3008 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3009 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3010 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3011 w_3407323_687499# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3012 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3013 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3014 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3015 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3016 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3017 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3018 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3019 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3020 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3021 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3022 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3023 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3024 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3025 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3026 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3027 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3028 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3029 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3030 a_3394410_687695# a_3394410_687695# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3031 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3032 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3033 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3034 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3035 a_3335479_772599# a_3359810_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3036 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3037 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3038 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3039 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3040 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3041 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3042 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3043 a_3367712_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X3044 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3045 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3046 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3047 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3048 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3049 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3050 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3051 w_3185490_798160# a_3403286_703346# a_3403286_704090# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3052 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3053 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3054 a_3366260_744206# a_3369760_747574# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3055 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3056 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3057 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3058 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3059 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3060 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3061 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3062 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3063 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3064 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3065 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3066 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3067 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3068 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3069 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3070 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3071 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3072 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3073 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3074 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3075 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3076 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3077 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3078 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3079 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3080 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3081 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3082 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3083 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3084 w_3403067_702950# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3085 w_3403067_702950# a_3403001_700774# a_3403286_703346# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3086 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3087 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3088 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3089 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3090 v2 a_3359810_749958# a_3335479_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3091 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3092 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3093 w_3685938_581428# w_3185490_798160# sky130_fd_pr__diode_pd2nw_05v5 area=2.25e+16p
X3094 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3095 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3096 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3097 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3098 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3099 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3100 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3101 v2 a_3442918_747574# a_3439418_744112# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3102 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3103 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3104 w_3403067_716474# a_3403189_717414# a_3403286_717614# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3105 a_3400801_715182# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3106 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X3107 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3108 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3109 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3110 w_3263498_541854# a_3400801_701658# w_3403067_702950# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3111 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3112 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3113 w_3185490_798160# a_3366260_744206# a_3369760_754598# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3114 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3115 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3116 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3117 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3118 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3119 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3120 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3121 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3122 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3123 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3124 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3125 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3126 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3127 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3128 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3129 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3130 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3131 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3132 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3133 w_3185490_798160# a_3359810_749958# a_3335479_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3134 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3135 w_3185490_798160# a_3427310_772647# sky130_fd_pr__diode_pw2nd_05v5 area=2.25e+16p
X3136 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3137 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3138 w_3185490_798160# a_3366260_744206# a_3369760_754598# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3139 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3140 a_3420293_704737# a_3381563_702505# w_3422393_701565# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3141 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3142 w_3185490_798160# a_3381660_701961# a_3381660_702705# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3143 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3144 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3145 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3146 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3147 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3148 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3149 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3150 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3151 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3152 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3153 w_3403067_716474# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3154 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3155 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3156 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3157 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3158 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3159 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3160 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3161 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3162 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3163 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3164 w_3263498_541854# a_3400801_715182# a_3400801_715182# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3165 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3166 a_3362906_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X3167 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3168 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3169 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3170 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3171 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3172 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3173 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3174 v2 a_3366260_744206# a_3369760_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3175 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3176 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3177 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3178 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3179 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3180 w_3263498_541854# a_3400801_715182# w_3403067_716474# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3181 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3182 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3183 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3184 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3185 a_3362834_747994# a_3362906_746854# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3186 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3187 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3188 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3189 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3190 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3191 a_3403286_716870# a_3381563_702505# w_3403067_716474# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3192 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3193 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3194 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3195 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3196 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3197 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3198 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3199 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3200 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3201 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3202 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3203 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3204 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3205 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3206 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3207 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3208 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3209 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3210 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3211 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3212 w_3263498_541854# a_3379175_700273# a_3379175_700273# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3213 a_3381660_718033# a_3381563_717833# w_3381441_717637# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3214 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3215 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3216 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3217 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3218 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3219 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3220 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3221 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3222 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3223 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3224 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3225 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3226 w_3263498_541854# a_3379175_716345# a_3379175_716345# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3227 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3228 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3229 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3230 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3231 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3232 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3233 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3234 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3235 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3236 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3237 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3238 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3239 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3240 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3241 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3242 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3243 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3244 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3245 w_3381441_701565# a_3381563_702505# a_3381660_702705# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3246 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3247 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3248 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3249 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3250 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3251 a_3407435_674425# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3252 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3253 a_3403286_704090# a_3381563_702505# w_3403067_702950# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3254 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3255 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3256 w_3263498_541854# a_3400801_701658# w_3403067_702950# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3257 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3258 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3259 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3260 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3261 w_3185490_798160# a_3394410_687695# a_3394410_687695# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3262 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3263 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3264 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3265 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3266 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3267 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3268 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3269 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3270 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3271 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3272 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3273 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3274 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3275 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3276 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3277 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3278 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3279 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3280 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3281 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3282 a_3403286_716870# a_3403286_716870# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3283 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3284 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3285 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3286 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3287 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3288 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3289 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3290 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3291 a_3381660_718033# a_3381660_718033# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3292 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3293 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3294 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3295 a_3379175_716345# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X3296 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3297 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3298 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3299 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3300 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3301 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3302 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3303 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3304 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3305 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3306 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3307 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3308 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3309 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3310 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3311 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3312 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3313 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3314 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3315 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3316 w_3422393_701565# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3317 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3318 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3319 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3320 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3321 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3322 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3323 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3324 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3325 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3326 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3327 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3328 w_3403067_716474# a_3381563_702505# a_3403286_716870# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3329 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3330 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3331 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3332 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3333 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3334 a_3405057_686207# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3335 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3336 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3337 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3338 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3339 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3340 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3341 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3342 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3343 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3344 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3345 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3346 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3347 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3348 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3349 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3350 v2 a_3439418_744112# a_3443016_749796# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3351 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3352 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3353 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3354 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3355 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3356 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3357 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3358 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3359 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3360 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3361 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3362 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3363 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3364 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3365 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3366 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3367 a_3420293_704737# a_3381563_702505# w_3422393_701565# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3368 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3369 w_3263498_541854# a_3408579_674425# a_3408579_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3370 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3371 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3372 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3373 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3374 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3375 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3376 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3377 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3378 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3379 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3380 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3381 a_3408579_674425# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3382 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3383 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3384 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3385 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3386 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3387 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3388 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3389 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3390 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3391 a_3379175_716345# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3392 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3393 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3394 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3395 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3396 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3397 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3398 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3399 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3400 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3401 w_3263498_541854# a_3407435_674425# a_3407435_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3402 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3403 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3404 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3405 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3406 a_3366260_744206# a_3369760_747574# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3407 a_3359810_749958# a_3362834_747994# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3408 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3409 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3410 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3411 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3412 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3413 a_3440870_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X3414 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3415 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3416 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3417 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3418 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3419 w_3263498_541854# a_3405057_686207# w_3407323_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3420 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3421 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3422 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3423 a_3401256_686207# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3424 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3425 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3426 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3427 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3428 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3429 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3430 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3431 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3432 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3433 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3434 a_3440870_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X3435 w_3422394_717637# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3436 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3437 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3438 a_3407542_687895# a_3407542_687895# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3439 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3440 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3441 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3442 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3443 v2 a_3434368_749958# a_3428294_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3444 w_3185490_798160# a_3381660_701961# a_3381660_701961# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3445 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3446 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3447 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3448 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3449 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3450 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3451 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3452 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3453 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3454 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3455 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3456 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3457 a_3403286_703346# a_3403001_700774# w_3403067_702950# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3458 w_3263498_541854# a_3400801_715182# w_3403067_716474# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3459 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3460 a_3420293_701761# a_3422243_697443# w_3422393_701565# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3461 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
R3 w_3185490_798160# m3_3657454_970934# sky130_fd_pr__res_generic_m4 w=7.4e+07u l=1.68e+07u
X3462 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3463 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3464 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3465 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3466 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3467 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3468 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3469 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X3470 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3471 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3472 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3473 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3474 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3475 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3476 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3477 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3478 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3479 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3480 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3481 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3482 w_3185490_798160# a_3381660_718033# a_3381660_718033# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3483 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3484 a_3335479_772599# a_3359810_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3485 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3486 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3487 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3488 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3489 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3490 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3491 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3492 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3493 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3494 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3495 a_3381660_718777# a_3381660_718033# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3496 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3497 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3498 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3499 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3500 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3501 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3502 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3503 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3504 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3505 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3506 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3507 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3508 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3509 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3510 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3511 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3512 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3513 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3514 a_3440870_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X3515 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3516 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3517 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3518 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3519 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3520 a_3367712_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X3521 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3522 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3523 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3524 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3525 a_3407435_674425# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3526 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3527 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3528 a_3335479_772599# a_3359810_749958# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3529 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3530 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3531 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3532 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3533 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3534 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3535 a_3379175_700273# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3536 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3537 w_3263498_541854# a_3405057_686207# w_3407323_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3538 w_3381441_701565# a_3361095_699281# a_3381660_701961# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3539 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3540 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3541 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3542 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3543 w_3422393_701565# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3544 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3545 w_3185490_798160# a_3403286_703346# a_3403286_704090# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3546 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3547 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3548 w_3407323_687499# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3549 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3550 a_3440870_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X3551 w_3396510_687499# a_3387775_698875# a_3394410_687695# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3552 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3553 a_3367712_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X3554 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3555 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3556 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3557 a_3403001_700774# a_3381563_717833# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X3558 w_3185490_798160# a_3434368_749958# a_3428294_754598# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3559 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3560 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3561 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3562 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3563 a_3407542_688639# a_3381563_702505# w_3407323_687499# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3564 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3565 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X3566 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3567 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3568 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3569 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3570 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3571 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3572 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3573 a_3369760_754598# a_3366260_744206# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3574 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3575 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3576 w_3185490_798160# a_3403286_703346# a_3403286_703346# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3577 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3578 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3579 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3580 w_3185490_798160# a_3439418_744112# a_3443016_749796# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3581 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3582 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3583 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3584 a_3420293_701761# a_3420293_701761# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3585 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3586 a_3381660_701961# a_3381660_701961# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3587 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3588 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3589 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3590 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3591 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3592 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3593 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3594 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3595 w_3185490_798160# a_3399027_674337# a_3407435_674425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X3596 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3597 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3598 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3599 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3600 w_3263498_541854# a_3379175_716345# w_3381441_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3601 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3602 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3603 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3604 a_3420294_717833# a_3381563_717833# w_3422394_717637# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3605 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3606 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3607 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3608 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3609 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3610 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3611 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3612 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3613 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3614 a_3379175_716345# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3615 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3616 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3617 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3618 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3619 a_3400801_701658# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X3620 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3621 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3622 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3623 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3624 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3625 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3626 a_3421607_697443# a_3421925_698875# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X3627 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3628 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3629 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3630 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3631 a_3407542_687895# a_3407282_686697# w_3407323_687499# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3632 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3633 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3634 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3635 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3636 a_3381660_702705# a_3381563_702505# w_3381441_701565# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3637 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3638 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3639 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3640 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3641 w_3263498_541854# a_3405057_686207# a_3405057_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3642 a_3394410_690671# a_3394410_687695# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3643 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3644 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3645 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3646 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3647 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3648 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3649 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3650 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3651 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3652 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3653 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3654 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3655 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3656 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3657 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3658 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3659 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3660 w_3185490_798160# a_3399027_674337# a_3401256_686207# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X3661 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3662 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3663 a_3367712_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X3664 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3665 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3666 a_3381660_718033# a_3381563_717833# w_3381441_717637# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3667 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3668 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3669 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3670 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3671 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3672 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3673 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X3674 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3675 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3676 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3677 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3678 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3679 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3680 a_3407542_688639# a_3407542_687895# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3681 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X3682 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3683 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3684 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3685 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3686 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3687 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3688 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3689 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3690 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3691 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3692 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3693 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3694 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3695 w_3422394_717637# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3696 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3697 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3698 w_3422394_717637# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3699 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3700 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3701 w_3263498_541854# a_3400801_715182# a_3400801_715182# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3702 v2 a_3439418_744112# a_3443016_749796# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3703 a_3428294_754598# a_3434368_749958# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3704 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3705 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3706 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3707 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3708 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3709 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3710 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3711 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3712 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3713 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3714 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3715 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3716 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3717 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3718 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3719 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3720 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3721 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3722 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3723 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3724 a_3422243_697443# a_3420381_704937# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X3725 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3726 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3727 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3728 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3729 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3730 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3731 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3732 a_3440870_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X3733 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3734 w_3407323_687499# a_3407282_686697# a_3407542_687895# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3735 a_3407542_687895# a_3407542_687895# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3736 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3737 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3738 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3739 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3740 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3741 w_3381441_717637# a_3379272_706425# a_3381660_718777# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3742 w_3396510_687499# a_3387775_698875# a_3394410_687695# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3743 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3744 a_3428294_754598# a_3434368_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3745 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3746 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3747 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3748 w_3396510_687499# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3749 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3750 v2 a_3366260_744206# a_3369760_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3751 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3752 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3753 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3754 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3755 a_3440870_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X3756 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3757 w_3263498_541854# a_3401256_686207# a_3401256_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3758 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3759 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3760 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3761 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3762 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3763 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3764 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3765 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3766 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3767 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3768 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3769 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3770 v2 a_3366260_744206# a_3369760_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3771 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3772 w_3263498_541854# a_3400801_701658# w_3403067_702950# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3773 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3774 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3775 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3776 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3777 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3778 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3779 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3780 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3781 v2 a_3366260_744206# a_3362906_746854# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3782 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3783 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3784 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3785 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3786 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3787 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3788 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3789 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3790 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3791 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3792 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3793 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3794 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3795 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3796 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3797 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3798 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3799 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3800 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3801 a_3407435_674425# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X3802 a_3403001_700774# a_3381563_717833# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X3803 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3804 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3805 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3806 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3807 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3808 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3809 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3810 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3811 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3812 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3813 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3814 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3815 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3816 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3817 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3818 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3819 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3820 w_3422394_717637# a_3381563_717833# a_3420294_717833# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3821 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3822 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3823 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3824 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3825 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3826 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3827 a_3403286_717614# a_3403286_716870# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3828 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3829 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3830 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3831 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3832 v2 a_3359810_749958# a_3335479_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3833 a_3420294_720809# a_3420381_704937# w_3422394_717637# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3834 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3835 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3836 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3837 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3838 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3839 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3840 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3841 w_3263498_541854# a_3379175_716345# w_3381441_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3842 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3843 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3844 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3845 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3846 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3847 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3848 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3849 w_3185490_798160# a_3399027_674337# a_3399027_674337# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X3850 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3851 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3852 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3853 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3854 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3855 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3856 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3857 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3858 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3859 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3860 w_3381441_701565# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3861 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3862 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3863 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3864 w_3407323_687499# a_3407282_686697# a_3407542_687895# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3865 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3866 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3867 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3868 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3869 v2 a_3359810_749958# a_3335479_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3870 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3871 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3872 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3873 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3874 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3875 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3876 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3877 w_3396510_687499# a_3263636_541992# a_3394410_690671# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3878 a_3405057_686207# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3879 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3880 a_3367712_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X3881 a_3381660_702705# a_3381563_702505# w_3381441_701565# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3882 v2 a_3434368_749958# a_3428294_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3883 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3884 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3885 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3886 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3887 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3888 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3889 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3890 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3891 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3892 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3893 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3894 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3895 w_3381441_717637# a_3381563_717833# a_3381660_718033# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3896 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3897 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3898 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3899 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3900 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3901 a_3381660_718777# a_3379272_706425# w_3381441_717637# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3902 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3903 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3904 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3905 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3906 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3907 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3908 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3909 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3910 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3911 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3912 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3913 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3914 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3915 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3916 w_3263498_541854# a_3401256_686207# w_3396510_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3917 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3918 a_3439418_744112# a_3442918_747574# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3919 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3920 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3921 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3922 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3923 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3924 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3925 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3926 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3927 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3928 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3929 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3930 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3931 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3932 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3933 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3934 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3935 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3936 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3937 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3938 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3939 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3940 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3941 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3942 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3943 w_3185490_798160# a_3407542_687895# a_3407542_687895# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3944 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3945 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3946 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3947 a_3369760_754598# a_3366260_744206# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3948 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3949 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3950 w_3185490_798160# a_3403286_703346# a_3403286_704090# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3951 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3952 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3953 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3954 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3955 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3956 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3957 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3958 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3959 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3960 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3961 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3962 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3963 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3964 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3965 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3966 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3967 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3968 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3969 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3970 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3971 w_3185490_798160# a_3403286_703346# a_3403286_703346# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3972 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3973 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3974 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3975 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3976 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3977 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3978 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3979 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3980 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3981 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3982 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3983 w_3185490_798160# a_3381660_701961# a_3381660_702705# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3984 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3985 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3986 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3987 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3988 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3989 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3990 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3991 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3992 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3993 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3994 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3995 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3996 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3997 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3998 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3999 w_3263498_541854# a_3400801_715182# w_3403067_716474# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4000 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4001 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4002 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4003 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4004 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4005 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4006 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4007 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4008 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4009 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4010 a_3361095_699281# a_3385867_698875# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X4011 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4012 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4013 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4014 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4015 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4016 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4017 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4018 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4019 a_3361095_699281# a_3379272_706425# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X4020 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4021 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4022 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4023 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4024 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4025 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4026 w_3263498_541854# a_3379175_700273# a_3379175_700273# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4027 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4028 w_3407323_687499# a_3381563_702505# a_3407542_688639# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4029 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4030 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4031 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4032 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4033 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4034 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4035 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4036 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4037 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4038 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4039 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4040 w_3396510_687499# a_3263636_541992# a_3394410_690671# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4041 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4042 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4043 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4044 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4045 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4046 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4047 a_3403286_717614# a_3403286_716870# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4048 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4049 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4050 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4051 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4052 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4053 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4054 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4055 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4056 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4057 a_3407435_674425# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4058 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4059 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4060 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4061 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4062 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4063 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4064 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4065 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4066 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4067 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4068 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4069 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4070 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4071 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4072 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4073 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4074 w_3381441_701565# a_3381563_702505# a_3381660_702705# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4075 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4076 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4077 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4078 w_3422393_701565# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4079 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4080 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4081 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4082 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4083 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4084 w_3185490_798160# a_3403286_703346# a_3403286_703346# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4085 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4086 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4087 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4088 w_3263498_541854# a_3400801_701658# a_3400801_701658# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4089 w_3396510_687499# a_3263636_541992# a_3394410_690671# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4090 w_3185490_798160# a_3399027_674337# a_3407435_674425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X4091 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4092 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4093 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4094 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4095 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4096 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4097 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4098 a_3443016_749796# a_3439418_744112# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4099 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4100 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4101 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4102 a_3394410_690671# a_3394410_687695# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4103 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4104 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4105 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4106 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4107 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4108 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4109 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4110 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4111 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4112 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4113 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4114 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4115 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4116 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4117 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4118 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4119 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4120 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4121 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4122 a_3400801_701658# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X4123 a_3394410_687695# a_3394410_687695# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4124 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4125 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4126 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4127 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4128 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4129 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4130 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4131 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4132 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4133 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4134 w_3263498_541854# a_3379175_716345# w_3381441_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4135 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4136 w_3263498_541854# a_3401256_686207# a_3401256_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4137 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4138 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4139 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4140 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4141 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4142 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4143 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4144 w_3403067_702950# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4145 w_3381441_717637# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4146 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4147 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4148 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4149 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4150 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4151 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4152 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4153 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4154 w_3403067_702950# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4155 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4156 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4157 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4158 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4159 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4160 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4161 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4162 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4163 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4164 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4165 w_3185490_798160# a_3399027_674337# a_3401256_686207# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X4166 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4167 a_3381660_701961# a_3361095_699281# w_3381441_701565# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4168 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4169 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4170 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4171 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4172 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4173 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4174 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4175 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4176 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4177 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4178 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4179 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4180 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4181 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4182 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4183 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4184 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4185 a_3420293_701761# a_3420293_701761# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4186 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4187 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4188 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4189 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4190 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4191 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4192 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4193 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4194 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4195 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4196 w_3185490_798160# a_3381563_702505# sky130_fd_pr__diode_pw2nd_05v5 area=2.25e+16p
X4197 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4198 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4199 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4200 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4201 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4202 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4203 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4204 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4205 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4206 w_3263498_541854# a_3408579_674425# a_3408579_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4207 a_3436064_746854# a_3439418_744112# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4208 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4209 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4210 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4211 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4212 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4213 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4214 a_3408579_674425# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4215 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4216 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4217 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4218 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4219 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4220 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4221 w_3185490_798160# a_3381660_701961# a_3381660_701961# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4222 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4223 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4224 a_3407542_687895# a_3407542_687895# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4225 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4226 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4227 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4228 w_3403067_716474# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4229 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4230 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4231 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4232 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4233 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4234 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4235 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4236 w_3263498_541854# a_3400801_715182# a_3400801_715182# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4237 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4238 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4239 a_3420293_701761# a_3422243_697443# w_3422393_701565# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4240 w_3185490_798160# a_3362834_747994# a_3359810_749958# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4241 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4242 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4243 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4244 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4245 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4246 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4247 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4248 w_3185490_798160# a_3420293_701761# a_3420293_704737# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4249 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4250 a_3404273_699542# a_3404591_700774# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X4251 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4252 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4253 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4254 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4255 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4256 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4257 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4258 a_3428294_754598# a_3434368_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4259 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4260 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4261 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4262 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4263 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4264 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4265 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4266 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4267 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4268 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4269 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4270 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4271 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4272 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4273 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4274 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4275 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4276 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4277 w_3407323_687499# a_3381563_702505# a_3407542_688639# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4278 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4279 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4280 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4281 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4282 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4283 a_3428294_754598# a_3434368_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4284 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4285 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4286 w_3263498_541854# a_3379175_700273# a_3379175_700273# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4287 a_3441490_744142# a_3440844_744112# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4288 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4289 w_3396510_687499# a_3263636_541992# a_3394410_690671# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4290 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4291 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4292 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4293 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4294 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4295 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4296 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4297 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4298 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4299 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4300 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4301 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4302 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4303 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4304 a_3386821_697443# a_3386503_698875# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X4305 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4306 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4307 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4308 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4309 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4310 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4311 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4312 w_3185490_798160# a_3399027_674337# a_3379175_716345# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X4313 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4314 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4315 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4316 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4317 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4318 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4319 w_3381441_701565# a_3361095_699281# a_3381660_701961# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4320 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4321 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4322 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4323 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4324 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4325 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4326 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4327 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4328 a_3407435_674425# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4329 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4330 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4331 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4332 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4333 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4334 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4335 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4336 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4337 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4338 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4339 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4340 a_3420294_717833# a_3420294_717833# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4341 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4342 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4343 v2 a_3359810_749958# a_3335479_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4344 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4345 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4346 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4347 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4348 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4349 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4350 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4351 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4352 a_3362906_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X4353 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4354 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4355 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4356 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4357 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4358 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4359 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4360 a_3405389_721804# a_3403286_717614# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=500000u
X4361 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4362 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4363 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4364 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4365 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4366 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4367 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4368 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4369 w_3185490_798160# a_3394410_687695# a_3394410_687695# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4370 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4371 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4372 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4373 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4374 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4375 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4376 a_3381660_718777# a_3381660_718033# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4377 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4378 a_3401256_686207# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4379 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4380 w_3185490_798160# a_3359810_749958# a_3335479_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4381 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4382 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4383 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4384 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4385 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4386 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4387 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4388 a_3403286_716870# a_3403286_716870# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4389 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4390 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4391 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4392 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4393 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4394 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4395 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4396 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4397 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4398 w_3263498_541854# a_3379175_716345# w_3381441_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4399 w_3185490_798160# a_3420294_717833# a_3420294_720809# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4400 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4401 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4402 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4403 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4404 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4405 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4406 w_3422393_701565# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4407 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4408 w_3381441_717637# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4409 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4410 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4411 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4412 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4413 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4414 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4415 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4416 w_3422393_701565# a_3381563_702505# a_3420293_704737# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4417 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4418 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4419 w_3381441_701565# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4420 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4421 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4422 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4423 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4424 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4425 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4426 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4427 a_3405057_686207# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4428 v2 a_3366260_744206# a_3369760_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4429 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4430 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4431 w_3403067_702950# a_3381563_702505# a_3403286_704090# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4432 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4433 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4434 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4435 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4436 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4437 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4438 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4439 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4440 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4441 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4442 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4443 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4444 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4445 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4446 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4447 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4448 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4449 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4450 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4451 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4452 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4453 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4454 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4455 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4456 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4457 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4458 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4459 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4460 a_3443016_749796# a_3439418_744112# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4461 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4462 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4463 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4464 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4465 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4466 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4467 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4468 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4469 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4470 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4471 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4472 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4473 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4474 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4475 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4476 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4477 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4478 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4479 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4480 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4481 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4482 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4483 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4484 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4485 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4486 a_3422243_697443# a_3420381_704937# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X4487 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4488 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4489 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4490 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4491 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4492 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4493 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4494 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4495 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4496 a_3446663_700871# a_3448095_700553# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X4497 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4498 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4499 a_3420335_697443# a_3420653_698875# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X4500 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4501 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4502 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4503 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4504 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4505 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4506 w_3263498_541854# a_3407435_674425# a_3407435_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4507 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4508 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4509 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4510 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4511 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4512 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4513 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4514 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4515 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4516 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4517 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4518 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4519 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4520 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4521 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4522 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4523 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4524 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4525 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4526 w_3185490_798160# a_3399027_674337# a_3400801_701658# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X4527 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4528 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4529 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4530 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4531 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4532 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4533 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4534 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4535 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4536 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4537 w_3185490_798160# a_3434368_749958# a_3428294_754598# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4538 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4539 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4540 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4541 w_3422394_717637# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4542 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4543 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4544 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4545 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4546 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4547 w_3422394_717637# a_3420381_704937# a_3420294_720809# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4548 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4549 w_3185490_798160# a_3420294_717833# a_3420294_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4550 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4551 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4552 w_3263498_541854# a_3400801_715182# w_3403067_716474# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4553 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4554 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4555 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4556 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4557 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4558 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4559 a_3400801_715182# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X4560 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4561 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4562 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4563 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
R4 a_3285528_930602# m3_3215040_970024# sky130_fd_pr__res_generic_m3 w=2.505e+07u l=6.55e+06u
X4564 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4565 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4566 a_3420294_720809# a_3420294_717833# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4567 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4568 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4569 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4570 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4571 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4572 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4573 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4574 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4575 w_3185490_798160# a_3420293_701761# a_3420293_701761# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4576 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4577 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4578 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4579 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4580 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4581 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4582 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4583 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4584 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4585 w_3185490_798160# a_3381660_718033# a_3381660_718777# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4586 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4587 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4588 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4589 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4590 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4591 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4592 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4593 v2 a_3434368_749958# a_3428294_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4594 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4595 w_3263498_541854# a_3379175_700273# a_3379175_700273# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4596 w_3422393_701565# a_3381563_702505# a_3420293_704737# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4597 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4598 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4599 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4600 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4601 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4602 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4603 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4604 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4605 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4606 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4607 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4608 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4609 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4610 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4611 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4612 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4613 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4614 a_3369760_754598# a_3366260_744206# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4615 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4616 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4617 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4618 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4619 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4620 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4621 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4622 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4623 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4624 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4625 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4626 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4627 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4628 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4629 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4630 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4631 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4632 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4633 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4634 a_3379175_700273# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4635 w_3263498_541854# a_3408579_674425# a_3408579_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4636 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4637 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4638 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4639 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4640 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4641 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4642 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4643 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4644 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4645 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4646 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4647 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4648 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4649 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4650 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4651 a_3368332_744142# a_3359810_749958# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4652 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4653 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4654 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4655 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4656 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4657 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4658 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4659 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4660 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4661 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4662 a_3403001_700774# a_3381563_717833# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X4663 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4664 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4665 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4666 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4667 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4668 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4669 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4670 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4671 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4672 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4673 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4674 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4675 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4676 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4677 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4678 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4679 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4680 w_3185490_798160# a_3263636_541992# sky130_fd_pr__diode_pw2nd_05v5 area=2.25e+16p
X4681 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4682 a_3420294_720809# a_3420381_704937# w_3422394_717637# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4683 a_3443016_749796# a_3439418_744112# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4684 a_3335479_772599# a_3359810_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4685 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4686 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4687 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4688 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4689 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4690 a_3263636_541992# a_3408714_686379# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X4691 w_3185490_798160# a_3420294_717833# a_3420294_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4692 w_3185490_798160# a_3381660_701961# a_3381660_702705# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4693 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4694 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4695 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4696 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4697 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4698 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4699 a_3428294_754598# a_3434368_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4700 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4701 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4702 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4703 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4704 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4705 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4706 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4707 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4708 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4709 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4710 w_3422393_701565# a_3422243_697443# a_3420293_701761# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4711 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4712 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4713 w_3422394_717637# a_3420381_704937# a_3420294_720809# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4714 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4715 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4716 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4717 w_3407323_687499# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4718 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4719 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4720 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4721 a_3407542_688639# a_3381563_702505# w_3407323_687499# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4722 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4723 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4724 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4725 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4726 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4727 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4728 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4729 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4730 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4731 w_3263498_541854# a_3405057_686207# a_3405057_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4732 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4733 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4734 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4735 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4736 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4737 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4738 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4739 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4740 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4741 v2 a_3442918_747574# a_3439418_744112# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4742 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4743 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4744 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4745 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4746 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4747 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4748 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4749 a_3381660_718777# a_3379272_706425# w_3381441_717637# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4750 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4751 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4752 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4753 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4754 w_3185490_798160# a_3394410_687695# a_3394410_687695# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4755 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4756 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4757 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4758 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4759 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4760 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4761 w_3263498_541854# a_3400801_715182# a_3400801_715182# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4762 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4763 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4764 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4765 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4766 w_3185490_798160# a_3369760_747574# a_3366260_744206# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4767 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4768 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4769 a_3394410_687695# a_3387775_698875# w_3396510_687499# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4770 w_3263498_541854# a_3400801_715182# a_3400801_715182# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4771 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4772 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4773 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4774 a_3361095_699281# a_3379272_706425# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X4775 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4776 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4777 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4778 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4779 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4780 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4781 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4782 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4783 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4784 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4785 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4786 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4787 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4788 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4789 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4790 w_3185490_798160# a_3399027_674337# a_3379175_716345# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X4791 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4792 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4793 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4794 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4795 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4796 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4797 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4798 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4799 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4800 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4801 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4802 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4803 a_3407542_688639# a_3407542_687895# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4804 w_3263498_541854# a_3379175_700273# a_3379175_700273# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4805 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4806 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4807 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4808 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4809 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4810 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4811 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4812 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4813 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4814 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4815 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4816 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4817 v2 a_3434368_749958# a_3440870_744142# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4818 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4819 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4820 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4821 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4822 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4823 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4824 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4825 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4826 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4827 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4828 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4829 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4830 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4831 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4832 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4833 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4834 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4835 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4836 w_3263498_541854# a_3408579_674425# w_3422394_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4837 w_3422394_717637# a_3381563_717833# a_3420294_717833# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4838 a_3407435_674425# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4839 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4840 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4841 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4842 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4843 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4844 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4845 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4846 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4847 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4848 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4849 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4850 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4851 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4852 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4853 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4854 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4855 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4856 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4857 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4858 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4859 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4860 w_3185490_798160# a_3381660_718033# a_3381660_718033# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4861 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4862 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4863 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4864 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4865 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4866 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4867 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4868 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4869 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4870 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4871 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4872 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4873 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4874 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4875 w_3422393_701565# a_3422243_697443# a_3420293_701761# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4876 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4877 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4878 a_3401256_686207# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4879 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4880 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4881 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4882 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4883 a_3440870_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X4884 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4885 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4886 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4887 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4888 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4889 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4890 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4891 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4892 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4893 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4894 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4895 a_3400801_701658# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4896 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4897 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4898 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4899 w_3422393_701565# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4900 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4901 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4902 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4903 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4904 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4905 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4906 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4907 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4908 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4909 a_3440870_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X4910 a_3381660_701961# a_3361095_699281# w_3381441_701565# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4911 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4912 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4913 v2 a_3439418_744112# a_3443016_749796# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4914 a_3428294_754598# a_3434368_749958# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4915 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4916 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4917 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4918 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4919 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4920 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4921 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4922 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4923 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4924 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4925 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4926 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4927 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4928 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4929 a_3420293_701761# a_3420293_701761# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4930 w_3403067_702950# a_3403001_700774# a_3403286_703346# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4931 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4932 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4933 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4934 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4935 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4936 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4937 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4938 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4939 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4940 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4941 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4942 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4943 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4944 a_3383521_705357# a_3379272_706425# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=1.4e+07u
X4945 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4946 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4947 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4948 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4949 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4950 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4951 a_3420294_717833# a_3420294_717833# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4952 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4953 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4954 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4955 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4956 a_3422243_697443# a_3420381_704937# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X4957 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4958 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4959 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4960 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4961 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4962 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4963 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4964 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4965 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4966 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4967 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4968 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4969 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4970 w_3396510_687499# a_3387775_698875# a_3394410_687695# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4971 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4972 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4973 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4974 a_3366260_744112# a_3366422_743586# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4975 w_3185490_798160# a_3399027_674337# a_3400801_701658# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X4976 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4977 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4978 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4979 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4980 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4981 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4982 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4983 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4984 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4985 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4986 w_3185490_798160# a_3381660_701961# a_3381660_701961# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4987 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4988 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4989 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4990 w_3263498_541854# a_3407435_674425# a_3407435_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4991 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4992 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4993 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4994 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4995 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4996 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4997 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4998 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4999 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5000 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5001 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5002 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5003 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5004 w_3422394_717637# a_3381563_717833# a_3420294_717833# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5005 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5006 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5007 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5008 a_3400801_715182# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5009 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5010 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5011 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5012 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5013 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5014 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X5015 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5016 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5017 a_3367712_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X5018 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5019 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5020 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5021 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5022 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5023 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5024 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5025 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5026 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5027 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5028 a_3381660_718033# a_3381563_717833# w_3381441_717637# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5029 w_3185490_798160# a_3403286_703346# a_3403286_704090# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5030 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
R5 w_3185490_798160# m3_3713300_450024# sky130_fd_pr__res_generic_m4 w=7.815e+07u l=1.755e+07u
X5031 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5032 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5033 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5034 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5035 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5036 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5037 w_3185490_798160# a_3394410_687695# a_3394410_690671# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5038 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5039 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5040 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5041 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5042 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5043 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5044 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5045 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5046 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5047 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5048 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5049 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X5050 v2 a_3434368_749958# a_3428294_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5051 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5052 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5053 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5054 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5055 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5056 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5057 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5058 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5059 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5060 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5061 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5062 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5063 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5064 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5065 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5066 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5067 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5068 w_3185490_798160# a_3420293_701761# a_3420293_704737# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5069 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5070 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5071 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5072 w_3263498_541854# a_3405057_686207# a_3405057_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5073 w_3381441_701565# a_3381563_702505# a_3381660_702705# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5074 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5075 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5076 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5077 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5078 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5079 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5080 v2 a_3434368_749958# a_3428294_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5081 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5082 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5083 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5084 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5085 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5086 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5087 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5088 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5089 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5090 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5091 a_3403286_716870# a_3403286_716870# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5092 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5093 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5094 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5095 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5096 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5097 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5098 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5099 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5100 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5101 a_3335479_772599# a_3359810_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5102 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5103 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5104 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5105 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5106 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5107 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5108 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5109 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5110 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5111 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5112 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5113 a_3407435_674425# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5114 a_3335479_772599# a_3359810_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5115 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5116 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5117 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5118 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5119 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5120 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5121 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5122 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5123 a_3379175_700273# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5124 w_3263498_541854# a_3408579_674425# a_3408579_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5125 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5126 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5127 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5128 a_3335479_772599# a_3359810_749958# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5129 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5130 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5131 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5132 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5133 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5134 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5135 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X5136 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5137 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5138 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X5139 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5140 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5141 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5142 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5143 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5144 a_3335479_772599# a_3359810_749958# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5145 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5146 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5147 a_3369760_754598# a_3366260_744206# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5148 v2 a_3366422_743586# a_3367712_744142# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5149 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5150 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5151 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5152 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5153 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5154 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5155 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5156 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5157 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5158 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5159 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5160 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5161 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5162 a_3369760_754598# a_3366260_744206# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5163 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5164 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5165 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5166 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5167 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5168 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5169 w_3396510_687499# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5170 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5171 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5172 a_3394410_690671# a_3394410_687695# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5173 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5174 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5175 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5176 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5177 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5178 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5179 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5180 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5181 w_3263498_541854# a_3400801_715182# w_3403067_716474# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5182 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5183 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5184 w_3263498_541854# a_3401256_686207# a_3401256_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5185 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5186 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5187 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5188 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5189 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5190 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5191 w_3403067_702950# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5192 a_3369760_754598# a_3366260_744206# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5193 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5194 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5195 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5196 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5197 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5198 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5199 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5200 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5201 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5202 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5203 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5204 a_3407542_688639# a_3407542_687895# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5205 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5206 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5207 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5208 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5209 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5210 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5211 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5212 w_3422393_701565# a_3381563_702505# a_3420293_704737# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5213 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5214 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5215 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5216 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5217 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5218 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5219 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5220 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5221 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5222 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5223 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5224 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5225 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5226 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5227 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5228 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5229 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5230 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5231 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5232 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5233 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5234 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5235 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5236 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5237 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5238 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5239 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5240 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5241 v2 a_3439418_744112# a_3443016_749796# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5242 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5243 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5244 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5245 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X5246 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5247 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5248 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X5249 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5250 w_3396510_687499# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5251 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5252 a_3361095_699281# a_3379272_706425# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X5253 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5254 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5255 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5256 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5257 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5258 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5259 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5260 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5261 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5262 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5263 a_3407542_687895# a_3407542_687895# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5264 w_3185490_798160# a_3394410_687695# a_3394410_690671# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5265 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5266 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5267 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5268 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5269 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5270 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5271 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5272 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5273 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5274 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5275 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5276 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5277 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5278 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5279 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5280 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5281 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5282 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5283 a_3403637_699542# a_3403955_700774# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X5284 w_3263498_541854# a_3400801_715182# a_3400801_715182# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5285 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5286 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5287 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5288 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5289 a_3399027_674337# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5290 w_3185490_798160# a_3420293_701761# a_3420293_701761# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5291 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5292 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5293 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5294 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5295 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5296 w_3185490_798160# a_3366260_744206# a_3369760_754598# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5297 a_3366260_744112# a_3366422_743586# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5298 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5299 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5300 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5301 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5302 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5303 w_3403067_716474# a_3403189_717414# a_3403286_717614# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5304 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5305 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5306 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5307 a_3405532_706743# a_3403286_704090# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=1.4e+06u
X5308 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5309 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5310 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5311 w_3263498_541854# a_3379175_700273# w_3381441_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5312 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5313 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5314 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5315 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5316 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5317 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5318 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5319 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5320 w_3185490_798160# a_3399027_674337# a_3379175_700273# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5321 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5322 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5323 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5324 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5325 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5326 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5327 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5328 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5329 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5330 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5331 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5332 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5333 a_3369760_747574# a_3367712_744142# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5334 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5335 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5336 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5337 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5338 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5339 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5340 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5341 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5342 a_3408579_674425# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5343 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5344 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5345 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5346 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5347 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5348 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5349 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5350 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5351 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X5352 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5353 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5354 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5355 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5356 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5357 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5358 w_3263498_541854# a_3408579_674425# w_3422394_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5359 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5360 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5361 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5362 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5363 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5364 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5365 w_3263498_541854# a_3405057_686207# a_3405057_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5366 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5367 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5368 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5369 w_3263498_541854# a_3400801_701658# w_3403067_702950# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5370 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5371 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5372 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5373 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5374 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5375 a_3420294_720809# a_3420294_717833# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5376 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5377 a_3422243_697443# a_3448095_699281# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X5378 a_3443016_749796# a_3439418_744112# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5379 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5380 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5381 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5382 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5383 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5384 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5385 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5386 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5387 w_3381441_701565# a_3361095_699281# a_3381660_701961# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5388 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5389 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5390 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5391 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5392 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5393 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5394 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5395 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5396 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5397 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5398 a_3420294_717833# a_3420294_717833# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5399 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5400 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5401 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5402 w_3422393_701565# a_3381563_702505# a_3420293_704737# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5403 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5404 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5405 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5406 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5407 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5408 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5409 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5410 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5411 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5412 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5413 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5414 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5415 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5416 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5417 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5418 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5419 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5420 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5421 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5422 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5423 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5424 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5425 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5426 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5427 a_3422243_697443# a_3420381_704937# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X5428 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5429 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5430 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5431 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5432 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5433 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5434 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5435 a_3400801_701658# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5436 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5437 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5438 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5439 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5440 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5441 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5442 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5443 w_3263498_541854# a_3400801_715182# w_3403067_716474# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5444 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5445 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5446 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5447 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5448 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5449 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5450 w_3422393_701565# a_3422243_697443# a_3420293_701761# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5451 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5452 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5453 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5454 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5455 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5456 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5457 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5458 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5459 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5460 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5461 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5462 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5463 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5464 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5465 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5466 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5467 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5468 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5469 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5470 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5471 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5472 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5473 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5474 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5475 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5476 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5477 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5478 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5479 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5480 w_3185490_798160# a_3407542_687895# a_3407542_687895# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5481 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5482 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5483 w_3185490_798160# a_3420294_717833# a_3420294_720809# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5484 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5485 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5486 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5487 w_3403067_716474# a_3403189_717414# a_3403286_717614# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5488 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5489 a_3420293_701761# a_3422243_697443# w_3422393_701565# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5490 w_3185490_798160# a_3439418_744112# a_3443016_749796# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5491 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5492 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5493 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5494 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5495 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5496 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5497 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5498 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5499 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5500 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5501 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5502 w_3185490_798160# a_3399027_674337# a_3400801_715182# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5503 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5504 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5505 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5506 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5507 v2 a_3434368_749958# a_3428294_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5508 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5509 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5510 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5511 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5512 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5513 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5514 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5515 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5516 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5517 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5518 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5519 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5520 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5521 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5522 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5523 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5524 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5525 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5526 w_3185490_798160# a_3381660_701961# a_3381660_702705# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5527 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5528 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5529 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5530 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5531 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5532 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5533 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5534 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5535 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5536 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5537 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5538 w_3381441_717637# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5539 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5540 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5541 a_3379175_700273# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5542 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5543 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5544 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5545 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5546 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5547 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5548 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5549 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5550 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5551 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5552 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5553 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5554 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5555 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5556 w_3263498_541854# a_3379175_700273# w_3381441_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5557 a_3359663_700553# a_3361095_700871# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X5558 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5559 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5560 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5561 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5562 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5563 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5564 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5565 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5566 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5567 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5568 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5569 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5570 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5571 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5572 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5573 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5574 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5575 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5576 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5577 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5578 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5579 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5580 a_3366260_744206# a_3369760_747574# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5581 w_3185490_798160# a_3399027_674337# a_3408579_674425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5582 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5583 w_3381441_717637# a_3379272_706425# a_3381660_718777# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5584 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5585 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5586 a_3381660_718033# a_3381660_718033# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5587 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5588 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5589 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5590 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5591 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5592 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5593 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5594 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5595 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5596 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5597 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5598 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5599 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5600 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5601 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5602 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5603 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5604 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5605 a_3403286_704090# a_3381563_702505# w_3403067_702950# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5606 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5607 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5608 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5609 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5610 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5611 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5612 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5613 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5614 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5615 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5616 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5617 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5618 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5619 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5620 a_3405057_686207# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5621 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5622 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5623 w_3185490_798160# a_3420294_717833# a_3420294_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5624 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5625 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5626 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5627 w_3403067_716474# a_3381563_702505# a_3403286_716870# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5628 a_3443016_749796# a_3439418_744112# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5629 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5630 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5631 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5632 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5633 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5634 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5635 a_3420294_720809# a_3420294_717833# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5636 v2 a_3440870_744142# a_3442918_747574# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5637 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5638 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5639 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5640 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5641 a_3420294_717833# a_3381563_717833# w_3422394_717637# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5642 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5643 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5644 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5645 w_3422393_701565# a_3422243_697443# a_3420293_701761# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5646 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5647 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5648 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5649 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5650 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5651 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5652 a_3394410_690671# a_3263636_541992# w_3396510_687499# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5653 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5654 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5655 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5656 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5657 a_3446663_699599# a_3448095_699917# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X5658 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5659 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5660 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5661 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5662 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5663 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5664 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5665 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5666 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5667 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5668 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5669 a_3407435_674425# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5670 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5671 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5672 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5673 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5674 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5675 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5676 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5677 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5678 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5679 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5680 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5681 a_3408579_674425# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5682 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5683 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5684 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5685 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5686 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5687 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5688 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5689 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5690 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5691 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5692 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5693 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5694 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5695 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5696 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5697 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5698 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5699 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5700 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5701 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5702 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5703 a_3422243_697443# a_3420381_704937# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X5704 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5705 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5706 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5707 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5708 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5709 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5710 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5711 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5712 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5713 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5714 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5715 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5716 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5717 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5718 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5719 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5720 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5721 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5722 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5723 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5724 a_3443016_749796# a_3439418_744112# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5725 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5726 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5727 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5728 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5729 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5730 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5731 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5732 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5733 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5734 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5735 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5736 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5737 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5738 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5739 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5740 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5741 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5742 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5743 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5744 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5745 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5746 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5747 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5748 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5749 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5750 a_3443016_749796# a_3439418_744112# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5751 w_3185490_798160# a_3434368_749958# a_3428294_754598# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5752 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5753 a_3361095_699281# a_3379272_706425# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X5754 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5755 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5756 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5757 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5758 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5759 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5760 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5761 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5762 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5763 w_3185490_798160# a_3381660_701961# a_3381660_701961# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5764 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5765 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5766 a_3407542_687895# a_3407542_687895# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5767 w_3403067_702950# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5768 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5769 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5770 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5771 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5772 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5773 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5774 w_3263498_541854# a_3407435_674425# w_3422393_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5775 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5776 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X5777 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5778 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5779 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5780 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5781 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5782 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5783 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5784 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5785 a_3403286_703346# a_3403001_700774# w_3403067_702950# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5786 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5787 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5788 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5789 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5790 a_3398102_692829# a_3387775_698875# sky130_fd_pr__cap_mim_m3_1 l=1.4e+07u w=1.4e+07u
X5791 w_3381441_717637# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5792 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5793 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5794 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5795 a_3399027_674337# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5796 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5797 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5798 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5799 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5800 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5801 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5802 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5803 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5804 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5805 w_3185490_798160# a_3381660_718033# a_3381660_718033# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5806 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5807 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5808 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5809 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5810 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5811 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5812 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5813 w_3403067_716474# a_3381563_702505# a_3403286_716870# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5814 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5815 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5816 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5817 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5818 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5819 a_3381660_718777# a_3381660_718033# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5820 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5821 w_3185628_834308# w_3185490_798160# sky130_fd_pr__diode_pd2nw_05v5 area=2.25e+16p
X5822 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5823 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5824 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5825 a_3407542_688639# a_3381563_702505# w_3407323_687499# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5826 a_3369760_754598# a_3366260_744206# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5827 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5828 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5829 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5830 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5831 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5832 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5833 w_3185490_798160# a_3399027_674337# a_3379175_700273# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5834 w_3263498_541854# a_3400801_715182# a_3400801_715182# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5835 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5836 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5837 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5838 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5839 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5840 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5841 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5842 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5843 a_3394410_690671# a_3263636_541992# w_3396510_687499# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5844 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5845 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5846 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5847 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5848 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5849 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5850 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5851 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5852 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5853 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5854 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5855 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5856 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5857 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5858 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5859 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5860 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5861 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5862 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5863 w_3422394_717637# a_3381563_717833# a_3420294_717833# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5864 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5865 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5866 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5867 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5868 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5869 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5870 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5871 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5872 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5873 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5874 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5875 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X5876 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5877 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5878 a_3420294_720809# a_3420381_704937# w_3422394_717637# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5879 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5880 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5881 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5882 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5883 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5884 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5885 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5886 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5887 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5888 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5889 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5890 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X5891 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5892 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5893 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5894 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5895 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5896 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5897 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5898 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5899 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
R6 v2 m3_3722410_898374# sky130_fd_pr__res_generic_m5 w=7.42e+07u l=1.77e+07u
X5900 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5901 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5902 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5903 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5904 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5905 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5906 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5907 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5908 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5909 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5910 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5911 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5912 a_3408579_674425# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5913 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5914 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5915 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5916 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5917 w_3185490_798160# a_3381660_718033# a_3381660_718777# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5918 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5919 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5920 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5921 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5922 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5923 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5924 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5925 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5926 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5927 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5928 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5929 a_3335479_772599# a_3359810_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5930 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5931 w_3263498_541854# a_3405057_686207# a_3405057_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5932 a_3428294_754598# a_3434368_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5933 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5934 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5935 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5936 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5937 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5938 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5939 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5940 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5941 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5942 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5943 a_3428294_754598# a_3434368_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5944 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5945 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5946 w_3381441_701565# a_3381563_702505# a_3381660_702705# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5947 v2 a_3359810_749958# a_3335479_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5948 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5949 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5950 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5951 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5952 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5953 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5954 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5955 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5956 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5957 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5958 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5959 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5960 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5961 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5962 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5963 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5964 v2 a_3366260_744206# a_3369760_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5965 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5966 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5967 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5968 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5969 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5970 a_3361095_699281# a_3379272_706425# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X5971 v2 a_3359810_749958# a_3335479_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5972 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5973 a_3403286_703346# a_3403001_700774# w_3403067_702950# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5974 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5975 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5976 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5977 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5978 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5979 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5980 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5981 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5982 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5983 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5984 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5985 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X5986 w_3185490_798160# a_3359810_749958# a_3335479_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5987 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X5988 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5989 a_3400801_701658# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5990 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5991 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5992 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5993 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5994 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5995 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5996 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5997 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5998 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5999 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6000 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6001 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6002 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6003 w_3381441_717637# a_3379272_706425# a_3381660_718777# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6004 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6005 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6006 w_3185490_798160# a_3359810_749958# a_3335479_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6007 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6008 w_3185490_798160# a_3403286_716870# a_3403286_717614# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6009 a_3285528_930602# v2 sky130_fd_pr__diode_pd2nw_05v5 area=2.25e+16p
X6010 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6011 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6012 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6013 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6014 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6015 w_3185490_798160# a_3366260_744206# a_3369760_754598# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6016 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6017 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6018 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6019 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6020 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6021 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6022 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6023 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6024 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6025 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6026 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6027 a_3361095_699281# a_3379272_706425# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X6028 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6029 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6030 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6031 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6032 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6033 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6034 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6035 a_3381660_701961# a_3361095_699281# w_3381441_701565# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6036 v2 a_3366260_744206# a_3369760_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6037 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6038 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6039 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6040 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6041 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6042 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6043 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6044 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6045 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6046 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6047 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6048 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6049 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6050 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6051 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6052 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6053 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6054 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6055 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6056 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6057 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6058 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6059 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6060 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6061 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6062 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6063 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6064 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6065 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6066 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6067 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6068 v2 a_3366260_744206# a_3369760_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6069 v2 a_3359810_749958# a_3335479_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6070 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6071 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6072 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6073 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6074 a_3407542_687895# a_3407542_687895# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6075 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6076 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6077 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6078 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6079 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6080 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6081 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6082 a_3400801_715182# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6083 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6084 a_3381660_702705# a_3381660_701961# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6085 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6086 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6087 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6088 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6089 a_3408579_674425# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6090 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6091 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6092 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6093 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6094 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6095 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6096 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6097 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6098 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6099 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6100 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6101 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6102 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6103 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6104 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6105 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6106 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6107 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6108 w_3185490_798160# a_3399027_674337# a_3408579_674425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6109 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6110 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6111 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6112 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6113 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6114 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6115 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6116 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6117 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6118 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6119 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6120 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6121 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6122 a_3439418_744112# a_3442918_747574# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6123 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6124 w_3396510_687499# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6125 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6126 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6127 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6128 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6129 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6130 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6131 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6132 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6133 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6134 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6135 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6136 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6137 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6138 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6139 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6140 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6141 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6142 a_3401256_686207# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6143 a_3405057_686207# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6144 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6145 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6146 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6147 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6148 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6149 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6150 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6151 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6152 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6153 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6154 a_3369760_754598# a_3366260_744206# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6155 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6156 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6157 w_3263498_541854# a_3405057_686207# w_3407323_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6158 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6159 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6160 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6161 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6162 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6163 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6164 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6165 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6166 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6167 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6168 w_3381441_701565# a_3361095_699281# a_3381660_701961# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6169 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6170 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6171 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6172 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6173 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6174 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6175 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6176 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6177 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6178 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6179 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6180 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6181 w_3403067_716474# a_3403189_717414# a_3403286_717614# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6182 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6183 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6184 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6185 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6186 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6187 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6188 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6189 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6190 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6191 a_3408579_674425# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6192 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6193 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6194 a_3420293_704737# a_3420293_701761# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6195 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6196 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6197 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6198 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6199 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6200 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6201 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6202 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6203 a_3394410_687695# a_3387775_698875# w_3396510_687499# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6204 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6205 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6206 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6207 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6208 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6209 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6210 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6211 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6212 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6213 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6214 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6215 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6216 a_3403286_716870# a_3403286_716870# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6217 a_3422243_697443# a_3420381_704937# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X6218 a_3439418_744112# a_3442918_747574# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6219 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6220 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6221 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6222 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6223 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6224 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6225 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6226 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6227 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6228 a_3401256_686207# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6229 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6230 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6231 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6232 w_3263498_541854# a_3405057_686207# a_3405057_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6233 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6234 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6235 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6236 v2 a_3439418_744112# a_3443016_749796# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6237 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6238 w_3185490_798160# a_3381660_718033# a_3381660_718033# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6239 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6240 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6241 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6242 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6243 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6244 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6245 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6246 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6247 w_3263498_541854# a_3408579_674425# a_3408579_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6248 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6249 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6250 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6251 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6252 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6253 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6254 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6255 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6256 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6257 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6258 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6259 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6260 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6261 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6262 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6263 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6264 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6265 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6266 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6267 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6268 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6269 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6270 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6271 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6272 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6273 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6274 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6275 w_3185490_798160# a_3407542_687895# a_3407542_687895# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6276 a_3420293_701761# a_3422243_697443# w_3422393_701565# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6277 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6278 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6279 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6280 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6281 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6282 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6283 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6284 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6285 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6286 w_3263498_541854# a_3408579_674425# w_3422394_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6287 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6288 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6289 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6290 a_3381660_702705# a_3381660_701961# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6291 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6292 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6293 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6294 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6295 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6296 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6297 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6298 w_3263498_541854# a_3400801_715182# w_3403067_716474# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6299 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6300 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6301 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6302 w_3263498_541854# a_3379175_716345# a_3379175_716345# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6303 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6304 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6305 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6306 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6307 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6308 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6309 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6310 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6311 a_3379175_716345# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6312 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6313 w_3381441_717637# a_3381563_717833# a_3381660_718033# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6314 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6315 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6316 a_3403286_704090# a_3381563_702505# w_3403067_702950# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6317 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6318 w_3185490_798160# a_3403286_716870# a_3403286_716870# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6319 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6320 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6321 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6322 w_3185490_798160# a_3403286_703346# a_3403286_704090# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6323 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6324 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6325 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6326 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6327 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6328 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6329 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6330 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6331 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6332 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6333 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6334 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6335 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6336 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6337 w_3396510_687499# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6338 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6339 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6340 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6341 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6342 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6343 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6344 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6345 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6346 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6347 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6348 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6349 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6350 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6351 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6352 w_3403067_716474# a_3403189_717414# a_3403286_717614# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6353 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6354 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6355 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6356 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6357 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6358 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X6359 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6360 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6361 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6362 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6363 a_3407542_688639# a_3407542_687895# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6364 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6365 a_3407542_687895# a_3407282_686697# w_3407323_687499# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6366 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6367 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6368 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6369 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6370 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6371 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6372 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6373 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6374 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6375 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6376 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6377 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6378 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6379 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6380 w_3263498_541854# a_3400801_715182# a_3400801_715182# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6381 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6382 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6383 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6384 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6385 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6386 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6387 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6388 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6389 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6390 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6391 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6392 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6393 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6394 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6395 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6396 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6397 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6398 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6399 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6400 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6401 w_3403067_716474# a_3381563_702505# a_3403286_716870# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6402 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6403 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6404 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6405 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6406 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6407 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6408 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6409 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6410 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6411 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6412 w_3263498_541854# a_3379175_700273# w_3381441_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6413 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6414 a_3420293_704737# a_3420293_701761# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6415 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6416 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6417 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6418 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6419 w_3185490_798160# a_3369760_747574# a_3366260_744206# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6420 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6421 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6422 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6423 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6424 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6425 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6426 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6427 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6428 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6429 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6430 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6431 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6432 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6433 w_3403067_702950# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6434 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6435 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6436 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6437 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6438 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6439 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6440 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6441 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6442 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6443 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6444 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6445 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6446 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6447 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6448 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6449 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6450 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6451 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6452 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6453 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6454 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6455 w_3185490_798160# a_3439418_744112# a_3443016_749796# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6456 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6457 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6458 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6459 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6460 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6461 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6462 a_3403286_703346# a_3403286_703346# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6463 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6464 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6465 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6466 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6467 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6468 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X6469 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6470 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6471 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6472 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6473 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6474 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6475 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6476 a_3420294_720809# a_3420294_717833# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6477 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6478 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6479 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6480 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6481 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6482 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6483 w_3185490_798160# a_3399027_674337# a_3405057_686207# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6484 a_3359663_699281# a_3361095_699281# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X6485 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6486 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6487 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6488 a_3403286_704090# a_3381563_702505# w_3403067_702950# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6489 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6490 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6491 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6492 w_3403067_716474# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6493 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6494 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6495 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6496 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6497 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6498 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6499 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6500 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6501 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6502 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6503 w_3185490_798160# a_3403286_716870# a_3403286_717614# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6504 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6505 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6506 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6507 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6508 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6509 a_3403286_717614# a_3403189_717414# w_3403067_716474# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6510 w_3263498_541854# a_3400801_715182# a_3400801_715182# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6511 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6512 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6513 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6514 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6515 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6516 a_3400801_701658# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6517 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6518 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6519 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6520 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6521 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6522 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6523 a_3400801_701658# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6524 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6525 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6526 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6527 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6528 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6529 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6530 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6531 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6532 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6533 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6534 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6535 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6536 a_3403286_703346# a_3403001_700774# w_3403067_702950# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6537 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6538 v2 a_3439418_744112# a_3443016_749796# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6539 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6540 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6541 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6542 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6543 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6544 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6545 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6546 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6547 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6548 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6549 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6550 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6551 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6552 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6553 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6554 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6555 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6556 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6557 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6558 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6559 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6560 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6561 v2 a_3439418_744112# a_3443016_749796# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6562 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6563 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6564 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6565 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6566 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6567 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6568 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6569 w_3403067_716474# a_3381563_702505# a_3403286_716870# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6570 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6571 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6572 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6573 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6574 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6575 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6576 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X6577 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6578 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6579 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6580 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6581 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6582 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6583 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6584 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6585 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6586 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6587 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6588 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6589 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6590 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6591 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6592 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6593 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6594 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6595 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6596 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6597 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6598 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6599 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6600 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6601 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6602 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6603 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6604 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6605 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6606 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6607 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6608 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6609 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6610 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6611 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6612 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6613 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6614 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6615 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6616 w_3381441_717637# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6617 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6618 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6619 a_3443016_749796# a_3439418_744112# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6620 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6621 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6622 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6623 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6624 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6625 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6626 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6627 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6628 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6629 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6630 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6631 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6632 w_3263498_541854# a_3379175_700273# w_3381441_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6633 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6634 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6635 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6636 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6637 a_3401256_686207# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6638 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6639 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6640 v2 a_3366260_744206# a_3369760_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6641 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6642 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6643 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6644 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6645 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6646 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6647 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6648 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6649 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6650 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6651 a_3440844_744112# a_3420382_721009# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6652 w_3403067_702950# a_3403001_700774# a_3403286_703346# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6653 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6654 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6655 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6656 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6657 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6658 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6659 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6660 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6661 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6662 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6663 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6664 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6665 a_3381660_718777# a_3381660_718033# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6666 a_3366286_744142# a_3366260_744112# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6667 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6668 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6669 w_3263498_541854# a_3405057_686207# w_3407323_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6670 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6671 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6672 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6673 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6674 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6675 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6676 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6677 a_3422243_697443# a_3420381_704937# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X6678 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6679 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6680 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6681 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6682 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6683 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6684 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6685 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6686 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6687 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6688 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6689 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6690 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6691 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6692 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6693 a_3401256_686207# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6694 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6695 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6696 a_3361095_699281# a_3379272_706425# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X6697 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6698 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6699 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6700 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6701 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6702 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6703 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6704 a_3420294_720809# a_3420381_704937# w_3422394_717637# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6705 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6706 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6707 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6708 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6709 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6710 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6711 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6712 a_3403286_703346# a_3403001_700774# w_3403067_702950# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6713 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6714 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6715 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6716 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6717 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6718 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6719 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6720 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6721 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6722 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6723 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6724 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6725 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6726 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6727 a_3394410_690671# a_3398102_692829# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=500000u
X6728 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6729 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6730 v2 a_3359810_749958# a_3335479_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6731 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6732 a_3403286_717614# a_3403189_717414# w_3403067_716474# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6733 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6734 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6735 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6736 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6737 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6738 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6739 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6740 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6741 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6742 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6743 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6744 v2 a_3434368_749958# a_3428294_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6745 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6746 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6747 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6748 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6749 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6750 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6751 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6752 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6753 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6754 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6755 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6756 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6757 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6758 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6759 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6760 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6761 a_3359663_699917# a_3361095_699599# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X6762 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6763 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6764 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6765 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6766 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6767 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6768 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6769 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6770 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6771 a_3381660_701961# a_3361095_699281# w_3381441_701565# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6772 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6773 a_3369760_754598# a_3366260_744206# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6774 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6775 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6776 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6777 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6778 a_3335479_772599# a_3359810_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6779 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6780 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6781 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6782 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6783 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6784 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6785 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6786 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6787 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6788 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6789 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6790 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6791 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6792 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6793 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6794 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6795 w_3263498_541854# a_3379175_716345# a_3379175_716345# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6796 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6797 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6798 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6799 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6800 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6801 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6802 w_3263498_541854# a_3408579_674425# w_3422394_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6803 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6804 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6805 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6806 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6807 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6808 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6809 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6810 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6811 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6812 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6813 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6814 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6815 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6816 w_3422394_717637# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6817 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6818 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6819 w_3263498_541854# a_3400801_715182# w_3403067_716474# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6820 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6821 w_3185490_798160# a_3403286_716870# a_3403286_716870# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6822 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6823 a_3335479_772599# a_3359810_749958# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6824 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6825 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6826 a_3446663_700235# a_3448095_700553# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X6827 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6828 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6829 w_3403067_702950# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6830 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6831 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6832 a_3379175_716345# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6833 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6834 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6835 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6836 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6837 w_3263498_541854# a_3407435_674425# w_3422393_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6838 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6839 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6840 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6841 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6842 a_3428294_754598# a_3434368_749958# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6843 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6844 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6845 w_3185490_798160# a_3403286_716870# a_3403286_717614# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6846 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6847 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6848 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6849 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6850 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6851 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6852 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6853 w_3185490_798160# a_3403286_703346# a_3403286_703346# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6854 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6855 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6856 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6857 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6858 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X6859 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6860 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6861 w_3263498_541854# a_3401256_686207# w_3396510_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6862 a_3369760_754598# a_3366260_744206# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6863 a_3335479_772599# a_3359810_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6864 a_3443016_749796# a_3439418_744112# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6865 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6866 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6867 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6868 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6869 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6870 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6871 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6872 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6873 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6874 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6875 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6876 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6877 w_3396510_687499# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6878 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6879 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6880 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6881 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6882 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6883 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6884 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6885 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6886 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6887 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6888 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6889 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6890 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6891 a_3408579_674425# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6892 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6893 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6894 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6895 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6896 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6897 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6898 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6899 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6900 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6901 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6902 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6903 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6904 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6905 a_3434368_749958# a_3435992_747994# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6906 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6907 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6908 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6909 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6910 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6911 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6912 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6913 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6914 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6915 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6916 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6917 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6918 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6919 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6920 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6921 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6922 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6923 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6924 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6925 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6926 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6927 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6928 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6929 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6930 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6931 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6932 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6933 a_3381660_718033# a_3381563_717833# w_3381441_717637# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6934 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6935 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6936 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6937 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6938 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6939 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6940 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6941 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6942 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6943 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6944 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6945 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6946 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6947 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6948 a_3422243_697443# a_3420381_704937# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X6949 a_3401256_686207# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6950 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6951 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6952 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6953 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6954 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6955 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6956 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6957 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6958 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6959 w_3185490_798160# a_3366260_744206# a_3369760_754598# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6960 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6961 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6962 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X6963 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6964 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6965 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6966 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6967 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6968 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6969 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6970 w_3263498_541854# a_3407435_674425# w_3422393_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6971 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6972 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6973 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6974 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6975 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6976 a_3403286_703346# a_3403286_703346# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6977 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6978 w_3263498_541854# a_3405057_686207# w_3407323_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6979 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6980 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6981 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6982 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6983 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6984 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6985 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6986 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6987 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6988 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6989 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6990 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6991 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6992 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6993 w_3185490_798160# a_3399027_674337# a_3405057_686207# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6994 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6995 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6996 w_3407323_687499# a_3407282_686697# a_3407542_687895# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6997 a_3362906_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X6998 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6999 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7000 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7001 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7002 a_3361095_699281# a_3379272_706425# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X7003 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7004 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7005 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7006 a_3403286_704090# a_3403286_703346# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7007 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7008 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7009 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7010 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7011 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7012 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7013 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7014 w_3185490_798160# a_3420293_701761# a_3420293_704737# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7015 w_3185490_798160# a_3381660_701961# a_3381660_702705# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7016 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7017 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7018 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7019 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7020 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X7021 a_3362906_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X7022 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7023 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7024 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7025 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7026 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7027 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7028 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7029 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7030 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7031 w_3263498_541854# a_3379175_716345# w_3381441_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7032 a_3420971_697443# a_3420653_698875# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X7033 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7034 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7035 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7036 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7037 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7038 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7039 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7040 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7041 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7042 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7043 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
R7 a_3427310_772647# m3_3612250_970254# sky130_fd_pr__res_generic_m3 w=2.505e+07u l=4.15e+06u
X7044 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7045 w_3263498_541854# a_3379175_716345# a_3379175_716345# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7046 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7047 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7048 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7049 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7050 a_3403286_716870# a_3381563_702505# w_3403067_716474# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7051 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7052 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7053 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7054 w_3263498_541854# a_3400801_715182# a_3400801_715182# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7055 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7056 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7057 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X7058 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7059 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7060 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7061 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7062 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7063 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7064 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7065 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7066 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7067 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7068 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7069 a_3400801_701658# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7070 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7071 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7072 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7073 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7074 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7075 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7076 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7077 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7078 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7079 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7080 w_3407323_687499# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7081 w_3185490_798160# a_3394410_687695# a_3394410_687695# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7082 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7083 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7084 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7085 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7086 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7087 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7088 w_3185490_798160# a_3403286_716870# a_3403286_716870# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7089 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7090 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7091 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7092 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7093 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7094 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7095 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7096 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7097 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7098 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7099 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7100 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7101 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7102 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7103 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7104 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7105 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7106 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7107 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7108 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7109 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7110 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7111 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7112 w_3263498_541854# a_3408579_674425# w_3422394_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7113 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7114 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7115 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7116 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7117 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7118 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7119 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7120 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7121 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7122 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7123 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7124 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7125 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7126 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7127 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7128 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7129 a_3400801_715182# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7130 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7131 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7132 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7133 a_3407542_688639# a_3407542_687895# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7134 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7135 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7136 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7137 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7138 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7139 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7140 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7141 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7142 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7143 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7144 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7145 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7146 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7147 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7148 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7149 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7150 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7151 w_3381441_717637# a_3381563_717833# a_3381660_718033# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7152 a_3428294_754598# a_3434368_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7153 w_3185490_798160# a_3399027_674337# a_3407435_674425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X7154 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7155 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7156 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7157 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7158 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7159 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7160 a_3381660_718777# a_3379272_706425# w_3381441_717637# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7161 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7162 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X7163 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7164 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7165 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7166 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7167 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7168 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7169 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7170 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7171 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7172 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7173 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7174 w_3396510_687499# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7175 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7176 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7177 a_3400801_701658# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X7178 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7179 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7180 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7181 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7182 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7183 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7184 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7185 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7186 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7187 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7188 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7189 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7190 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7191 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7192 a_3361095_699281# a_3379272_706425# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X7193 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7194 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7195 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7196 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7197 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7198 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7199 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7200 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7201 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7202 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7203 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7204 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7205 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7206 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7207 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7208 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7209 w_3185490_798160# a_3399027_674337# a_3401256_686207# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X7210 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7211 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7212 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7213 a_3403286_703346# a_3403286_703346# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7214 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7215 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7216 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7217 a_3399027_674337# w_3474538_503344# sky130_fd_pr__diode_pd2nw_05v5 area=2.25e+16p
X7218 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7219 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7220 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7221 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7222 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7223 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7224 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7225 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7226 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7227 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7228 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7229 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7230 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7231 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7232 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7233 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7234 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7235 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7236 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7237 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7238 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7239 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7240 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7241 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7242 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7243 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7244 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7245 w_3263498_541854# a_3379175_716345# w_3381441_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7246 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7247 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7248 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7249 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7250 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7251 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7252 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7253 w_3263498_541854# a_3379175_700273# w_3381441_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7254 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7255 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7256 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7257 a_3420294_717833# a_3420294_717833# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7258 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7259 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7260 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7261 v2 a_3434368_749958# a_3428294_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7262 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7263 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7264 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7265 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7266 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7267 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7268 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7269 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7270 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7271 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7272 w_3403067_702950# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7273 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7274 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7275 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7276 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7277 w_3407323_687499# a_3381563_702505# a_3407542_688639# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7278 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7279 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7280 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7281 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7282 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7283 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7284 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7285 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7286 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7287 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7288 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7289 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7290 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7291 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7292 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7293 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7294 w_3185490_798160# a_3420293_701761# a_3420293_701761# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7295 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7296 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7297 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7298 w_3185490_798160# a_3381660_701961# a_3381660_701961# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7299 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7300 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7301 a_3379175_716345# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X7302 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7303 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7304 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7305 a_3383521_705357# a_3379272_706425# sky130_fd_pr__cap_mim_m3_1 l=1.4e+07u w=3e+07u
X7306 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7307 w_3263498_541854# a_3379175_716345# a_3379175_716345# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7308 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7309 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7310 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7311 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7312 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7313 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7314 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7315 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7316 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7317 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7318 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7319 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7320 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7321 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7322 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7323 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7324 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7325 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7326 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7327 w_3185490_798160# a_3403286_716870# a_3403286_717614# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7328 w_3403067_716474# a_3403189_717414# a_3403286_717614# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7329 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7330 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7331 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7332 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7333 a_3407435_674425# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X7334 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7335 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7336 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7337 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7338 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7339 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7340 a_3369760_754598# a_3366260_744206# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7341 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7342 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7343 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7344 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7345 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7346 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7347 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7348 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7349 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7350 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7351 w_3185490_798160# a_3394410_687695# a_3394410_690671# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7352 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7353 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7354 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7355 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7356 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7357 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7358 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7359 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7360 a_3443016_749796# a_3439418_744112# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7361 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7362 w_3185490_798160# a_3399027_674337# a_3399027_674337# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X7363 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7364 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7365 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7366 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7367 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7368 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7369 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7370 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7371 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7372 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7373 a_3381660_702705# a_3381660_701961# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7374 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7375 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7376 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7377 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7378 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7379 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7380 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7381 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7382 w_3185490_798160# a_3403286_703346# a_3403286_704090# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7383 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7384 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7385 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7386 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7387 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7388 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7389 a_3420294_717833# a_3381563_717833# w_3422394_717637# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7390 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7391 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7392 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7393 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7394 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7395 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7396 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7397 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7398 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7399 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X7400 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7401 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7402 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7403 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7404 v2 a_3439418_744112# a_3443016_749796# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7405 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7406 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7407 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7408 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7409 w_3381441_701565# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7410 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7411 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7412 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7413 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7414 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7415 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7416 w_3185490_798160# a_3381660_718033# a_3381660_718777# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7417 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7418 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7419 a_3381660_718033# a_3381660_718033# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7420 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7421 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7422 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7423 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7424 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7425 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7426 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7427 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7428 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7429 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7430 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7431 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7432 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7433 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7434 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7435 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7436 a_3401256_686207# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7437 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7438 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7439 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7440 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7441 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7442 a_3381660_702705# a_3381563_702505# w_3381441_701565# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7443 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7444 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7445 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7446 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7447 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7448 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7449 w_3263498_541854# a_3407435_674425# w_3422393_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7450 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7451 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7452 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7453 a_3403286_704090# a_3403286_703346# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7454 w_3263498_541854# a_3405057_686207# w_3407323_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7455 w_3403067_702950# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7456 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7457 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7458 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7459 a_3394410_690671# a_3263636_541992# w_3396510_687499# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7460 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7461 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7462 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7463 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7464 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7465 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7466 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7467 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7468 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7469 w_3185490_798160# a_3394410_687695# a_3394410_687695# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7470 w_3407323_687499# a_3381563_702505# a_3407542_688639# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7471 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7472 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7473 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7474 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7475 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7476 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7477 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7478 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7479 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7480 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7481 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7482 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7483 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7484 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7485 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7486 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7487 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7488 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7489 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7490 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7491 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7492 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7493 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7494 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7495 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7496 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7497 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7498 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7499 a_3379175_716345# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7500 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7501 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7502 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7503 w_3396510_687499# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7504 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7505 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7506 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7507 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7508 w_3263498_541854# a_3379175_716345# w_3381441_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7509 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7510 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7511 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7512 w_3185490_798160# a_3442918_747574# a_3439418_744112# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7513 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7514 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7515 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7516 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7517 w_3263498_541854# a_3401256_686207# a_3387775_698875# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7518 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7519 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7520 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7521 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7522 w_3263498_541854# a_3379175_716345# a_3379175_716345# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7523 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7524 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7525 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7526 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7527 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7528 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7529 w_3185490_798160# a_3403286_716870# a_3403286_716870# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7530 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7531 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7532 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7533 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7534 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7535 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7536 a_3400801_701658# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7537 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7538 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7539 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7540 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7541 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7542 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7543 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7544 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7545 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7546 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7547 w_3185490_798160# a_3394410_687695# a_3394410_690671# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7548 a_3407542_687895# a_3407542_687895# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7549 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7550 v2 a_3366260_744206# a_3369760_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7551 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7552 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7553 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7554 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7555 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7556 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7557 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7558 a_3420294_717833# a_3381563_717833# w_3422394_717637# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7559 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7560 a_3362906_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X7561 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7562 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7563 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7564 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7565 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7566 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7567 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7568 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7569 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7570 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7571 a_3381660_702705# a_3381660_701961# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7572 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7573 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7574 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7575 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7576 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7577 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7578 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7579 w_3263498_541854# a_3408579_674425# w_3422394_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7580 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7581 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7582 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7583 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7584 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7585 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7586 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7587 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7588 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7589 w_3422393_701565# a_3381563_702505# a_3420293_704737# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7590 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7591 a_3362906_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X7592 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7593 w_3422394_717637# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7594 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7595 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7596 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7597 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7598 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7599 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7600 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7601 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7602 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7603 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7604 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7605 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7606 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7607 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7608 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7609 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X7610 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7611 w_3185490_798160# a_3434368_749958# a_3428294_754598# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7612 w_3403067_716474# a_3381563_702505# a_3403286_716870# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7613 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7614 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7615 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7616 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7617 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7618 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7619 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7620 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7621 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7622 a_3407542_688639# a_3381563_702505# w_3407323_687499# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7623 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7624 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7625 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7626 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7627 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7628 w_3381441_701565# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7629 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7630 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7631 a_3361095_699281# a_3379272_706425# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X7632 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7633 v2 a_3359810_749958# a_3335479_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7634 w_3185490_798160# a_3439418_744112# a_3443016_749796# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7635 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7636 a_3394410_690671# a_3263636_541992# w_3396510_687499# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7637 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7638 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7639 w_3263498_541854# a_3401256_686207# w_3396510_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7640 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7641 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7642 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7643 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7644 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7645 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7646 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7647 w_3396510_687499# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7648 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7649 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7650 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7651 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7652 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7653 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7654 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7655 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7656 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7657 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7658 a_3381660_702705# a_3381563_702505# w_3381441_701565# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7659 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7660 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7661 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7662 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7663 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7664 w_3263498_541854# a_3407435_674425# a_3407435_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7665 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7666 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7667 a_3403286_703346# a_3403286_703346# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7668 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7669 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7670 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7671 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7672 w_3403067_702950# a_3381563_702505# a_3403286_704090# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7673 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7674 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7675 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7676 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7677 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7678 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7679 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7680 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7681 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7682 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7683 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7684 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7685 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7686 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7687 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7688 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7689 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7690 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7691 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7692 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7693 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7694 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7695 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7696 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7697 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7698 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7699 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7700 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7701 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X7702 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7703 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7704 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7705 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7706 a_3359810_749958# a_3362834_747994# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7707 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7708 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7709 w_3185490_798160# a_3381660_718033# a_3381660_718033# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7710 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7711 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7712 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7713 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7714 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7715 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7716 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7717 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7718 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7719 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7720 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7721 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7722 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7723 w_3422394_717637# a_3420381_704937# a_3420294_720809# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7724 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7725 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7726 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7727 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7728 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7729 a_3379175_716345# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7730 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7731 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7732 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7733 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7734 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7735 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7736 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7737 w_3263498_541854# a_3407435_674425# w_3422393_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7738 a_3428294_754598# a_3434368_749958# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7739 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7740 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7741 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7742 w_3263498_541854# a_3379175_716345# w_3381441_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7743 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7744 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7745 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7746 w_3263498_541854# a_3379175_700273# w_3381441_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7747 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7748 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7749 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7750 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7751 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7752 a_3386821_697443# a_3387139_698875# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X7753 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7754 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7755 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7756 a_3362906_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X7757 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7758 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7759 w_3185490_798160# a_3407542_687895# a_3407542_687895# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7760 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7761 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7762 a_3403286_703346# a_3403001_700774# w_3403067_702950# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7763 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7764 w_3185490_798160# a_3420294_717833# a_3420294_720809# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7765 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7766 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7767 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7768 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7769 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7770 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7771 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7772 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7773 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7774 w_3185490_798160# a_3394410_687695# a_3394410_690671# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7775 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7776 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7777 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7778 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7779 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7780 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7781 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7782 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7783 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7784 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7785 a_3362906_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X7786 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7787 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7788 w_3185490_798160# a_3399027_674337# a_3379175_716345# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X7789 a_3428294_754598# a_3434368_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7790 a_3366260_744206# a_3369760_747574# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7791 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7792 a_3407435_674425# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X7793 w_3381441_717637# a_3379272_706425# a_3381660_718777# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7794 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7795 w_3185490_798160# a_3420293_701761# a_3420293_704737# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7796 w_3185490_798160# a_3381660_701961# a_3381660_702705# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7797 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7798 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7799 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7800 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7801 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7802 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7803 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7804 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7805 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7806 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7807 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7808 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7809 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7810 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7811 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7812 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7813 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7814 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7815 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7816 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7817 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7818 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7819 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7820 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7821 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7822 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7823 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7824 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7825 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7826 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7827 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7828 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7829 w_3185490_798160# a_3399027_674337# a_3399027_674337# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X7830 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7831 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7832 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7833 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7834 w_3422393_701565# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7835 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7836 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7837 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
R8 m3_3146060_431482# w_3185490_798160# sky130_fd_pr__res_generic_m3 w=7.4e+07u l=2.055e+07u
X7838 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7839 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7840 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7841 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7842 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7843 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7844 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7845 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7846 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7847 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7848 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7849 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7850 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7851 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7852 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7853 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7854 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7855 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7856 a_3405057_686207# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7857 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7858 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7859 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7860 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7861 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7862 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7863 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7864 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7865 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7866 a_3427310_772647# v2 sky130_fd_pr__diode_pd2nw_05v5 area=2.25e+16p
X7867 a_3422243_697443# a_3420381_704937# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X7868 a_3359663_700553# a_3361095_700235# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X7869 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7870 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7871 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7872 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7873 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7874 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7875 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7876 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7877 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7878 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7879 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7880 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7881 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7882 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7883 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7884 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7885 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7886 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X7887 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7888 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7889 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7890 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7891 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7892 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7893 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7894 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7895 w_3185490_798160# a_3403286_703346# a_3403286_703346# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7896 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7897 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7898 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7899 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7900 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7901 w_3422393_701565# a_3422243_697443# a_3420293_701761# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7902 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7903 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7904 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7905 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7906 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7907 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7908 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7909 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7910 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7911 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7912 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7913 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7914 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7915 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7916 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7917 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7918 v2 a_3434368_749958# a_3428294_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7919 w_3422394_717637# a_3420381_704937# a_3420294_720809# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7920 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7921 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7922 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7923 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7924 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7925 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7926 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7927 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7928 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7929 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7930 w_3381441_701565# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7931 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7932 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7933 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7934 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7935 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7936 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7937 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7938 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7939 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7940 w_3185490_798160# a_3381660_718033# a_3381660_718777# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7941 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7942 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7943 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7944 a_3381660_718777# a_3379272_706425# w_3381441_717637# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7945 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7946 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7947 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7948 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7949 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7950 a_3369760_754598# a_3366260_744206# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7951 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7952 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7953 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7954 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7955 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7956 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7957 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7958 a_3335479_772599# a_3359810_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7959 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7960 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7961 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7962 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7963 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7964 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7965 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7966 a_3394410_687695# a_3387775_698875# w_3396510_687499# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7967 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7968 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7969 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7970 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7971 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7972 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7973 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7974 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7975 w_3263498_541854# a_3379175_700273# a_3379175_700273# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7976 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7977 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7978 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7979 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7980 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7981 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7982 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7983 a_3394410_687695# a_3387775_698875# w_3396510_687499# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7984 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X7985 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7986 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7987 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7988 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7989 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7990 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7991 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7992 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7993 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7994 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7995 w_3185490_798160# a_3399027_674337# a_3400801_701658# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X7996 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7997 v2 a_3420382_721009# a_3436064_746854# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7998 w_3185490_798160# a_3394410_687695# a_3394410_690671# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7999 a_3335479_772599# a_3359810_749958# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8000 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8001 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8002 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8003 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8004 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8005 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8006 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8007 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8008 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8009 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8010 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8011 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8012 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8013 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8014 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8015 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8016 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8017 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8018 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8019 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8020 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8021 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8022 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8023 w_3185490_798160# a_3420293_701761# a_3420293_701761# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8024 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8025 w_3185490_798160# a_3381660_701961# a_3381660_701961# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8026 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8027 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8028 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8029 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8030 a_3400801_715182# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X8031 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8032 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8033 a_3379175_716345# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8034 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8035 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8036 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8037 a_3436064_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X8038 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8039 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8040 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8041 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8042 w_3422394_717637# a_3381563_717833# a_3420294_717833# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8043 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8044 a_3369760_754598# a_3366260_744206# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8045 a_3335479_772599# a_3359810_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8046 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8047 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8048 a_3428294_754598# a_3434368_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8049 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8050 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8051 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8052 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8053 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8054 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8055 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8056 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8057 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8058 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8059 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8060 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8061 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8062 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8063 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8064 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8065 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8066 a_3436064_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X8067 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8068 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8069 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8070 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8071 w_3263498_541854# a_3400801_715182# a_3400801_715182# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8072 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8073 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8074 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8075 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8076 a_3400801_701658# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8077 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8078 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8079 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8080 a_3440870_744142# a_3434368_749958# a_3441490_744142# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8081 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8082 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8083 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8084 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8085 w_3407323_687499# a_3407282_686697# a_3407542_687895# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8086 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8087 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8088 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8089 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8090 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8091 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8092 a_3422243_697443# a_3420381_704937# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X8093 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8094 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8095 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8096 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8097 a_3405154_692359# a_3409354_691535# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X8098 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8099 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8100 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8101 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8102 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8103 w_3407323_687499# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8104 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X8105 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8106 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8107 v2 a_3359810_749958# a_3335479_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8108 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8109 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8110 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8111 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8112 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8113 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8114 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8115 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8116 a_3442918_747574# a_3440870_744142# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8117 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8118 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8119 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8120 w_3422394_717637# a_3420381_704937# a_3420294_720809# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8121 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8122 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8123 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8124 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8125 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8126 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8127 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8128 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8129 w_3381441_717637# a_3381563_717833# a_3381660_718033# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8130 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8131 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8132 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8133 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8134 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8135 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8136 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8137 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8138 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8139 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8140 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8141 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8142 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8143 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8144 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8145 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8146 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8147 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8148 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8149 w_3185490_798160# a_3359810_749958# a_3335479_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8150 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8151 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8152 w_3185490_798160# a_3366260_744206# a_3369760_754598# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8153 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8154 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8155 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8156 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8157 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8158 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8159 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8160 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8161 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8162 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8163 a_3407542_687895# a_3407282_686697# w_3407323_687499# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8164 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8165 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8166 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8167 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8168 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8169 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8170 w_3403067_716474# a_3403189_717414# a_3403286_717614# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8171 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8172 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8173 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8174 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8175 a_3379175_700273# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8176 a_3407542_687895# a_3407282_686697# w_3407323_687499# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8177 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8178 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8179 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8180 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8181 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8182 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8183 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8184 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8185 w_3185490_798160# a_3407542_687895# a_3407542_687895# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8186 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8187 w_3381441_701565# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8188 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8189 a_3394410_687695# a_3387775_698875# w_3396510_687499# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8190 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8191 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8192 v2 a_3366260_744206# a_3369760_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8193 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8194 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8195 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8196 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8197 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8198 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8199 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8200 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8201 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8202 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8203 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8204 w_3396510_687499# a_3387775_698875# a_3394410_687695# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8205 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8206 a_3443016_749796# a_3439418_744112# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8207 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8208 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8209 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8210 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8211 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8212 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8213 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8214 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8215 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8216 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8217 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8218 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8219 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8220 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8221 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8222 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8223 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8224 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8225 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8226 w_3263498_541854# a_3407435_674425# a_3407435_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8227 v2 a_3435992_747994# a_3434368_749958# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8228 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8229 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8230 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8231 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8232 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8233 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8234 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8235 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8236 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8237 a_3400801_701658# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8238 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8239 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8240 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8241 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8242 a_3443016_749796# a_3439418_744112# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8243 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8244 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X8245 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8246 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8247 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8248 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8249 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8250 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8251 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8252 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8253 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8254 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8255 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8256 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8257 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8258 w_3263498_541854# a_3405057_686207# w_3407323_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8259 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8260 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8261 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8262 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8263 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8264 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8265 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8266 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8267 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8268 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8269 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8270 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8271 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8272 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8273 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8274 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8275 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8276 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8277 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8278 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8279 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8280 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8281 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8282 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8283 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8284 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8285 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8286 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8287 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8288 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8289 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8290 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8291 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8292 a_3379175_716345# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8293 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8294 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8295 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8296 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8297 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8298 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8299 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8300 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8301 w_3263498_541854# a_3407435_674425# w_3422393_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8302 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8303 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8304 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8305 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8306 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8307 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8308 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8309 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8310 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8311 w_3381441_701565# a_3381563_702505# a_3381660_702705# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8312 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8313 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8314 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8315 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8316 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8317 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8318 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8319 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8320 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8321 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8322 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8323 w_3185490_798160# a_3420293_701761# a_3420293_704737# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8324 a_3403286_704090# a_3381563_702505# w_3403067_702950# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8325 w_3403067_702950# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8326 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8327 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8328 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8329 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8330 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8331 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8332 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8333 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8334 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8335 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8336 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8337 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8338 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8339 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8340 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8341 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8342 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8343 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8344 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8345 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8346 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8347 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8348 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8349 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8350 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8351 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8352 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8353 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8354 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8355 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8356 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8357 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8358 a_3439418_744112# a_3442918_747574# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8359 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8360 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8361 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8362 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8363 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8364 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8365 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8366 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8367 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8368 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8369 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8370 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8371 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8372 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8373 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8374 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8375 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8376 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8377 a_3401256_686207# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8378 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8379 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8380 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8381 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8382 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8383 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8384 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8385 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8386 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8387 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8388 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8389 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8390 w_3263498_541854# a_3379175_716345# a_3379175_716345# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8391 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8392 w_3407323_687499# a_3407282_686697# a_3407542_687895# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8393 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8394 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8395 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8396 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8397 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8398 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8399 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8400 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8401 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8402 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8403 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8404 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8405 a_3381660_701961# a_3381660_701961# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8406 w_3422393_701565# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8407 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8408 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8409 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8410 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8411 w_3403067_716474# a_3381563_702505# a_3403286_716870# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8412 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8413 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8414 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8415 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8416 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8417 w_3407323_687499# a_3381563_702505# a_3407542_688639# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8418 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8419 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8420 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8421 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8422 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8423 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8424 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8425 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8426 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8427 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8428 a_3405057_686207# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8429 a_3379175_700273# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8430 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8431 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8432 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8433 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8434 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8435 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8436 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8437 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8438 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8439 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8440 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8441 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8442 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8443 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8444 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8445 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8446 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8447 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8448 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8449 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8450 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8451 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8452 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8453 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8454 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8455 a_3424227_705357# a_3420381_704937# sky130_fd_pr__cap_mim_m3_1 l=1.4e+07u w=3e+07u
X8456 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8457 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8458 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8459 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8460 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8461 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8462 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8463 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8464 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8465 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8466 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8467 a_3443016_749796# a_3439418_744112# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8468 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8469 a_3367712_744142# a_3366422_743586# a_3368332_744142# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8470 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8471 w_3185490_798160# a_3420294_717833# a_3420294_720809# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8472 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8473 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8474 w_3422393_701565# a_3381563_702505# a_3420293_704737# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8475 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8476 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8477 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8478 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8479 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8480 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8481 a_3420293_704737# a_3420293_701761# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8482 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8483 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8484 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8485 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8486 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8487 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8488 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8489 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8490 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8491 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8492 w_3263498_541854# a_3405057_686207# a_3405057_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8493 a_3443016_749796# a_3439418_744112# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8494 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8495 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8496 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8497 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8498 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8499 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8500 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8501 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8502 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8503 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8504 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8505 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8506 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8507 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8508 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8509 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8510 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8511 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8512 w_3185490_798160# a_3407542_687895# a_3407542_688639# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8513 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8514 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8515 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8516 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8517 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8518 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8519 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8520 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8521 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8522 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8523 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8524 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8525 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8526 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8527 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8528 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8529 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8530 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X8531 a_3420293_701761# a_3420293_701761# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8532 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8533 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8534 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8535 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8536 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8537 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8538 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8539 w_3263498_541854# a_3407435_674425# a_3407435_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8540 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8541 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8542 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8543 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8544 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8545 w_3263498_541854# a_3379175_700273# a_3379175_700273# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8546 w_3422394_717637# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8547 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8548 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8549 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8550 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8551 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8552 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8553 a_3403286_703346# a_3403001_700774# w_3403067_702950# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8554 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8555 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8556 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8557 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8558 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8559 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8560 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8561 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8562 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8563 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8564 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8565 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8566 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8567 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8568 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8569 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8570 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8571 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8572 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8573 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8574 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8575 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8576 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8577 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8578 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8579 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8580 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8581 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8582 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8583 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8584 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8585 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8586 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8587 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8588 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8589 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8590 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8591 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8592 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8593 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8594 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8595 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8596 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8597 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8598 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8599 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8600 w_3185490_798160# a_3394410_687695# a_3394410_687695# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8601 w_3185490_798160# a_3434368_749958# a_3428294_754598# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8602 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8603 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8604 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8605 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8606 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8607 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8608 a_3443016_749796# a_3439418_744112# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8609 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8610 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8611 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8612 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8613 w_3396510_687499# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8614 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8615 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8616 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8617 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8618 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8619 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8620 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8621 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8622 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8623 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8624 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8625 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8626 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8627 w_3263498_541854# a_3379175_716345# a_3379175_716345# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8628 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8629 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8630 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8631 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X8632 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8633 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8634 a_3407435_674425# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8635 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8636 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8637 a_3420293_704737# a_3381563_702505# w_3422393_701565# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8638 w_3381441_701565# a_3361095_699281# a_3381660_701961# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8639 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8640 w_3263498_541854# a_3400801_715182# a_3400801_715182# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8641 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8642 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8643 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8644 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8645 w_3263498_541854# a_3405057_686207# w_3407323_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8646 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8647 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8648 w_3407323_687499# a_3381563_702505# a_3407542_688639# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8649 w_3185490_798160# a_3420293_701761# a_3420293_701761# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8650 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8651 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8652 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8653 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8654 v2 a_3434368_749958# a_3428294_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8655 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8656 v2 a_3435992_747994# a_3434368_749958# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8657 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8658 w_3407323_687499# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8659 a_3407542_688639# a_3407542_687895# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8660 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8661 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8662 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8663 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8664 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8665 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8666 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8667 a_3403286_704090# a_3381563_702505# w_3403067_702950# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8668 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8669 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8670 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8671 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8672 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8673 a_3420294_717833# a_3420294_717833# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8674 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8675 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8676 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8677 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8678 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8679 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8680 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8681 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8682 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8683 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8684 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8685 a_3394410_690671# a_3394410_687695# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8686 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8687 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8688 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8689 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8690 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8691 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8692 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8693 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8694 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8695 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8696 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8697 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8698 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8699 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8700 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8701 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8702 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8703 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8704 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8705 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8706 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8707 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8708 a_3436064_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X8709 w_3422393_701565# a_3422243_697443# a_3420293_701761# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8710 w_3403067_716474# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8711 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8712 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8713 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8714 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8715 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8716 a_3420293_704737# a_3420293_701761# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8717 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8718 a_3405057_686207# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8719 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8720 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8721 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8722 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8723 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8724 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8725 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8726 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8727 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8728 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8729 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8730 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8731 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8732 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8733 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8734 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8735 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8736 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8737 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8738 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X8739 a_3379175_700273# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8740 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8741 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8742 a_3436064_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X8743 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8744 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8745 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8746 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8747 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8748 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8749 v2 a_3439418_744112# a_3443016_749796# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8750 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8751 w_3185490_798160# a_3407542_687895# a_3407542_688639# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8752 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8753 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8754 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8755 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8756 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8757 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8758 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8759 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8760 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8761 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8762 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8763 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8764 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8765 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8766 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8767 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8768 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8769 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8770 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8771 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8772 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8773 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8774 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8775 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8776 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8777 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8778 a_3381660_718033# a_3381563_717833# w_3381441_717637# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8779 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8780 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8781 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8782 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8783 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8784 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8785 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8786 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8787 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8788 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8789 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8790 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8791 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8792 a_3428294_754598# a_3434368_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8793 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8794 a_3400801_701658# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8795 a_3381660_718033# a_3381660_718033# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8796 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8797 w_3185490_798160# a_3420294_717833# a_3420294_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8798 w_3263498_541854# a_3408579_674425# a_3420382_721009# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8799 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8800 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8801 w_3422394_717637# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8802 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8803 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8804 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8805 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8806 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8807 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8808 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8809 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8810 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8811 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8812 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8813 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8814 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8815 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8816 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8817 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8818 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8819 v2 a_3366260_744206# a_3369760_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8820 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8821 a_3420293_704737# a_3381563_702505# w_3422393_701565# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8822 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8823 v2 a_3359810_749958# a_3335479_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8824 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8825 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8826 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8827 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8828 a_3435992_747994# a_3436064_746854# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8829 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8830 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8831 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X8832 a_3399027_674337# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X8833 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8834 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8835 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8836 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8837 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8838 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8839 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8840 w_3263498_541854# a_3400801_701658# a_3400801_701658# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8841 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8842 a_3403286_704090# a_3381563_702505# w_3403067_702950# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8843 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8844 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8845 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8846 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8847 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8848 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8849 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8850 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8851 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8852 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8853 w_3185490_798160# a_3359810_749958# a_3335479_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8854 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8855 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8856 a_3420293_704737# a_3381563_702505# w_3422393_701565# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8857 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8858 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8859 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8860 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8861 a_3403286_716870# a_3381563_702505# w_3403067_716474# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8862 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8863 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8864 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8865 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8866 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8867 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8868 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8869 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8870 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8871 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8872 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8873 w_3185490_798160# a_3399027_674337# a_3379175_700273# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X8874 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8875 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8876 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8877 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8878 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8879 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8880 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8881 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8882 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8883 a_3381660_718033# a_3381563_717833# w_3381441_717637# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8884 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8885 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8886 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8887 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8888 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8889 w_3185490_798160# a_3420294_717833# a_3420294_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8890 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8891 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8892 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8893 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8894 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8895 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8896 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8897 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8898 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8899 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8900 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8901 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8902 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8903 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8904 a_3420294_720809# a_3420294_717833# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8905 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8906 a_3436064_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X8907 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8908 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8909 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8910 v2 a_3366260_744206# a_3369760_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8911 v2 a_3359810_749958# a_3335479_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8912 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8913 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8914 v2 a_3434368_749958# a_3428294_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8915 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8916 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8917 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8918 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8919 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8920 w_3185490_798160# a_3394410_687695# a_3394410_690671# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8921 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8922 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8923 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8924 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8925 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8926 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8927 a_3401256_686207# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8928 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8929 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8930 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8931 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8932 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8933 a_3400801_715182# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8934 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8935 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8936 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8937 a_3436064_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X8938 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8939 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8940 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8941 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8942 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8943 a_3381660_702705# a_3381660_701961# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8944 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8945 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8946 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8947 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8948 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8949 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8950 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8951 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8952 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8953 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8954 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8955 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8956 a_3335479_772599# a_3359810_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8957 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8958 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8959 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8960 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8961 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8962 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8963 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8964 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8965 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8966 a_3362906_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X8967 a_3379175_700273# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8968 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8969 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8970 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8971 a_3379175_716345# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8972 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8973 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8974 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8975 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8976 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8977 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8978 w_3381441_717637# a_3381563_717833# a_3381660_718033# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8979 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8980 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8981 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8982 a_3335479_772599# a_3359810_749958# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8983 a_3381660_718777# a_3379272_706425# w_3381441_717637# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8984 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8985 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8986 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8987 a_3362906_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X8988 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8989 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8990 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8991 a_3409645_692829# a_3407542_688639# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=500000u
X8992 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8993 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8994 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8995 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8996 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8997 w_3185490_798160# a_3399027_674337# sky130_fd_pr__diode_pw2nd_05v5 area=2.25e+16p
X8998 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8999 w_3685938_617428# w_3685938_581428# sky130_fd_pr__diode_pd2nw_05v5 area=2.25e+16p
X9000 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9001 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9002 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9003 a_3428294_754598# a_3434368_749958# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9004 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9005 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9006 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9007 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9008 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9009 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9010 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9011 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9012 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9013 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9014 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9015 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9016 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9017 a_3369760_754598# a_3366260_744206# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9018 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9019 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9020 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9021 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9022 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9023 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9024 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9025 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9026 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9027 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9028 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9029 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9030 a_3420293_704737# a_3381563_702505# w_3422393_701565# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9031 w_3381441_701565# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9032 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9033 v2 a_3439418_744112# a_3443016_749796# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9034 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9035 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9036 w_3185490_798160# a_3399027_674337# a_3400801_715182# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X9037 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9038 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9039 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9040 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9041 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9042 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9043 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9044 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9045 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9046 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9047 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9048 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9049 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9050 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9051 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9052 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9053 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9054 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9055 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9056 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9057 a_3434368_749958# a_3435992_747994# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9058 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9059 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9060 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9061 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9062 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9063 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9064 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9065 w_3263498_541854# a_3407435_674425# a_3407435_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9066 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9067 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9068 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9069 v2 a_3439418_744112# a_3443016_749796# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9070 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9071 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9072 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9073 a_3404909_699542# a_3400898_721334# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X9074 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9075 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9076 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9077 a_3394410_690671# a_3263636_541992# w_3396510_687499# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9078 a_3379175_700273# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X9079 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9080 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9081 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9082 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9083 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9084 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9085 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9086 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9087 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9088 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9089 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9090 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9091 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9092 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9093 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9094 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9095 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9096 w_3263498_541854# a_3405057_686207# w_3407323_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9097 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9098 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9099 w_3403067_702950# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9100 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9101 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9102 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9103 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9104 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9105 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9106 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9107 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9108 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9109 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X9110 v2 a_3362834_747994# a_3359810_749958# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9111 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9112 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9113 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9114 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9115 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9116 w_3185490_798160# a_3399027_674337# a_3408579_674425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X9117 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9118 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9119 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9120 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9121 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9122 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9123 w_3263498_541854# a_3401256_686207# w_3396510_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9124 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9125 w_3185490_798160# a_3394410_687695# a_3394410_690671# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9126 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9127 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9128 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9129 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9130 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9131 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9132 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9133 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9134 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9135 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9136 w_3396510_687499# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9137 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9138 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9139 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9140 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9141 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9142 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9143 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9144 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9145 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9146 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9147 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9148 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9149 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9150 a_3405057_686207# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X9151 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9152 a_3381660_702705# a_3381660_701961# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9153 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9154 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9155 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9156 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9157 a_3381660_701961# a_3381660_701961# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9158 a_3407435_674425# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9159 w_3381441_701565# a_3381563_702505# a_3381660_702705# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9160 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9161 a_3446663_700235# a_3448095_699917# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X9162 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9163 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9164 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9165 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9166 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9167 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9168 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9169 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9170 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9171 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9172 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9173 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9174 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9175 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9176 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9177 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9178 w_3185490_798160# a_3420293_701761# a_3420293_704737# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9179 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9180 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9181 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9182 w_3263498_541854# a_3379175_716345# w_3381441_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9183 w_3185490_798160# a_3442918_747574# a_3439418_744112# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9184 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9185 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9186 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9187 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9188 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9189 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9190 v2 a_3369760_747574# a_3366260_744206# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9191 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9192 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9193 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9194 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9195 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9196 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9197 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9198 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9199 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9200 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9201 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9202 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9203 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9204 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9205 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9206 a_3394410_687695# a_3394410_687695# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9207 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9208 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9209 a_3408579_674425# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X9210 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9211 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9212 w_3263498_541854# a_3401256_686207# a_3401256_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9213 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9214 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9215 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9216 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9217 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9218 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9219 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9220 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9221 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9222 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9223 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9224 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9225 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9226 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9227 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9228 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9229 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9230 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9231 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9232 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9233 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X9234 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9235 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9236 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9237 w_3185490_798160# a_3381660_718777# a_3366422_743586# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9238 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9239 w_3396510_687499# a_3387775_698875# a_3394410_687695# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9240 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9241 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9242 a_3405057_686207# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9243 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9244 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9245 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9246 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9247 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9248 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9249 a_3407542_688639# a_3381563_702505# w_3407323_687499# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9250 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9251 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9252 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9253 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9254 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9255 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9256 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9257 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9258 w_3185490_798160# a_3403286_716870# a_3403286_717614# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9259 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9260 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9261 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9262 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9263 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9264 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9265 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9266 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9267 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9268 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9269 a_3369760_754598# a_3366260_744206# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9270 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9271 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9272 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9273 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9274 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9275 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9276 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9277 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9278 w_3381441_701565# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9279 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9280 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9281 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9282 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9283 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9284 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9285 w_3185490_798160# a_3439418_744112# a_3443016_749796# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9286 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9287 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9288 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9289 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9290 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9291 a_3420293_701761# a_3420293_701761# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9292 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9293 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9294 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9295 w_3263498_541854# a_3408579_674425# a_3408579_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9296 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9297 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9298 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9299 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9300 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9301 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9302 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9303 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9304 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9305 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9306 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9307 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9308 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9309 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9310 a_3408579_674425# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9311 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9312 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9313 w_3185490_798160# a_3439418_744112# a_3443016_749796# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9314 a_3428294_754598# a_3434368_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9315 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9316 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9317 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9318 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9319 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9320 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9321 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9322 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9323 w_3263498_541854# a_3407435_674425# a_3407435_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9324 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9325 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9326 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9327 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9328 w_3263498_541854# a_3405057_686207# a_3405057_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9329 w_3185490_798160# a_3381660_718033# a_3381660_718777# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9330 a_3381660_702705# a_3381563_702505# w_3381441_701565# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9331 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9332 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9333 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9334 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9335 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9336 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9337 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9338 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9339 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9340 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X9341 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9342 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9343 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9344 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9345 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9346 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9347 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9348 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9349 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9350 a_3403286_704090# a_3403286_703346# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9351 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9352 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9353 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9354 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9355 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9356 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9357 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9358 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9359 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9360 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9361 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9362 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9363 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9364 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9365 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9366 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9367 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9368 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9369 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9370 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9371 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9372 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9373 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9374 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9375 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9376 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9377 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9378 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9379 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9380 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9381 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9382 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9383 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9384 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9385 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9386 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9387 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9388 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9389 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9390 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9391 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9392 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9393 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9394 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9395 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9396 a_3400801_715182# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9397 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9398 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9399 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9400 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9401 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9402 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9403 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9404 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9405 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9406 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9407 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9408 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9409 w_3381441_701565# a_3361095_699281# a_3381660_701961# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9410 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9411 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9412 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9413 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9414 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9415 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9416 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9417 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9418 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9419 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9420 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9421 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9422 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9423 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9424 w_3185490_798160# a_3285528_930602# sky130_fd_pr__diode_pw2nd_05v5 area=2.25e+16p
X9425 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9426 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9427 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9428 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9429 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9430 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9431 w_3185490_798160# a_3420293_701761# a_3420293_701761# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9432 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9433 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9434 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9435 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9436 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9437 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9438 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9439 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9440 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9441 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9442 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9443 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9444 w_3381441_717637# a_3379272_706425# a_3381660_718777# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9445 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9446 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9447 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9448 v2 a_3439418_744112# a_3443016_749796# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9449 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9450 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9451 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9452 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9453 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9454 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9455 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9456 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9457 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X9458 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9459 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9460 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9461 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9462 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9463 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9464 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9465 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9466 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9467 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9468 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9469 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9470 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9471 a_3439444_744142# a_3439418_744112# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9472 a_3403001_700774# a_3381563_717833# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X9473 a_3405532_706743# a_3381563_717833# sky130_fd_pr__cap_mim_m3_1 l=2.7e+07u w=1.8e+07u
X9474 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9475 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9476 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9477 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9478 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9479 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9480 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9481 w_3263498_541854# a_3408579_674425# a_3408579_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9482 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9483 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9484 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9485 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9486 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9487 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9488 a_3400801_715182# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9489 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9490 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9491 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9492 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9493 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9494 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9495 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9496 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9497 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9498 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9499 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9500 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9501 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9502 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9503 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9504 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9505 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9506 w_3422393_701565# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9507 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9508 a_3403189_717414# a_3381563_717833# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X9509 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9510 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9511 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9512 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9513 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9514 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9515 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9516 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9517 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9518 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9519 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9520 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9521 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9522 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9523 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9524 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9525 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9526 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9527 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9528 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9529 w_3263498_541854# a_3401256_686207# a_3401256_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9530 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9531 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9532 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9533 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9534 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9535 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9536 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9537 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9538 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9539 v2 a_3362834_747994# a_3359810_749958# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9540 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9541 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9542 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9543 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9544 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9545 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9546 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9547 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9548 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9549 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9550 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9551 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9552 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9553 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9554 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9555 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9556 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9557 a_3405057_686207# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9558 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9559 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9560 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9561 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9562 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9563 w_3185490_798160# a_3399027_674337# a_3400801_715182# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X9564 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9565 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9566 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9567 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9568 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9569 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9570 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9571 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9572 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9573 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9574 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9575 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9576 w_3396510_687499# a_3263636_541992# a_3394410_690671# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9577 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9578 a_3436064_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X9579 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9580 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9581 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9582 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9583 w_3407323_687499# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9584 a_3381660_702705# a_3381563_702505# w_3381441_701565# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9585 a_3443016_749796# a_3439418_744112# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9586 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9587 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9588 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9589 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9590 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9591 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9592 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9593 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9594 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9595 a_3403286_717614# a_3403189_717414# w_3403067_716474# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9596 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9597 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9598 w_3263498_541854# a_3405057_686207# a_3405057_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9599 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9600 w_3185490_798160# a_3420294_717833# a_3420294_720809# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9601 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9602 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9603 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9604 a_3379175_700273# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X9605 w_3185490_798160# a_3403286_716870# a_3403286_716870# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9606 w_3381441_701565# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9607 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9608 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9609 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9610 a_3436064_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X9611 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9612 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9613 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9614 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9615 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9616 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9617 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9618 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9619 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9620 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9621 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9622 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9623 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9624 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9625 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9626 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9627 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9628 v2 a_3369760_747574# a_3366260_744206# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9629 v2 a_3434368_749958# a_3428294_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9630 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9631 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9632 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9633 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9634 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9635 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9636 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9637 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9638 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9639 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9640 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9641 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9642 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9643 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9644 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9645 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9646 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9647 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9648 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9649 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X9650 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9651 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9652 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9653 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9654 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9655 w_3422394_717637# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9656 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9657 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9658 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9659 w_3263498_541854# a_3379175_700273# a_3379175_700273# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9660 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9661 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9662 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9663 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9664 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9665 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9666 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9667 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9668 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9669 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9670 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9671 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9672 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9673 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9674 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9675 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9676 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9677 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9678 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9679 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9680 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9681 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9682 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9683 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9684 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9685 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9686 w_3422393_701565# a_3381563_702505# a_3420293_704737# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9687 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9688 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9689 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9690 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9691 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9692 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9693 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9694 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9695 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9696 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9697 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9698 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9699 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9700 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9701 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9702 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9703 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9704 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9705 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9706 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9707 w_3263498_541854# a_3408579_674425# w_3422394_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9708 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9709 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9710 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9711 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9712 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9713 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9714 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9715 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9716 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9717 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9718 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9719 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9720 w_3263498_541854# a_3400801_701658# w_3403067_702950# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9721 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9722 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9723 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9724 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9725 a_3362834_747994# a_3362906_746854# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9726 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9727 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9728 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9729 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9730 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9731 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9732 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9733 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9734 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9735 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9736 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9737 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9738 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9739 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X9740 w_3403067_702950# a_3403001_700774# a_3403286_703346# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9741 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9742 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X9743 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9744 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9745 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9746 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9747 a_3403286_703346# a_3403286_703346# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9748 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9749 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9750 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9751 w_3263498_541854# a_3379175_716345# w_3381441_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9752 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9753 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9754 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9755 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9756 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9757 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9758 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9759 w_3381441_717637# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9760 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9761 a_3401256_686207# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X9762 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9763 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9764 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9765 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9766 a_3420294_720809# a_3420294_717833# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9767 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9768 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9769 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9770 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9771 a_3403286_717614# a_3403189_717414# w_3403067_716474# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9772 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9773 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9774 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9775 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9776 a_3381660_701961# a_3381660_701961# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9777 w_3185490_798160# a_3381660_718033# a_3381660_718777# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9778 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9779 w_3185628_906308# w_3185628_870308# sky130_fd_pr__diode_pd2nw_05v5 area=2.25e+16p
X9780 w_3185490_798160# a_3407542_687895# a_3407542_687895# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9781 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9782 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9783 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9784 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9785 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9786 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9787 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9788 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9789 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9790 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9791 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9792 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9793 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9794 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9795 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9796 w_3403067_716474# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9797 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9798 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9799 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X9800 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9801 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9802 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9803 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9804 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9805 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9806 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9807 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9808 v2 a_3359810_749958# a_3335479_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9809 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9810 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9811 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9812 w_3396510_687499# a_3263636_541992# a_3394410_690671# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9813 w_3403067_716474# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9814 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9815 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9816 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9817 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9818 a_3369760_747574# a_3367712_744142# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9819 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9820 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9821 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9822 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9823 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9824 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9825 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9826 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9827 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9828 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9829 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9830 a_3403286_717614# a_3403189_717414# w_3403067_716474# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9831 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9832 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9833 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9834 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9835 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9836 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9837 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9838 w_3422394_717637# a_3420381_704937# a_3420294_720809# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9839 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X9840 a_3379175_700273# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9841 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9842 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9843 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9844 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9845 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9846 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9847 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9848 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9849 w_3185490_798160# a_3359810_749958# a_3335479_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9850 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9851 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9852 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9853 w_3381441_701565# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9854 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9855 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9856 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9857 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9858 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X9859 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9860 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9861 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9862 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9863 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9864 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9865 w_3185490_798160# a_3434368_749958# a_3428294_754598# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9866 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9867 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9868 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9869 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9870 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9871 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9872 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9873 a_3381660_718777# a_3379272_706425# w_3381441_717637# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9874 w_3185490_798160# a_3403286_704090# a_3381563_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9875 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9876 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9877 a_3434368_749958# a_3435992_747994# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9878 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9879 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9880 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9881 a_3381660_701961# a_3361095_699281# w_3381441_701565# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9882 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9883 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9884 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9885 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9886 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9887 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9888 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9889 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9890 w_3263498_541854# a_3407435_674425# a_3407435_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9891 a_3381563_717833# a_3403286_704090# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9892 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9893 a_3403286_704090# a_3403286_703346# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9894 v2 a_3366260_744206# a_3369760_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9895 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9896 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9897 a_3400801_701658# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9898 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9899 a_3394410_687695# a_3387775_698875# w_3396510_687499# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9900 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9901 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9902 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9903 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9904 a_3362906_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X9905 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9906 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9907 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9908 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9909 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9910 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9911 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9912 w_3185490_798160# a_3420294_717833# a_3420294_717833# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9913 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9914 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9915 v2 a_3435992_747994# a_3434368_749958# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9916 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9917 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9918 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9919 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9920 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9921 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9922 w_3403067_702950# a_3403001_700774# a_3403286_703346# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9923 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9924 a_3443016_749796# a_3439418_744112# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9925 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9926 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9927 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9928 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9929 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9930 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9931 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9932 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9933 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9934 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9935 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9936 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9937 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9938 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9939 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9940 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9941 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9942 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9943 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9944 w_3263498_541854# a_3400801_701658# a_3400801_701658# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9945 a_3369760_754598# a_3366260_744206# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9946 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9947 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9948 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9949 w_3263498_541854# a_3400801_701658# a_3400801_701658# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9950 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9951 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9952 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9953 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9954 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9955 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9956 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9957 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9958 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9959 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9960 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9961 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9962 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9963 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9964 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9965 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9966 a_3359810_749958# a_3362834_747994# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9967 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9968 w_3185490_798160# a_3407542_688639# a_3405154_692359# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9969 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9970 w_3263498_541854# a_3400801_701658# a_3381563_717833# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9971 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9972 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9973 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9974 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9975 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9976 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9977 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9978 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9979 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9980 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X9981 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9982 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9983 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9984 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9985 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9986 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9987 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9988 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9989 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9990 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9991 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9992 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9993 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9994 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9995 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9996 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9997 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9998 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9999 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10000 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10001 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10002 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10003 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10004 a_3403286_717614# a_3403189_717414# w_3403067_716474# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10005 w_3422393_701565# a_3422243_697443# a_3420293_701761# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10006 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10007 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10008 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10009 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10010 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10011 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10012 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10013 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10014 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10015 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10016 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10017 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10018 a_3420382_721009# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10019 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10020 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10021 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10022 w_3263498_541854# a_3408579_674425# a_3408579_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10023 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
R9 w_3263498_541854# w_3474538_503344# sky130_fd_pr__res_generic_m5 w=7.4e+07u l=1.005e+07u
X10024 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10025 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10026 a_3400801_715182# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10027 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10028 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10029 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10030 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10031 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10032 a_3335479_772599# a_3359810_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10033 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10034 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10035 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10036 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X10037 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10038 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10039 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10040 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10041 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10042 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10043 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10044 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10045 a_3428294_754598# a_3434368_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10046 a_3366260_744206# a_3369760_747574# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10047 w_3422393_701565# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10048 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10049 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10050 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10051 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10052 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10053 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10054 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10055 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10056 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10057 w_3185490_798160# a_3399027_674337# a_3405057_686207# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X10058 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10059 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10060 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10061 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10062 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10063 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10064 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10065 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10066 a_3407542_687895# a_3407282_686697# w_3407323_687499# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10067 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10068 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10069 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10070 a_3379175_700273# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10071 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10072 a_3394410_687695# a_3387775_698875# w_3396510_687499# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10073 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10074 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10075 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10076 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10077 w_3263498_541854# a_3401256_686207# a_3401256_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10078 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10079 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10080 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10081 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10082 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10083 w_3185490_798160# a_3407542_687895# a_3407542_688639# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10084 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10085 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10086 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10087 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10088 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10089 a_3436064_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X10090 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10091 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10092 w_3185490_798160# a_3381660_718033# a_3381660_718033# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10093 a_3405057_686207# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10094 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10095 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10096 w_3396510_687499# a_3387775_698875# a_3394410_687695# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10097 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10098 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10099 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10100 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10101 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10102 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10103 w_3403067_702950# a_3381563_702505# a_3403286_704090# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10104 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10105 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10106 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10107 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10108 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10109 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10110 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10111 w_3185490_798160# a_3366260_744206# a_3369760_754598# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10112 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10113 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10114 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10115 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10116 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10117 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10118 a_3436064_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X10119 a_3403286_716870# a_3381563_702505# w_3403067_716474# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10120 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10121 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10122 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10123 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10124 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10125 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10126 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10127 w_3185490_798160# a_3403286_716870# a_3403286_717614# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10128 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10129 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10130 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10131 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10132 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10133 w_3422394_717637# a_3381563_717833# a_3420294_717833# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10134 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10135 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10136 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10137 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10138 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10139 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10140 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10141 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10142 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10143 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10144 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10145 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10146 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10147 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10148 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10149 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10150 a_3443016_749796# a_3439418_744112# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10151 v2 a_3434368_749958# a_3428294_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10152 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10153 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10154 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10155 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10156 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10157 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10158 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10159 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10160 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10161 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10162 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10163 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10164 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10165 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10166 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10167 w_3263498_541854# a_3407435_674425# a_3407435_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10168 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10169 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10170 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10171 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10172 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10173 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10174 a_3381563_717833# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10175 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10176 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10177 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10178 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10179 w_3263498_541854# a_3379175_700273# a_3379175_700273# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10180 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10181 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10182 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10183 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10184 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10185 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10186 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10187 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10188 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10189 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10190 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10191 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10192 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10193 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10194 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10195 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10196 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10197 w_3381441_701565# a_3381563_702505# a_3381660_702705# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10198 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10199 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10200 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10201 a_3436064_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X10202 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10203 a_3335479_772599# a_3359810_749958# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10204 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10205 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10206 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10207 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10208 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10209 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10210 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10211 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10212 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10213 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10214 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10215 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10216 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10217 a_3408579_674425# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10218 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10219 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10220 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10221 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10222 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10223 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10224 a_3436064_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X10225 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10226 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10227 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10228 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10229 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10230 w_3263498_541854# a_3408579_674425# w_3422394_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10231 a_3446663_700871# a_3427310_772647# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X10232 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10233 a_3369760_754598# a_3366260_744206# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10234 a_3335479_772599# a_3359810_749958# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10235 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X10236 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10237 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10238 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10239 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10240 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10241 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10242 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10243 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10244 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10245 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10246 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10247 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10248 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10249 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10250 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10251 a_3407435_674425# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10252 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10253 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10254 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10255 a_3403286_717614# a_3403286_716870# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10256 w_3407323_687499# a_3407282_686697# a_3407542_687895# w_3407323_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10257 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10258 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10259 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10260 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10261 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10262 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10263 a_3403286_704090# a_3403286_703346# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10264 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10265 w_3396510_687499# a_3387775_698875# a_3394410_687695# w_3396510_687499# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10266 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10267 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10268 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10269 a_3369760_754598# a_3366260_744206# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10270 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10271 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10272 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10273 a_3359663_699917# a_3361095_700235# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X10274 w_3263498_541854# a_3401256_686207# w_3396510_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10275 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10276 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10277 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10278 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10279 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10280 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10281 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10282 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10283 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10284 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10285 a_3403286_716870# a_3381563_702505# w_3403067_716474# w_3403067_716474# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10286 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10287 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10288 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10289 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10290 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10291 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10292 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10293 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10294 w_3263498_541854# a_3408579_674425# a_3408579_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10295 w_3185490_798160# a_3407542_687895# a_3407542_688639# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10296 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10297 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10298 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10299 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10300 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10301 a_3420382_721009# a_3420294_720809# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10302 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10303 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10304 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10305 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10306 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10307 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10308 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10309 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10310 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10311 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10312 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10313 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10314 w_3403067_716474# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10315 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10316 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10317 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10318 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10319 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10320 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10321 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10322 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10323 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10324 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10325 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10326 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X10327 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10328 a_3400898_721334# a_3403286_717614# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10329 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10330 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X10331 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10332 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10333 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10334 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10335 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10336 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10337 w_3185490_798160# a_3403286_716870# a_3403286_716870# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10338 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10339 a_3379175_700273# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10340 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10341 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10342 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10343 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10344 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10345 a_3381660_718033# a_3381660_718033# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10346 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10347 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10348 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10349 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10350 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10351 w_3263498_541854# a_3401256_686207# a_3401256_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10352 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10353 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10354 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10355 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10356 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10357 a_3387457_697443# a_3387139_698875# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X10358 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10359 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10360 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10361 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10362 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10363 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10364 w_3185490_798160# a_3403286_716870# a_3403286_717614# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10365 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10366 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10367 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10368 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10369 a_3379175_716345# a_3399027_674337# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X10370 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10371 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X10372 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10373 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10374 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10375 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10376 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10377 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10378 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10379 a_3436064_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X10380 v2 a_3439418_744112# a_3443016_749796# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10381 a_3379272_706425# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10382 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10383 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10384 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10385 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10386 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10387 w_3407323_687499# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10388 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10389 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10390 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10391 a_3400801_701658# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10392 w_3185490_798160# a_3403286_703346# a_3403286_703346# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10393 a_3366422_743586# a_3381660_718777# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10394 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10395 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10396 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10397 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10398 w_3263498_541854# a_3405057_686207# a_3405057_686207# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10399 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10400 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10401 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10402 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10403 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10404 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X10405 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10406 a_3436064_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X10407 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10408 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10409 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10410 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10411 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10412 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10413 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10414 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10415 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10416 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10417 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10418 w_3185490_798160# a_3420293_704737# a_3420381_704937# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10419 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10420 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10421 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10422 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10423 w_3185490_798160# a_3381660_702705# a_3379272_706425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10424 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10425 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10426 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10427 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10428 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10429 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10430 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10431 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10432 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10433 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10434 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10435 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10436 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10437 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10438 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10439 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10440 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10441 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10442 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10443 w_3263498_541854# a_3400801_701658# a_3400801_701658# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10444 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10445 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10446 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10447 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10448 w_3263498_541854# a_3400801_715182# a_3400898_721334# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10449 w_3185490_798160# a_3403286_717614# a_3400898_721334# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10450 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10451 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10452 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10453 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10454 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10455 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10456 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10457 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10458 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10459 a_3403286_717614# a_3403286_716870# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10460 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10461 a_3405154_692359# a_3405057_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10462 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10463 a_3403286_703346# a_3403286_703346# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10464 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10465 a_3407282_686697# a_3409354_691535# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X10466 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10467 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10468 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10469 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10470 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10471 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10472 w_3381441_701565# a_3361095_699281# a_3381660_701961# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10473 a_3362906_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X10474 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10475 w_3263498_541854# w_3685938_653428# sky130_fd_pr__diode_pd2nw_05v5 area=2.25e+16p
X10476 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10477 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10478 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10479 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10480 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10481 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10482 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10483 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10484 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10485 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10486 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10487 w_3185490_798160# a_3394410_690671# a_3387775_698875# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10488 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10489 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10490 a_3362906_746854# a_3366260_744206# a_3366286_744142# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10491 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10492 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10493 w_3422393_701565# a_3381563_702505# a_3420293_704737# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10494 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10495 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X10496 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10497 a_3381660_701961# a_3381660_701961# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10498 w_3263498_541854# a_3408579_674425# w_3422394_717637# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10499 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10500 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10501 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10502 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10503 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10504 a_3361629_772599# a_3369760_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10505 w_3185490_798160# a_3407542_687895# a_3407542_687895# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10506 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10507 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10508 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10509 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10510 a_3400898_721334# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10511 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10512 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10513 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10514 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10515 a_3400801_715182# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10516 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10517 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10518 a_3420971_697443# a_3421289_698875# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X10519 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10520 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10521 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10522 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10523 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10524 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10525 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10526 a_3400801_715182# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10527 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10528 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10529 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10530 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10531 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10532 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10533 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10534 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10535 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10536 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10537 a_3422243_697443# a_3420381_704937# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X10538 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10539 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10540 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10541 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10542 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10543 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10544 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10545 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10546 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10547 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10548 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10549 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10550 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10551 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10552 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10553 a_3379175_700273# a_3379175_700273# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10554 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10555 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10556 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10557 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10558 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10559 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10560 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10561 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10562 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10563 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10564 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10565 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10566 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10567 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10568 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10569 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10570 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10571 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10572 a_3403001_700774# a_3381563_717833# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X10573 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10574 w_3263498_541854# a_3407435_674425# a_3420381_704937# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10575 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10576 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10577 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10578 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10579 a_3446663_699599# a_3448095_699281# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X10580 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10581 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10582 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10583 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10584 a_3381660_701961# a_3361095_699281# w_3381441_701565# w_3381441_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10585 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10586 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10587 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10588 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10589 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10590 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10591 w_3263498_541854# a_3407435_674425# w_3422393_701565# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10592 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10593 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10594 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10595 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10596 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10597 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10598 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10599 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10600 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10601 w_3403067_702950# a_3403001_700774# a_3403286_703346# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10602 w_3403067_702950# a_3400801_701658# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10603 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10604 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10605 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10606 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10607 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10608 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10609 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10610 a_3428294_754598# a_3434368_749958# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10611 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10612 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10613 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10614 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10615 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10616 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10617 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10618 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10619 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10620 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10621 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10622 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10623 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10624 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10625 a_3387775_698875# a_3394410_690671# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10626 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10627 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10628 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10629 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10630 a_3427213_772599# a_3428294_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10631 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10632 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10633 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10634 a_3387775_698875# a_3401256_686207# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10635 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10636 a_3428294_754598# a_3434368_749958# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10637 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10638 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10639 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10640 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10641 w_3263498_541854# a_3379175_716345# a_3366422_743586# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10642 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10643 a_3420294_717833# a_3381563_717833# w_3422394_717637# w_3422394_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10644 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10645 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10646 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10647 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10648 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10649 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10650 w_3185490_798160# a_3403286_716870# a_3403286_716870# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10651 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10652 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10653 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10654 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10655 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10656 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10657 a_3420381_704937# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10658 w_3185490_798160# a_3369760_754598# a_3361629_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10659 w_3263498_541854# a_3400801_701658# w_3403067_702950# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10660 w_3263498_541854# a_3407435_674425# a_3407435_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10661 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10662 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10663 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10664 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10665 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10666 a_3362906_746854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X10667 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10668 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10669 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10670 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10671 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10672 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10673 a_3403286_704090# a_3381563_702505# w_3403067_702950# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10674 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10675 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10676 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10677 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10678 a_3434368_749958# a_3435992_747994# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10679 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10680 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10681 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10682 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10683 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10684 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10685 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10686 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10687 w_3185490_798160# a_3420294_720809# a_3420382_721009# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10688 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10689 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10690 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10691 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10692 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10693 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10694 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10695 a_3362906_746854# a_3366260_744112# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10696 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10697 a_3361629_772599# a_3369760_754598# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10698 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10699 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10700 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10701 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10702 a_3381660_718033# a_3381563_717833# w_3381441_717637# w_3381441_717637# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10703 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10704 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10705 w_3381441_717637# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10706 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10707 w_3422393_701565# a_3422243_697443# a_3420293_701761# w_3422393_701565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10708 v2 a_3366260_744206# a_3369760_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10709 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10710 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10711 a_3408579_674425# a_3408579_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10712 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10713 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10714 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10715 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10716 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10717 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10718 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10719 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10720 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10721 a_3403286_717614# a_3403286_716870# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10722 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10723 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X10724 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10725 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10726 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10727 v2 a_3362834_747994# a_3359810_749958# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10728 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10729 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10730 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10731 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10732 w_3263498_541854# a_3400801_701658# w_3403067_702950# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10733 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10734 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10735 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10736 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10737 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10738 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10739 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10740 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10741 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10742 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10743 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10744 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10745 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10746 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10747 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10748 a_3407435_674425# a_3407435_674425# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10749 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10750 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10751 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10752 v2 a_3369760_754598# a_3361629_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10753 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10754 w_3263498_541854# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10755 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10756 v2 a_3428294_754598# a_3427213_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10757 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10758 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10759 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10760 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10761 a_3403286_716870# a_3403286_716870# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10762 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10763 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10764 w_3185490_798160# v2 sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X10765 w_3403067_702950# a_3381563_702505# a_3403286_704090# w_3403067_702950# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10766 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10767 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10768 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10769 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10770 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10771 a_3443016_749796# a_3439418_744112# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10772 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10773 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10774 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10775 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10776 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10777 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10778 w_3263498_541854# a_3379175_700273# a_3379272_706425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10779 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10780 a_3366422_743586# a_3379175_716345# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10781 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10782 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10783 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10784 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10785 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10786 a_3422243_697443# a_3421925_698875# w_3185490_798160# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X10787 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10788 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10789 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10790 w_3263498_541854# a_3401256_686207# w_3396510_687499# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10791 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10792 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10793 a_3405154_692359# a_3407542_688639# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10794 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10795 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10796 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10797 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10798 a_3285528_930602# a_3335479_772599# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10799 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10800 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10801 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10802 a_3427213_772599# a_3428294_754598# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10803 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10804 a_3403286_703346# a_3403286_703346# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10805 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10806 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10807 w_3263498_541854# a_3408579_674425# a_3408579_674425# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10808 v2 a_3359810_749958# a_3335479_772599# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10809 a_3379272_706425# a_3381660_702705# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10810 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10811 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10812 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10813 w_3185490_798160# a_3407542_687895# a_3407542_688639# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10814 a_3399027_674337# w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10815 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10816 w_3185490_798160# a_3443016_749796# a_3427310_772647# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10817 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10818 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10819 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10820 v2 a_3434368_749958# a_3428294_754598# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10821 v2 a_3369760_747574# a_3366260_744206# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10822 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10823 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10824 w_3185490_798160# a_3335479_772599# a_3285528_930602# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10825 w_3403067_716474# a_3400801_715182# w_3263498_541854# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10826 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10827 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10828 a_3427310_772647# a_3443016_749796# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10829 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10830 w_3185490_798160# a_3399027_674337# a_3407435_674425# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X10831 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10832 a_3367712_744142# w_3185490_798160# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X10833 a_3420381_704937# a_3420293_704737# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10834 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10835 a_3285528_930602# a_3361629_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10836 v2 w_3185490_798160# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10837 w_3263498_541854# a_3405057_686207# a_3405154_692359# w_3263498_541854# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10838 v2 a_3361629_772599# a_3285528_930602# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10839 a_3420293_701761# a_3420293_701761# w_3185490_798160# w_3185490_798160# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10840 w_3185490_798160# a_3428294_754598# a_3427213_772599# w_3185490_798160# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10841 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10842 a_3427310_772647# a_3427213_772599# v2 v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10843 v2 a_3427213_772599# a_3427310_772647# v2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
.end

