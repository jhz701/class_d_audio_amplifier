* NGSPICE file created from triangle_revised_flat.ext - technology: sky130A


* Top level circuit triangle_revised_flat

X0 vdd vbias2 vbias2 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u M=24
X1 w_1705_3239# vbias1 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u M=24
X2 a_1901_1139# a_1901_1139# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u M=16
X3 vdd vbias2 vsquare vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u M=48
X4 vss a_15425_1139# a_15425_1139# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u M=16
X5 vss a_16369_1227# vsquare vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u M=64
X6 vdd vbias1 vt vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u M=48
X7 vss a_2845_1227# vt vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u M=64
X8 a_16369_1227# vref w_15229_3239# w_15229_3239# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u M=16
X9 a_n1703_5991# a_n471_5673# vss sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X10 vdd vbias2 w_15229_3239# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u M=24
X11 a_1901_1139# vref w_1705_3239# w_1705_3239# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u M=16
X12 a_15425_1139# vref w_15229_3239# w_15229_3239# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u M=16
X13 a_2845_1227# a_1901_1139# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u M=16
X14 a_16369_1227# a_20559_4831# vss sky130_fd_pr__res_xhigh_po w=350000u l=500000u
X15 w_1705_3239# vref a_2845_1227# w_1705_3239# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u M=16
X16 vref vt sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X17 a_n1703_6627# a_n471_6309# vss sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X18 vref vt sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X19 vdd vbias1 vbias1 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u M=24
X20 vref vt sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X21 a_2845_1227# a_5497_5073# vss sky130_fd_pr__res_xhigh_po w=350000u l=2.8e+06u
X22 vref vt sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X23 a_n1703_5355# a_n471_5673# vss sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X24 a_16369_1227# a_15425_1139# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u M=16
X25 vref vt sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X26 a_n1703_5991# a_n471_6309# vss sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X27 vt vref vss sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X28 a_n1703_5355# vsquare vss sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X29 a_n1703_7263# vref vss sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X30 vref vsquare vss sky130_fd_pr__res_xhigh_po w=350000u l=9e+06u
X31 vref vt sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X32 vref vt sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X33 a_n1703_7263# a_n471_6945# vss sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X34 a_20559_4831# vsquare sky130_fd_pr__cap_mim_m3_1 l=1.4e+07u w=1.4e+07u
X35 a_5497_5073# vt sky130_fd_pr__cap_mim_m3_1 l=1.8e+07u w=2.7e+07u
X36 a_n1703_6627# a_n471_6945# vss sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X37 vref vt sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
.end

