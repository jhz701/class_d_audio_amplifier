* NGSPICE file created from half_driver_revised.ext - technology: sky130A

.subckt half_driver_post vdd vss vp_p out_p vp_n
X0 vdd.t2999 vp_p.t0 out_p.t2284 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1 vdd.t2998 vp_p.t1 out_p.t2283 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2 out_p.t2282 vp_p.t2 vdd.t2997 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3 out_p.t422 vp_n.t0 vss.t599 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4 vdd.t2996 vp_p.t3 out_p.t2281 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5 out_p.t2280 vp_p.t4 vdd.t2995 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6 vdd.t2994 vp_p.t5 out_p.t2262 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7 out_p.t2261 vp_p.t6 vdd.t2993 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8 out_p.t2260 vp_p.t7 vdd.t2992 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9 out_p.t2259 vp_p.t8 vdd.t2991 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10 out_p.t2258 vp_p.t9 vdd.t2990 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X11 out_p.t3468 vp_n.t1 vss.t598 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X12 out_p.t2257 vp_p.t10 vdd.t2989 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X13 out_p.t2248 vp_p.t11 vdd.t2988 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X14 vdd.t2987 vp_p.t12 out_p.t2247 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X15 vdd.t2986 vp_p.t13 out_p.t2246 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X16 out_p.t2245 vp_p.t14 vdd.t2985 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X17 out_p.t2244 vp_p.t15 vdd.t2984 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X18 vdd.t2983 vp_p.t16 out_p.t2243 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X19 out_p.t2225 vp_p.t17 vdd.t2982 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X20 vdd.t2981 vp_p.t18 out_p.t2224 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X21 vdd.t2980 vp_p.t19 out_p.t2223 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X22 out_p.t2222 vp_p.t20 vdd.t2979 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X23 out_p.t2221 vp_p.t21 vdd.t2978 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X24 vdd.t2977 vp_p.t22 out_p.t2220 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X25 out_p.t2212 vp_p.t23 vdd.t2976 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X26 out_p.t2211 vp_p.t24 vdd.t2975 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X27 out_p.t2210 vp_p.t25 vdd.t2974 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X28 out_p.t2209 vp_p.t26 vdd.t2973 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X29 vdd.t2972 vp_p.t27 out_p.t2208 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X30 out_p.t2207 vp_p.t28 vdd.t2971 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X31 vdd.t2970 vp_p.t29 out_p.t2199 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X32 vdd.t2969 vp_p.t30 out_p.t2198 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X33 out_p.t2197 vp_p.t31 vdd.t2968 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X34 out_p.t2196 vp_p.t32 vdd.t2967 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X35 out_p.t2195 vp_p.t33 vdd.t2966 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X36 vdd.t2965 vp_p.t34 out_p.t2194 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X37 vdd.t2964 vp_p.t35 out_p.t2176 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X38 out_p.t2175 vp_p.t36 vdd.t2963 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X39 out_p.t2174 vp_p.t37 vdd.t2962 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X40 vdd.t2961 vp_p.t38 out_p.t2173 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X41 out_p.t2172 vp_p.t39 vdd.t2960 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X42 vdd.t2959 vp_p.t40 out_p.t2171 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X43 vdd.t2958 vp_p.t41 out_p.t2163 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X44 vdd.t2957 vp_p.t42 out_p.t2162 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X45 vdd.t2956 vp_p.t43 out_p.t2161 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X46 out_p.t2160 vp_p.t44 vdd.t2955 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X47 vdd.t2954 vp_p.t45 out_p.t2159 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X48 out_p.t2158 vp_p.t46 vdd.t2953 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X49 out_p.t2140 vp_p.t47 vdd.t2952 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X50 out_p.t2139 vp_p.t48 vdd.t2951 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X51 out_p.t2138 vp_p.t49 vdd.t2950 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X52 vdd.t2949 vp_p.t50 out_p.t2137 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X53 out_p.t2136 vp_p.t51 vdd.t2948 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X54 out_p.t3467 vp_n.t2 vss.t597 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X55 vss.t596 vp_n.t3 out_p.t3460 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X56 vdd.t2947 vp_p.t52 out_p.t2135 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X57 out_p.t2117 vp_p.t53 vdd.t2946 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X58 vdd.t2945 vp_p.t54 out_p.t2116 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X59 out_p.t2115 vp_p.t55 vdd.t2944 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X60 vdd.t2943 vp_p.t56 out_p.t2114 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X61 out_p.t2113 vp_p.t57 vdd.t2942 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X62 out_p.t2112 vp_p.t58 vdd.t2941 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X63 vss.t595 vp_n.t4 out_p.t3456 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X64 out_p.t2093 vp_p.t59 vdd.t2940 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X65 out_p.t2092 vp_p.t60 vdd.t2939 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X66 out_p.t2091 vp_p.t61 vdd.t2938 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X67 out_p.t2090 vp_p.t62 vdd.t2937 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X68 vdd.t2936 vp_p.t63 out_p.t2089 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X69 out_p.t2088 vp_p.t64 vdd.t2935 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X70 out_p.t2070 vp_p.t65 vdd.t2934 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X71 out_p.t2069 vp_p.t66 vdd.t2933 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X72 vdd.t2932 vp_p.t67 out_p.t2068 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X73 vdd.t2931 vp_p.t68 out_p.t2067 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X74 out_p.t2066 vp_p.t69 vdd.t2930 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X75 out_p.t2065 vp_p.t70 vdd.t2929 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X76 vdd.t2928 vp_p.t71 out_p.t2047 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X77 out_p.t2046 vp_p.t72 vdd.t2927 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X78 out_p.t2045 vp_p.t73 vdd.t2926 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X79 vdd.t2925 vp_p.t74 out_p.t2044 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X80 out_p.t2043 vp_p.t75 vdd.t2924 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X81 vss.t594 vp_n.t5 out_p.t3472 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X82 vdd.t2923 vp_p.t76 out_p.t2042 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X83 out_p.t2024 vp_p.t77 vdd.t2922 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X84 vdd.t2921 vp_p.t78 out_p.t2023 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X85 vdd.t2920 vp_p.t79 out_p.t2022 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X86 vdd.t2919 vp_p.t80 out_p.t2021 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X87 vdd.t2918 vp_p.t81 out_p.t2020 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X88 vdd.t2917 vp_p.t82 out_p.t2019 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X89 vdd.t2916 vp_p.t83 out_p.t2001 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X90 vdd.t2915 vp_p.t84 out_p.t2000 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X91 out_p.t1999 vp_p.t85 vdd.t2914 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X92 out_p.t1998 vp_p.t86 vdd.t2913 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X93 out_p.t1997 vp_p.t87 vdd.t2912 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X94 vdd.t2911 vp_p.t88 out_p.t1996 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X95 vdd.t2910 vp_p.t89 out_p.t1978 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X96 out_p.t227 vp_n.t6 vss.t593 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X97 vdd.t2909 vp_p.t90 out_p.t1977 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X98 out_p.t1976 vp_p.t91 vdd.t2908 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X99 vdd.t2907 vp_p.t92 out_p.t1975 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X100 vdd.t2906 vp_p.t93 out_p.t1974 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X101 vdd.t2905 vp_p.t94 out_p.t1973 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X102 vdd.t2904 vp_p.t95 out_p.t1955 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X103 out_p.t1954 vp_p.t96 vdd.t2903 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X104 vdd.t2902 vp_p.t97 out_p.t1953 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X105 vss.t592 vp_n.t7 out_p.t236 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X106 vdd.t2901 vp_p.t98 out_p.t1952 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X107 vss.t591 vp_n.t8 out_p.t232 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X108 vdd.t2900 vp_p.t99 out_p.t1951 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X109 out_p.t1950 vp_p.t100 vdd.t2899 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X110 out_p.t1942 vp_p.t101 vdd.t2898 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X111 out_p.t1941 vp_p.t102 vdd.t2897 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X112 out_p.t230 vp_n.t9 vss.t590 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X113 out_p.t1940 vp_p.t103 vdd.t2896 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X114 vdd.t2895 vp_p.t104 out_p.t1939 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X115 vdd.t2894 vp_p.t105 out_p.t1938 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X116 vdd.t2893 vp_p.t106 out_p.t1937 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X117 out_p.t1919 vp_p.t107 vdd.t2892 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X118 out_p.t1918 vp_p.t108 vdd.t2891 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X119 vdd.t2890 vp_p.t109 out_p.t1917 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X120 out_p.t229 vp_n.t10 vss.t589 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X121 vdd.t2889 vp_p.t110 out_p.t1916 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X122 vdd.t2888 vp_p.t111 out_p.t1915 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X123 out_p.t1914 vp_p.t112 vdd.t2887 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X124 out_p.t1896 vp_p.t113 vdd.t2886 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X125 out_p.t1895 vp_p.t114 vdd.t2885 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X126 out_p.t1894 vp_p.t115 vdd.t2884 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X127 vdd.t2883 vp_p.t116 out_p.t1893 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X128 out_p.t1892 vp_p.t117 vdd.t2882 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X129 vdd.t2881 vp_p.t118 out_p.t1891 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X130 vdd.t2880 vp_p.t119 out_p.t1873 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X131 out_p.t1872 vp_p.t120 vdd.t2879 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X132 out_p.t1871 vp_p.t121 vdd.t2878 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X133 vdd.t2877 vp_p.t122 out_p.t1870 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X134 out_p.t1869 vp_p.t123 vdd.t2876 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X135 vss.t588 vp_n.t11 out_p.t231 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X136 out_p.t1868 vp_p.t124 vdd.t2875 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X137 vss.t587 vp_n.t12 out_p.t228 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X138 out_p.t226 vp_n.t13 vss.t586 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X139 vdd.t2874 vp_p.t125 out_p.t1850 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X140 vdd.t2873 vp_p.t126 out_p.t1849 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X141 vdd.t2872 vp_p.t127 out_p.t1848 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X142 vdd.t2871 vp_p.t128 out_p.t1847 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X143 vdd.t2870 vp_p.t129 out_p.t1846 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X144 out_p.t1845 vp_p.t130 vdd.t2869 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X145 vdd.t2868 vp_p.t131 out_p.t1837 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X146 out_p.t1836 vp_p.t132 vdd.t2867 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X147 out_p.t1835 vp_p.t133 vdd.t2866 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X148 vdd.t2865 vp_p.t134 out_p.t1834 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X149 vdd.t2864 vp_p.t135 out_p.t1833 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X150 out_p.t1832 vp_p.t136 vdd.t2863 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X151 out_p.t1814 vp_p.t137 vdd.t2862 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X152 vdd.t2861 vp_p.t138 out_p.t1813 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X153 vdd.t2860 vp_p.t139 out_p.t1812 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X154 out_p.t1811 vp_p.t140 vdd.t2859 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X155 out_p.t1810 vp_p.t141 vdd.t2858 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X156 out_p.t233 vp_n.t14 vss.t585 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X157 out_p.t243 vp_n.t15 vss.t584 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X158 out_p.t1809 vp_p.t142 vdd.t2857 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X159 vdd.t2856 vp_p.t143 out_p.t1791 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X160 out_p.t1790 vp_p.t144 vdd.t2855 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X161 out_p.t1789 vp_p.t145 vdd.t2854 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X162 vdd.t2853 vp_p.t146 out_p.t1788 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X163 vdd.t2852 vp_p.t147 out_p.t1787 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X164 out_p.t1786 vp_p.t148 vdd.t2851 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X165 vdd.t2850 vp_p.t149 out_p.t1767 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X166 out_p.t1766 vp_p.t150 vdd.t2849 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X167 vdd.t2848 vp_p.t151 out_p.t1765 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X168 vdd.t2847 vp_p.t152 out_p.t1764 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X169 vdd.t2846 vp_p.t153 out_p.t1763 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X170 vss.t583 vp_n.t16 out_p.t242 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X171 vdd.t2845 vp_p.t154 out_p.t1762 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X172 vdd.t2844 vp_p.t155 out_p.t1744 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X173 vdd.t2843 vp_p.t156 out_p.t1743 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X174 vdd.t2842 vp_p.t157 out_p.t1742 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X175 vdd.t2841 vp_p.t158 out_p.t1741 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X176 vdd.t2840 vp_p.t159 out_p.t1740 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X177 vdd.t2839 vp_p.t160 out_p.t1739 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X178 out_p.t1731 vp_p.t161 vdd.t2838 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X179 vdd.t2837 vp_p.t162 out_p.t1730 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X180 out_p.t1729 vp_p.t163 vdd.t2836 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X181 out_p.t1728 vp_p.t164 vdd.t2835 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X182 out_p.t1727 vp_p.t165 vdd.t2834 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X183 vss.t582 vp_n.t17 out_p.t240 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X184 out_p.t239 vp_n.t18 vss.t581 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X185 vdd.t2833 vp_p.t166 out_p.t1726 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X186 vdd.t2832 vp_p.t167 out_p.t1708 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X187 vdd.t2831 vp_p.t168 out_p.t1707 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X188 vdd.t2830 vp_p.t169 out_p.t1706 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X189 vdd.t2829 vp_p.t170 out_p.t1705 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X190 out_p.t1704 vp_p.t171 vdd.t2828 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X191 out_p.t1703 vp_p.t172 vdd.t2827 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X192 out_p.t238 vp_n.t19 vss.t580 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X193 out_p.t1685 vp_p.t173 vdd.t2826 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X194 vdd.t2825 vp_p.t174 out_p.t1684 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X195 vdd.t2824 vp_p.t175 out_p.t1683 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X196 vdd.t2823 vp_p.t176 out_p.t1682 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X197 vss.t579 vp_n.t20 out_p.t237 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X198 out_p.t1681 vp_p.t177 vdd.t2822 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X199 vdd.t2821 vp_p.t178 out_p.t1680 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X200 vss.t578 vp_n.t21 out_p.t235 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X201 vdd.t2820 vp_p.t179 out_p.t1662 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X202 out_p.t1661 vp_p.t180 vdd.t2819 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X203 out_p.t244 vp_n.t22 vss.t577 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X204 vdd.t2818 vp_p.t181 out_p.t1660 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X205 out_p.t1659 vp_p.t182 vdd.t2817 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X206 vdd.t2816 vp_p.t183 out_p.t1658 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X207 out_p.t1657 vp_p.t184 vdd.t2815 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X208 out_p.t1638 vp_p.t185 vdd.t2814 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X209 out_p.t1637 vp_p.t186 vdd.t2813 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X210 out_p.t256 vp_n.t23 vss.t576 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X211 vdd.t2812 vp_p.t187 out_p.t1636 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X212 vdd.t2811 vp_p.t188 out_p.t1635 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X213 out_p.t255 vp_n.t24 vss.t575 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X214 vss.t574 vp_n.t25 out_p.t3444 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X215 out_p.t1634 vp_p.t189 vdd.t2810 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X216 out_p.t1633 vp_p.t190 vdd.t2809 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X217 out_p.t1596 vp_p.t191 vdd.t2808 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X218 out_p.t1595 vp_p.t192 vdd.t2807 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X219 out_p.t1594 vp_p.t193 vdd.t2806 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X220 vdd.t2805 vp_p.t194 out_p.t1593 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X221 out_p.t253 vp_n.t26 vss.t573 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X222 out_p.t1592 vp_p.t195 vdd.t2804 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X223 out_p.t1591 vp_p.t196 vdd.t2803 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X224 vdd.t2802 vp_p.t197 out_p.t1573 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X225 vdd.t2801 vp_p.t198 out_p.t1572 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X226 vdd.t2800 vp_p.t199 out_p.t1571 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X227 vss.t572 vp_n.t27 out_p.t251 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X228 out_p.t1570 vp_p.t200 vdd.t2799 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X229 vss.t571 vp_n.t28 out_p.t249 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X230 out_p.t1569 vp_p.t201 vdd.t2798 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X231 vdd.t2797 vp_p.t202 out_p.t1568 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X232 out_p.t1550 vp_p.t203 vdd.t2796 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X233 vdd.t2795 vp_p.t204 out_p.t1549 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X234 out_p.t247 vp_n.t29 vss.t570 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X235 out_p.t1548 vp_p.t205 vdd.t2794 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X236 vdd.t2793 vp_p.t206 out_p.t1547 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X237 out_p.t1546 vp_p.t207 vdd.t2792 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X238 out_p.t260 vp_n.t30 vss.t569 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X239 out_p.t1545 vp_p.t208 vdd.t2791 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X240 vss.t568 vp_n.t31 out_p.t268 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X241 out_p.t1527 vp_p.t209 vdd.t2790 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X242 out_p.t1526 vp_p.t210 vdd.t2789 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X243 vdd.t2788 vp_p.t211 out_p.t1525 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X244 vdd.t2787 vp_p.t212 out_p.t1524 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X245 out_p.t265 vp_n.t32 vss.t567 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X246 out_p.t1523 vp_p.t213 vdd.t2786 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X247 vdd.t2785 vp_p.t214 out_p.t1522 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X248 vdd.t2784 vp_p.t215 out_p.t1514 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X249 out_p.t1513 vp_p.t216 vdd.t2783 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X250 vdd.t2782 vp_p.t217 out_p.t1512 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X251 vss.t566 vp_n.t33 out_p.t264 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X252 vdd.t2781 vp_p.t218 out_p.t1511 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X253 out_p.t1510 vp_p.t219 vdd.t2780 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X254 vss.t565 vp_n.t34 out_p.t263 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X255 vdd.t2779 vp_p.t220 out_p.t1509 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X256 out_p.t1473 vp_p.t221 vdd.t2778 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X257 out_p.t1472 vp_p.t222 vdd.t2777 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X258 out_p.t1471 vp_p.t223 vdd.t2776 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X259 out_p.t261 vp_n.t35 vss.t564 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X260 vdd.t2775 vp_p.t224 out_p.t1470 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X261 out_p.t1469 vp_p.t225 vdd.t2774 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X262 out_p.t345 vp_n.t36 vss.t563 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X263 vss.t562 vp_n.t37 out_p.t267 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X264 out_p.t1468 vp_p.t226 vdd.t2773 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X265 vdd.t2772 vp_p.t227 out_p.t1449 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X266 out_p.t250 vp_n.t38 vss.t561 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X267 out_p.t1448 vp_p.t228 vdd.t2771 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X268 vdd.t2770 vp_p.t229 out_p.t1447 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X269 out_p.t3500 vp_n.t39 vss.t560 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X270 out_p.t1446 vp_p.t230 vdd.t2769 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X271 vss.t559 vp_n.t40 out_p.t330 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X272 vdd.t2768 vp_p.t231 out_p.t1445 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X273 vss.t558 vp_n.t41 out_p.t157 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X274 out_p.t1444 vp_p.t232 vdd.t2767 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X275 vss.t557 vp_n.t42 out_p.t3578 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X276 out_p.t1407 vp_p.t233 vdd.t2766 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X277 out_p.t1406 vp_p.t234 vdd.t2765 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X278 vdd.t2764 vp_p.t235 out_p.t1405 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X279 vdd.t2763 vp_p.t236 out_p.t1404 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X280 vss.t556 vp_n.t43 out_p.t3572 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X281 vdd.t2762 vp_p.t237 out_p.t1403 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X282 vdd.t2761 vp_p.t238 out_p.t1402 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X283 out_p.t1365 vp_p.t239 vdd.t2760 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X284 out_p.t331 vp_n.t44 vss.t555 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X285 vdd.t2759 vp_p.t240 out_p.t1364 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X286 out_p.t1363 vp_p.t241 vdd.t2758 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X287 out_p.t1362 vp_p.t242 vdd.t2757 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X288 vss.t554 vp_n.t45 out_p.t332 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X289 vdd.t2756 vp_p.t243 out_p.t1361 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X290 vdd.t2755 vp_p.t244 out_p.t1360 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X291 out_p.t334 vp_n.t46 vss.t553 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X292 vdd.t2754 vp_p.t245 out_p.t2473 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X293 out_p.t2472 vp_p.t246 vdd.t2753 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X294 vss.t552 vp_n.t47 out_p.t320 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X295 out_p.t323 vp_n.t48 vss.t551 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X296 out_p.t325 vp_n.t49 vss.t550 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X297 vss.t549 vp_n.t50 out_p.t326 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X298 vdd.t2752 vp_p.t247 out_p.t2471 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X299 vss.t548 vp_n.t51 out_p.t337 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X300 out_p.t3523 vp_n.t52 vss.t547 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X301 out_p.t2470 vp_p.t248 vdd.t2751 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X302 vss.t546 vp_n.t53 out_p.t3515 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X303 out_p.t2469 vp_p.t249 vdd.t2750 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X304 vdd.t2749 vp_p.t250 out_p.t2468 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X305 vss.t545 vp_n.t54 out_p.t3505 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X306 vdd.t2748 vp_p.t251 out_p.t2462 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X307 vdd.t2747 vp_p.t252 out_p.t2461 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X308 vdd.t2746 vp_p.t253 out_p.t2460 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X309 out_p.t2459 vp_p.t254 vdd.t2745 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X310 vdd.t2744 vp_p.t255 out_p.t2458 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X311 out_p.t2457 vp_p.t256 vdd.t2743 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X312 vss.t544 vp_n.t55 out_p.t3499 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X313 out_p.t350 vp_n.t56 vss.t543 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X314 vdd.t2742 vp_p.t257 out_p.t2425 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X315 out_p.t2424 vp_p.t258 vdd.t2741 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X316 out_p.t2423 vp_p.t259 vdd.t2740 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X317 vdd.t2739 vp_p.t260 out_p.t2422 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X318 out_p.t2421 vp_p.t261 vdd.t2738 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X319 out_p.t2420 vp_p.t262 vdd.t2737 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X320 out_p.t351 vp_n.t57 vss.t542 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X321 vss.t541 vp_n.t58 out_p.t341 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X322 vss.t540 vp_n.t59 out_p.t342 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X323 vdd.t2736 vp_p.t263 out_p.t2414 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X324 vdd.t2735 vp_p.t264 out_p.t2413 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X325 out_p.t324 vp_n.t60 vss.t539 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X326 vdd.t2734 vp_p.t265 out_p.t2412 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X327 out_p.t2411 vp_p.t266 vdd.t2733 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X328 vss.t538 vp_n.t61 out_p.t3552 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X329 out_p.t2410 vp_p.t267 vdd.t2732 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X330 vdd.t2731 vp_p.t268 out_p.t2409 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X331 vss.t537 vp_n.t62 out_p.t3561 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X332 vdd.t2730 vp_p.t269 out_p.t2398 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X333 out_p.t2397 vp_p.t270 vdd.t2729 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X334 out_p.t2396 vp_p.t271 vdd.t2728 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X335 out_p.t2395 vp_p.t272 vdd.t2727 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X336 vss.t536 vp_n.t63 out_p.t258 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X337 out_p.t3564 vp_n.t64 vss.t535 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X338 vdd.t2726 vp_p.t273 out_p.t2394 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X339 vss.t534 vp_n.t65 out_p.t3524 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X340 vdd.t2725 vp_p.t274 out_p.t2393 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X341 vdd.t2724 vp_p.t275 out_p.t2387 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X342 out_p.t3506 vp_n.t66 vss.t533 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X343 vdd.t2723 vp_p.t276 out_p.t2386 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X344 out_p.t2385 vp_p.t277 vdd.t2722 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X345 out_p.t3508 vp_n.t67 vss.t532 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X346 vss.t531 vp_n.t68 out_p.t36 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X347 out_p.t2384 vp_p.t278 vdd.t2721 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X348 vdd.t2720 vp_p.t279 out_p.t2383 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X349 out_p.t2382 vp_p.t280 vdd.t2719 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X350 vdd.t2718 vp_p.t281 out_p.t2379 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X351 out_p.t158 vp_n.t69 vss.t530 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X352 out_p.t2378 vp_p.t282 vdd.t2717 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X353 out_p.t2377 vp_p.t283 vdd.t2716 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X354 out_p.t2376 vp_p.t284 vdd.t2715 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X355 vss.t529 vp_n.t70 out_p.t166 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X356 out_p.t171 vp_n.t71 vss.t528 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X357 out_p.t2375 vp_p.t285 vdd.t2714 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X358 vss.t527 vp_n.t72 out_p.t3567 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X359 out_p.t2374 vp_p.t286 vdd.t2713 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X360 vdd.t2712 vp_p.t287 out_p.t2368 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X361 vss.t526 vp_n.t73 out_p.t3529 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X362 out_p.t3537 vp_n.t74 vss.t525 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X363 out_p.t2367 vp_p.t288 vdd.t2711 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X364 vdd.t2710 vp_p.t289 out_p.t2366 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X365 out_p.t3542 vp_n.t75 vss.t524 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X366 out_p.t60 vp_n.t76 vss.t523 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X367 vss.t522 vp_n.t77 out_p.t57 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X368 out_p.t54 vp_n.t78 vss.t521 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X369 vdd.t2709 vp_p.t290 out_p.t2365 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X370 out_p.t2364 vp_p.t291 vdd.t2708 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X371 out_p.t2363 vp_p.t292 vdd.t2707 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X372 vdd.t2706 vp_p.t293 out_p.t2362 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X373 vdd.t2705 vp_p.t294 out_p.t2361 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X374 out_p.t51 vp_n.t79 vss.t520 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X375 vss.t519 vp_n.t80 out_p.t48 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X376 vdd.t2704 vp_p.t295 out_p.t2360 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X377 vdd.t2703 vp_p.t296 out_p.t2359 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X378 vss.t518 vp_n.t81 out_p.t45 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X379 out_p.t42 vp_n.t82 vss.t517 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X380 out_p.t2358 vp_p.t297 vdd.t2702 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X381 out_p.t2357 vp_p.t298 vdd.t2701 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X382 out_p.t2351 vp_p.t299 vdd.t2700 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X383 vdd.t2699 vp_p.t300 out_p.t2350 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X384 out_p.t2349 vp_p.t301 vdd.t2698 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X385 out_p.t2348 vp_p.t302 vdd.t2697 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X386 vdd.t2696 vp_p.t303 out_p.t2347 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X387 vss.t516 vp_n.t83 out_p.t39 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X388 out_p.t96 vp_n.t84 vss.t515 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X389 out_p.t2346 vp_p.t304 vdd.t2695 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X390 vdd.t2694 vp_p.t305 out_p.t2341 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X391 out_p.t2340 vp_p.t306 vdd.t2693 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X392 vdd.t2692 vp_p.t307 out_p.t2339 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X393 out_p.t2338 vp_p.t308 vdd.t2691 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X394 out_p.t2337 vp_p.t309 vdd.t2690 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X395 out_p.t93 vp_n.t85 vss.t514 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X396 out_p.t2336 vp_p.t310 vdd.t2689 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X397 out_p.t91 vp_n.t86 vss.t513 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X398 out_p.t2335 vp_p.t311 vdd.t2688 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X399 out_p.t2334 vp_p.t312 vdd.t2687 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X400 vdd.t2686 vp_p.t313 out_p.t2333 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X401 vdd.t2685 vp_p.t314 out_p.t2332 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X402 out_p.t2331 vp_p.t315 vdd.t2684 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X403 vdd.t2683 vp_p.t316 out_p.t2330 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X404 vdd.t2682 vp_p.t317 out_p.t2324 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X405 out_p.t88 vp_n.t87 vss.t512 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X406 out_p.t2323 vp_p.t318 vdd.t2681 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X407 out_p.t2322 vp_p.t319 vdd.t2680 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X408 out_p.t2321 vp_p.t320 vdd.t2679 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X409 vdd.t2678 vp_p.t321 out_p.t2320 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X410 vss.t511 vp_n.t88 out_p.t83 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X411 vdd.t2677 vp_p.t322 out_p.t2319 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X412 vdd.t2676 vp_p.t323 out_p.t2318 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X413 out_p.t71 vp_n.t89 vss.t510 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X414 vdd.t2675 vp_p.t324 out_p.t2317 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X415 out_p.t2316 vp_p.t325 vdd.t2674 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X416 vss.t509 vp_n.t90 out_p.t69 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X417 vdd.t2673 vp_p.t326 out_p.t2315 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X418 vdd.t2672 vp_p.t327 out_p.t2314 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X419 out_p.t2313 vp_p.t328 vdd.t2671 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X420 vdd.t2670 vp_p.t329 out_p.t2307 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X421 out_p.t2306 vp_p.t330 vdd.t2669 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X422 out_p.t2305 vp_p.t331 vdd.t2668 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X423 out_p.t63 vp_n.t91 vss.t508 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X424 vdd.t2667 vp_p.t332 out_p.t2304 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X425 vdd.t2666 vp_p.t333 out_p.t2303 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X426 vdd.t2665 vp_p.t334 out_p.t2302 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X427 vdd.t2664 vp_p.t335 out_p.t2301 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X428 out_p.t2300 vp_p.t336 vdd.t2663 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X429 vdd.t2662 vp_p.t337 out_p.t2299 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X430 out_p.t2298 vp_p.t338 vdd.t2661 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X431 vdd.t2660 vp_p.t339 out_p.t2297 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X432 vss.t507 vp_n.t92 out_p.t149 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X433 vdd.t2659 vp_p.t340 out_p.t2296 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X434 out_p.t2290 vp_p.t341 vdd.t2658 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X435 vdd.t2657 vp_p.t342 out_p.t2289 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X436 vss.t506 vp_n.t93 out_p.t121 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X437 out_p.t114 vp_n.t94 vss.t505 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X438 vdd.t2656 vp_p.t343 out_p.t2288 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X439 out_p.t2287 vp_p.t344 vdd.t2655 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X440 out_p.t2286 vp_p.t345 vdd.t2654 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X441 vdd.t2653 vp_p.t346 out_p.t2285 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X442 vdd.t2652 vp_p.t347 out_p.t2279 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X443 vss.t504 vp_n.t95 out_p.t109 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X444 out_p.t2278 vp_p.t348 vdd.t2651 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X445 vdd.t2650 vp_p.t349 out_p.t2277 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X446 out_p.t2276 vp_p.t350 vdd.t2649 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X447 out_p.t107 vp_n.t96 vss.t503 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X448 out_p.t2275 vp_p.t351 vdd.t2648 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X449 vdd.t2647 vp_p.t352 out_p.t2274 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X450 vss.t502 vp_n.t97 out_p.t103 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X451 vss.t501 vp_n.t98 out_p.t101 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X452 vdd.t2646 vp_p.t353 out_p.t2268 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X453 out_p.t2267 vp_p.t354 vdd.t2645 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X454 out_p.t98 vp_n.t99 vss.t500 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X455 vdd.t2644 vp_p.t355 out_p.t2266 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X456 vss.t499 vp_n.t100 out_p.t183 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X457 vdd.t2643 vp_p.t356 out_p.t2265 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X458 out_p.t2264 vp_p.t357 vdd.t2642 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X459 out_p.t2263 vp_p.t358 vdd.t2641 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X460 out_p.t147 vp_n.t101 vss.t498 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X461 out_p.t2254 vp_p.t359 vdd.t2640 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X462 vdd.t2639 vp_p.t360 out_p.t2253 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X463 vss.t497 vp_n.t102 out_p.t144 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X464 vdd.t2638 vp_p.t361 out_p.t2252 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X465 out_p.t2251 vp_p.t362 vdd.t2637 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X466 out_p.t134 vp_n.t103 vss.t496 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X467 vss.t495 vp_n.t104 out_p.t124 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X468 vss.t494 vp_n.t105 out_p.t131 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X469 out_p.t137 vp_n.t106 vss.t493 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X470 vdd.t2636 vp_p.t363 out_p.t2250 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X471 out_p.t2249 vp_p.t364 vdd.t2635 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X472 vdd.t2634 vp_p.t365 out_p.t2242 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X473 vdd.t2633 vp_p.t366 out_p.t2241 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X474 vdd.t2632 vp_p.t367 out_p.t2240 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X475 out_p.t2239 vp_p.t368 vdd.t2631 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X476 out_p.t2238 vp_p.t369 vdd.t2630 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X477 out_p.t2237 vp_p.t370 vdd.t2629 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X478 vss.t492 vp_n.t107 out_p.t140 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X479 out_p.t2231 vp_p.t371 vdd.t2628 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X480 vss.t491 vp_n.t108 out_p.t3490 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X481 vdd.t2627 vp_p.t372 out_p.t2230 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X482 out_p.t2229 vp_p.t373 vdd.t2626 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X483 vdd.t2625 vp_p.t374 out_p.t2228 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X484 vdd.t2624 vp_p.t375 out_p.t2227 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X485 out_p.t2226 vp_p.t376 vdd.t2623 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X486 out_p.t2218 vp_p.t377 vdd.t2622 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X487 vdd.t2621 vp_p.t378 out_p.t2217 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X488 out_p.t3497 vp_n.t109 vss.t490 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X489 vss.t489 vp_n.t110 out_p.t3494 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X490 vdd.t2620 vp_p.t379 out_p.t2216 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X491 vdd.t2619 vp_p.t380 out_p.t2215 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X492 out_p.t2214 vp_p.t381 vdd.t2618 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X493 out_p.t2213 vp_p.t382 vdd.t2617 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X494 out_p.t3455 vp_n.t111 vss.t488 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X495 vdd.t2616 vp_p.t383 out_p.t2205 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X496 vss.t487 vp_n.t112 out_p.t322 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X497 out_p.t2204 vp_p.t384 vdd.t2615 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X498 out_p.t13 vp_n.t113 vss.t486 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X499 out_p.t2203 vp_p.t385 vdd.t2614 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X500 vdd.t2613 vp_p.t386 out_p.t2202 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X501 vdd.t2612 vp_p.t387 out_p.t2201 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X502 vdd.t2611 vp_p.t388 out_p.t2200 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X503 vss.t485 vp_n.t114 out_p.t11 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X504 vdd.t2610 vp_p.t389 out_p.t2193 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X505 vdd.t2609 vp_p.t390 out_p.t2192 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X506 vdd.t2608 vp_p.t391 out_p.t2191 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X507 vdd.t2607 vp_p.t392 out_p.t2190 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X508 vss.t484 vp_n.t115 out_p.t8 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X509 vdd.t2606 vp_p.t393 out_p.t2189 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X510 out_p.t2188 vp_p.t394 vdd.t2605 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X511 vdd.t2604 vp_p.t395 out_p.t2182 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X512 out_p.t2181 vp_p.t396 vdd.t2603 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X513 out_p.t2180 vp_p.t397 vdd.t2602 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X514 out_p.t165 vp_n.t116 vss.t483 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X515 vss.t482 vp_n.t117 out_p.t164 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X516 out_p.t3 vp_n.t118 vss.t481 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X517 out_p.t2179 vp_p.t398 vdd.t2601 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X518 out_p.t2178 vp_p.t399 vdd.t2600 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X519 vss.t480 vp_n.t119 out_p.t1 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X520 vdd.t2599 vp_p.t400 out_p.t2177 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X521 vdd.t2598 vp_p.t401 out_p.t2169 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X522 out_p.t2168 vp_p.t402 vdd.t2597 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X523 out_p.t3487 vp_n.t120 vss.t479 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X524 vdd.t2596 vp_p.t403 out_p.t2167 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X525 vdd.t2595 vp_p.t404 out_p.t2166 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X526 out_p.t2165 vp_p.t405 vdd.t2594 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X527 out_p.t3486 vp_n.t121 vss.t478 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X528 vss.t477 vp_n.t122 out_p.t3484 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X529 out_p.t3492 vp_n.t123 vss.t476 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X530 vdd.t2593 vp_p.t406 out_p.t2164 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X531 vdd.t2592 vp_p.t407 out_p.t2157 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X532 out_p.t2156 vp_p.t408 vdd.t2591 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X533 vss.t475 vp_n.t124 out_p.t3541 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X534 vss.t474 vp_n.t125 out_p.t3539 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X535 vdd.t2590 vp_p.t409 out_p.t2155 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X536 out_p.t2154 vp_p.t410 vdd.t2589 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X537 out_p.t2153 vp_p.t411 vdd.t2588 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X538 vss.t473 vp_n.t126 out_p.t3546 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X539 out_p.t2152 vp_p.t412 vdd.t2587 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X540 vdd.t2586 vp_p.t413 out_p.t2146 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X541 out_p.t2145 vp_p.t414 vdd.t2585 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X542 out_p.t3544 vp_n.t127 vss.t472 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X543 out_p.t2144 vp_p.t415 vdd.t2584 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X544 out_p.t2143 vp_p.t416 vdd.t2583 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X545 vss.t471 vp_n.t128 out_p.t187 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X546 out_p.t185 vp_n.t129 vss.t470 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X547 out_p.t156 vp_n.t130 vss.t469 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X548 out_p.t2142 vp_p.t417 vdd.t2582 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X549 vdd.t2581 vp_p.t418 out_p.t2141 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X550 vdd.t2580 vp_p.t419 out_p.t2134 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X551 vss.t468 vp_n.t131 out_p.t153 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X552 out_p.t2133 vp_p.t420 vdd.t2579 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X553 vdd.t2578 vp_p.t421 out_p.t2132 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X554 out_p.t419 vp_n.t132 vss.t467 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X555 vss.t466 vp_n.t133 out_p.t3550 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X556 vdd.t2577 vp_p.t422 out_p.t2131 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X557 vdd.t2576 vp_p.t423 out_p.t2130 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X558 out_p.t2129 vp_p.t424 vdd.t2575 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X559 out_p.t2123 vp_p.t425 vdd.t2574 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X560 out_p.t2122 vp_p.t426 vdd.t2573 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X561 out_p.t2121 vp_p.t427 vdd.t2572 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X562 out_p.t2120 vp_p.t428 vdd.t2571 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X563 vdd.t2570 vp_p.t429 out_p.t2119 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X564 out_p.t3548 vp_n.t134 vss.t465 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X565 vdd.t2569 vp_p.t430 out_p.t2118 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X566 vss.t464 vp_n.t135 out_p.t3556 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X567 out_p.t2110 vp_p.t431 vdd.t2568 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X568 out_p.t2109 vp_p.t432 vdd.t2567 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X569 out_p.t2108 vp_p.t433 vdd.t2566 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X570 vdd.t2565 vp_p.t434 out_p.t2107 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X571 out_p.t2106 vp_p.t435 vdd.t2564 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X572 vdd.t2563 vp_p.t436 out_p.t2105 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X573 vdd.t2562 vp_p.t437 out_p.t2099 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X574 out_p.t2098 vp_p.t438 vdd.t2561 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X575 out_p.t2097 vp_p.t439 vdd.t2560 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X576 out_p.t2096 vp_p.t440 vdd.t2559 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X577 vdd.t2558 vp_p.t441 out_p.t2095 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X578 out_p.t2094 vp_p.t442 vdd.t2557 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X579 out_p.t2087 vp_p.t443 vdd.t2556 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X580 vss.t463 vp_n.t136 out_p.t3554 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X581 out_p.t2086 vp_p.t444 vdd.t2555 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X582 vdd.t2554 vp_p.t445 out_p.t2085 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X583 vdd.t2553 vp_p.t446 out_p.t2084 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X584 out_p.t3535 vp_n.t137 vss.t462 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X585 vdd.t2552 vp_p.t447 out_p.t2083 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X586 vdd.t2551 vp_p.t448 out_p.t2082 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X587 out_p.t2076 vp_p.t449 vdd.t2550 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X588 vdd.t2549 vp_p.t450 out_p.t2075 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X589 vdd.t2548 vp_p.t451 out_p.t2074 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X590 vdd.t2547 vp_p.t452 out_p.t2073 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X591 vss.t461 vp_n.t138 out_p.t3533 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X592 out_p.t3530 vp_n.t139 vss.t460 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X593 out_p.t2072 vp_p.t453 vdd.t2546 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X594 out_p.t2071 vp_p.t454 vdd.t2545 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X595 vss.t459 vp_n.t140 out_p.t321 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X596 vdd.t2544 vp_p.t455 out_p.t2064 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X597 vdd.t2543 vp_p.t456 out_p.t2063 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X598 vdd.t2542 vp_p.t457 out_p.t2062 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X599 out_p.t2061 vp_p.t458 vdd.t2541 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X600 vdd.t2540 vp_p.t459 out_p.t2060 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X601 vdd.t2539 vp_p.t460 out_p.t2059 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X602 out_p.t2053 vp_p.t461 vdd.t2538 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X603 vdd.t2537 vp_p.t462 out_p.t2052 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X604 vss.t458 vp_n.t141 out_p.t3568 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X605 out_p.t2051 vp_p.t463 vdd.t2536 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X606 out_p.t2050 vp_p.t464 vdd.t2535 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X607 vss.t457 vp_n.t142 out_p.t353 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X608 out_p.t3476 vp_n.t143 vss.t456 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X609 vdd.t2534 vp_p.t465 out_p.t2049 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X610 vdd.t2533 vp_p.t466 out_p.t2048 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X611 vdd.t2532 vp_p.t467 out_p.t2041 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X612 vdd.t2531 vp_p.t468 out_p.t2040 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X613 out_p.t2039 vp_p.t469 vdd.t2530 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X614 vss.t455 vp_n.t144 out_p.t3474 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X615 out_p.t2038 vp_p.t470 vdd.t2529 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X616 vdd.t2528 vp_p.t471 out_p.t2037 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X617 out_p.t2036 vp_p.t472 vdd.t2527 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X618 out_p.t2030 vp_p.t473 vdd.t2526 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X619 vdd.t2525 vp_p.t474 out_p.t2029 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X620 vss.t454 vp_n.t145 out_p.t3459 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X621 vdd.t2524 vp_p.t475 out_p.t2028 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X622 out_p.t2027 vp_p.t476 vdd.t2523 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X623 out_p.t3458 vp_n.t146 vss.t453 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X624 vdd.t2522 vp_p.t477 out_p.t2026 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X625 out_p.t2025 vp_p.t478 vdd.t2521 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X626 out_p.t2018 vp_p.t479 vdd.t2520 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X627 out_p.t421 vp_n.t147 vss.t452 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X628 out_p.t2017 vp_p.t480 vdd.t2519 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X629 vdd.t2518 vp_p.t481 out_p.t2016 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X630 out_p.t2015 vp_p.t482 vdd.t2517 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X631 out_p.t2014 vp_p.t483 vdd.t2516 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X632 vss.t451 vp_n.t148 out_p.t175 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X633 out_p.t2013 vp_p.t484 vdd.t2515 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X634 out_p.t2007 vp_p.t485 vdd.t2514 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X635 vss.t450 vp_n.t149 out_p.t3599 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X636 vdd.t2513 vp_p.t486 out_p.t2006 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X637 vdd.t2512 vp_p.t487 out_p.t2005 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X638 out_p.t2004 vp_p.t488 vdd.t2511 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X639 vdd.t2510 vp_p.t489 out_p.t2003 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X640 out_p.t2002 vp_p.t490 vdd.t2509 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X641 out_p.t1995 vp_p.t491 vdd.t2508 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X642 out_p.t3597 vp_n.t150 vss.t449 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X643 vss.t448 vp_n.t151 out_p.t3503 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X644 out_p.t1994 vp_p.t492 vdd.t2507 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X645 out_p.t1993 vp_p.t493 vdd.t2506 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X646 vdd.t2505 vp_p.t494 out_p.t1992 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X647 out_p.t1991 vp_p.t495 vdd.t2504 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X648 vdd.t2503 vp_p.t496 out_p.t1990 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X649 vss.t447 vp_n.t152 out_p.t3463 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X650 vdd.t2502 vp_p.t497 out_p.t1984 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X651 vdd.t2501 vp_p.t498 out_p.t1983 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X652 out_p.t1982 vp_p.t499 vdd.t2500 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X653 vdd.t2499 vp_p.t500 out_p.t1981 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X654 vss.t446 vp_n.t153 out_p.t257 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X655 out_p.t1980 vp_p.t501 vdd.t2498 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X656 out_p.t1979 vp_p.t502 vdd.t2497 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X657 vdd.t2496 vp_p.t503 out_p.t1972 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X658 out_p.t3461 vp_n.t154 vss.t445 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X659 out_p.t3570 vp_n.t155 vss.t444 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X660 out_p.t1971 vp_p.t504 vdd.t2495 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X661 vdd.t2494 vp_p.t505 out_p.t1970 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X662 vdd.t2493 vp_p.t506 out_p.t1969 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X663 out_p.t1968 vp_p.t507 vdd.t2492 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X664 vdd.t2491 vp_p.t508 out_p.t1967 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X665 vdd.t2490 vp_p.t509 out_p.t1961 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X666 out_p.t1960 vp_p.t510 vdd.t2489 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X667 out_p.t339 vp_n.t156 vss.t443 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X668 vdd.t2488 vp_p.t511 out_p.t1959 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X669 out_p.t1958 vp_p.t512 vdd.t2487 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X670 out_p.t1957 vp_p.t513 vdd.t2486 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X671 out_p.t1956 vp_p.t514 vdd.t2485 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X672 vdd.t2484 vp_p.t515 out_p.t1948 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X673 vss.t442 vp_n.t157 out_p.t340 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X674 vdd.t2483 vp_p.t516 out_p.t1947 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X675 out_p.t1946 vp_p.t517 vdd.t2482 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X676 vdd.t2481 vp_p.t518 out_p.t1945 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X677 vss.t441 vp_n.t158 out_p.t348 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X678 out_p.t1944 vp_p.t519 vdd.t2480 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X679 vdd.t2479 vp_p.t520 out_p.t1943 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X680 out_p.t1936 vp_p.t521 vdd.t2478 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X681 out_p.t1935 vp_p.t522 vdd.t2477 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X682 out_p.t1934 vp_p.t523 vdd.t2476 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X683 vdd.t2475 vp_p.t524 out_p.t1933 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X684 out_p.t1932 vp_p.t525 vdd.t2474 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X685 vss.t440 vp_n.t159 out_p.t344 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X686 out_p.t1931 vp_p.t526 vdd.t2473 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X687 out_p.t1925 vp_p.t527 vdd.t2472 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X688 out_p.t1924 vp_p.t528 vdd.t2471 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X689 out_p.t1923 vp_p.t529 vdd.t2470 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X690 vdd.t2469 vp_p.t530 out_p.t1922 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X691 out_p.t1921 vp_p.t531 vdd.t2468 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X692 out_p.t1920 vp_p.t532 vdd.t2467 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X693 out_p.t1913 vp_p.t533 vdd.t2466 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X694 out_p.t1912 vp_p.t534 vdd.t2465 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X695 out_p.t1911 vp_p.t535 vdd.t2464 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X696 out_p.t1910 vp_p.t536 vdd.t2463 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X697 out_p.t352 vp_n.t160 vss.t439 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X698 out_p.t1909 vp_p.t537 vdd.t2462 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X699 vss.t438 vp_n.t161 out_p.t180 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X700 vdd.t2461 vp_p.t538 out_p.t1908 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X701 vdd.t2460 vp_p.t539 out_p.t1902 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X702 vdd.t2459 vp_p.t540 out_p.t1901 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X703 out_p.t178 vp_n.t162 vss.t437 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X704 vdd.t2458 vp_p.t541 out_p.t1900 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X705 out_p.t1899 vp_p.t542 vdd.t2457 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X706 vss.t436 vp_n.t163 out_p.t177 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X707 vss.t435 vp_n.t164 out_p.t294 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X708 out_p.t1898 vp_p.t543 vdd.t2456 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X709 out_p.t1897 vp_p.t544 vdd.t2455 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X710 vdd.t2454 vp_p.t545 out_p.t1890 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X711 vdd.t2453 vp_p.t546 out_p.t1889 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X712 out_p.t1888 vp_p.t547 vdd.t2452 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X713 out_p.t1887 vp_p.t548 vdd.t2451 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X714 vdd.t2450 vp_p.t549 out_p.t1886 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X715 out_p.t310 vp_n.t165 vss.t434 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X716 vss.t433 vp_n.t166 out_p.t311 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X717 out_p.t1885 vp_p.t550 vdd.t2449 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X718 vdd.t2448 vp_p.t551 out_p.t1879 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X719 out_p.t1878 vp_p.t552 vdd.t2447 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X720 vdd.t2446 vp_p.t553 out_p.t1877 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X721 out_p.t1876 vp_p.t554 vdd.t2445 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X722 vdd.t2444 vp_p.t555 out_p.t1875 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X723 vss.t432 vp_n.t167 out_p.t312 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X724 out_p.t1874 vp_p.t556 vdd.t2443 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X725 out_p.t1867 vp_p.t557 vdd.t2442 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X726 out_p.t1866 vp_p.t558 vdd.t2441 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X727 out_p.t313 vp_n.t168 vss.t431 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X728 vdd.t2440 vp_p.t559 out_p.t1865 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X729 out_p.t1864 vp_p.t560 vdd.t2439 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X730 vss.t430 vp_n.t169 out_p.t328 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X731 vdd.t2438 vp_p.t561 out_p.t1863 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X732 out_p.t1862 vp_p.t562 vdd.t2437 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X733 out_p.t1856 vp_p.t563 vdd.t2436 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X734 out_p.t1855 vp_p.t564 vdd.t2435 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X735 vss.t429 vp_n.t170 out_p.t327 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X736 vdd.t2434 vp_p.t565 out_p.t1854 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X737 vdd.t2433 vp_p.t566 out_p.t1853 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X738 vdd.t2432 vp_p.t567 out_p.t1852 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X739 out_p.t333 vp_n.t171 vss.t428 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X740 out_p.t1851 vp_p.t568 vdd.t2431 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X741 out_p.t1843 vp_p.t569 vdd.t2430 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X742 out_p.t1842 vp_p.t570 vdd.t2429 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X743 out_p.t1841 vp_p.t571 vdd.t2428 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X744 vdd.t2427 vp_p.t572 out_p.t1840 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X745 out_p.t1839 vp_p.t573 vdd.t2426 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X746 vdd.t2425 vp_p.t574 out_p.t1838 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X747 out_p.t1831 vp_p.t575 vdd.t2424 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X748 vdd.t2423 vp_p.t576 out_p.t1830 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X749 out_p.t1829 vp_p.t577 vdd.t2422 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X750 out_p.t1828 vp_p.t578 vdd.t2421 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X751 vdd.t2420 vp_p.t579 out_p.t1827 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X752 out_p.t1826 vp_p.t580 vdd.t2419 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X753 out_p.t1820 vp_p.t581 vdd.t2418 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X754 vdd.t2417 vp_p.t582 out_p.t1819 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X755 vdd.t2416 vp_p.t583 out_p.t1818 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X756 vss.t427 vp_n.t172 out_p.t270 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X757 out_p.t273 vp_n.t173 vss.t426 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X758 vdd.t2415 vp_p.t584 out_p.t1817 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X759 out_p.t1816 vp_p.t585 vdd.t2414 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X760 vdd.t2413 vp_p.t586 out_p.t1815 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X761 out_p.t1808 vp_p.t587 vdd.t2412 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X762 vdd.t2411 vp_p.t588 out_p.t1807 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X763 vdd.t2410 vp_p.t589 out_p.t1806 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X764 vdd.t2409 vp_p.t590 out_p.t1805 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X765 out_p.t1804 vp_p.t591 vdd.t2408 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X766 out_p.t1803 vp_p.t592 vdd.t2407 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X767 out_p.t275 vp_n.t174 vss.t425 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X768 out_p.t1797 vp_p.t593 vdd.t2406 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X769 vss.t424 vp_n.t175 out_p.t279 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X770 out_p.t282 vp_n.t176 vss.t423 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X771 vdd.t2405 vp_p.t594 out_p.t1796 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X772 out_p.t1795 vp_p.t595 vdd.t2404 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X773 out_p.t1794 vp_p.t596 vdd.t2403 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X774 vdd.t2402 vp_p.t597 out_p.t1793 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X775 out_p.t285 vp_n.t177 vss.t422 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X776 vdd.t2401 vp_p.t598 out_p.t1792 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X777 vdd.t2400 vp_p.t599 out_p.t1784 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X778 out_p.t1783 vp_p.t600 vdd.t2399 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X779 out_p.t1782 vp_p.t601 vdd.t2398 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X780 out_p.t1781 vp_p.t602 vdd.t2397 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X781 vdd.t2396 vp_p.t603 out_p.t1780 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X782 out_p.t1779 vp_p.t604 vdd.t2395 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X783 out_p.t288 vp_n.t178 vss.t421 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X784 vdd.t2394 vp_p.t605 out_p.t1773 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X785 out_p.t1772 vp_p.t606 vdd.t2393 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X786 vss.t420 vp_n.t179 out_p.t290 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X787 out_p.t1771 vp_p.t607 vdd.t2392 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X788 out_p.t1770 vp_p.t608 vdd.t2391 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X789 vss.t419 vp_n.t180 out_p.t3528 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X790 out_p.t3525 vp_n.t181 vss.t418 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X791 out_p.t1769 vp_p.t609 vdd.t2390 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X792 out_p.t1768 vp_p.t610 vdd.t2389 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X793 vdd.t2388 vp_p.t611 out_p.t1761 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X794 vdd.t2387 vp_p.t612 out_p.t1760 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X795 out_p.t3526 vp_n.t182 vss.t417 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X796 out_p.t1759 vp_p.t613 vdd.t2386 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X797 out_p.t3521 vp_n.t183 vss.t416 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X798 out_p.t1758 vp_p.t614 vdd.t2385 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X799 vss.t415 vp_n.t184 out_p.t3522 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X800 vdd.t2384 vp_p.t615 out_p.t1757 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X801 vdd.t2383 vp_p.t616 out_p.t1756 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X802 out_p.t1750 vp_p.t617 vdd.t2382 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X803 vss.t414 vp_n.t185 out_p.t3516 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X804 out_p.t1749 vp_p.t618 vdd.t2381 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X805 vdd.t2380 vp_p.t619 out_p.t1748 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X806 out_p.t1747 vp_p.t620 vdd.t2379 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X807 out_p.t1746 vp_p.t621 vdd.t2378 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X808 out_p.t1745 vp_p.t622 vdd.t2377 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X809 out_p.t1737 vp_p.t623 vdd.t2376 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X810 out_p.t1736 vp_p.t624 vdd.t2375 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X811 out_p.t1735 vp_p.t625 vdd.t2374 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X812 out_p.t1734 vp_p.t626 vdd.t2373 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X813 out_p.t1733 vp_p.t627 vdd.t2372 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X814 out_p.t3509 vp_n.t186 vss.t413 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X815 out_p.t1732 vp_p.t628 vdd.t2371 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X816 vdd.t2370 vp_p.t629 out_p.t1725 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X817 out_p.t1724 vp_p.t630 vdd.t2369 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X818 vdd.t2368 vp_p.t631 out_p.t1723 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X819 out_p.t1722 vp_p.t632 vdd.t2367 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X820 vss.t412 vp_n.t187 out_p.t3510 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X821 vdd.t2366 vp_p.t633 out_p.t1721 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X822 out_p.t1720 vp_p.t634 vdd.t2365 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X823 vdd.t2364 vp_p.t635 out_p.t1714 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X824 out_p.t1713 vp_p.t636 vdd.t2363 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X825 vdd.t2362 vp_p.t637 out_p.t1712 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X826 vdd.t2361 vp_p.t638 out_p.t1711 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X827 out_p.t1710 vp_p.t639 vdd.t2360 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X828 vdd.t2359 vp_p.t640 out_p.t1709 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X829 vdd.t2358 vp_p.t641 out_p.t1702 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X830 out_p.t1701 vp_p.t642 vdd.t2357 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X831 vdd.t2356 vp_p.t643 out_p.t1700 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X832 out_p.t1699 vp_p.t644 vdd.t2355 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X833 vdd.t2354 vp_p.t645 out_p.t1698 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X834 vdd.t2353 vp_p.t646 out_p.t1697 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X835 vdd.t2352 vp_p.t647 out_p.t1691 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X836 out_p.t1690 vp_p.t648 vdd.t2351 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X837 out_p.t1689 vp_p.t649 vdd.t2350 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X838 out_p.t1688 vp_p.t650 vdd.t2349 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X839 out_p.t1687 vp_p.t651 vdd.t2348 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X840 vdd.t2347 vp_p.t652 out_p.t1686 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X841 out_p.t3491 vp_n.t188 vss.t411 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X842 out_p.t1679 vp_p.t653 vdd.t2346 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X843 vss.t410 vp_n.t189 out_p.t3488 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X844 out_p.t1678 vp_p.t654 vdd.t2345 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X845 vss.t409 vp_n.t190 out_p.t3495 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X846 out_p.t1677 vp_p.t655 vdd.t2344 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X847 vdd.t2343 vp_p.t656 out_p.t1676 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X848 out_p.t1675 vp_p.t657 vdd.t2342 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X849 vdd.t2341 vp_p.t658 out_p.t1674 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X850 out_p.t1668 vp_p.t659 vdd.t2340 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X851 vdd.t2339 vp_p.t660 out_p.t1667 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X852 out_p.t1666 vp_p.t661 vdd.t2338 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X853 out_p.t1665 vp_p.t662 vdd.t2337 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X854 out_p.t1664 vp_p.t663 vdd.t2336 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X855 vdd.t2335 vp_p.t664 out_p.t1663 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X856 out_p.t1655 vp_p.t665 vdd.t2334 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X857 vdd.t2333 vp_p.t666 out_p.t1654 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X858 vss.t408 vp_n.t191 out_p.t3493 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X859 vdd.t2332 vp_p.t667 out_p.t1653 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X860 out_p.t1652 vp_p.t668 vdd.t2331 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X861 vss.t407 vp_n.t192 out_p.t3454 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X862 out_p.t1651 vp_p.t669 vdd.t2330 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X863 vdd.t2329 vp_p.t670 out_p.t1650 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X864 out_p.t1644 vp_p.t671 vdd.t2328 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X865 out_p.t1643 vp_p.t672 vdd.t2327 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X866 out_p.t1642 vp_p.t673 vdd.t2326 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X867 out_p.t1641 vp_p.t674 vdd.t2325 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X868 vdd.t2324 vp_p.t675 out_p.t1640 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X869 vdd.t2323 vp_p.t676 out_p.t1639 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X870 out_p.t3595 vp_n.t193 vss.t406 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X871 out_p.t1632 vp_p.t677 vdd.t2322 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X872 out_p.t1631 vp_p.t678 vdd.t2321 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X873 out_p.t1630 vp_p.t679 vdd.t2320 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X874 vdd.t2319 vp_p.t680 out_p.t1629 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X875 vss.t405 vp_n.t194 out_p.t189 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X876 vdd.t2318 vp_p.t681 out_p.t1628 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X877 out_p.t1627 vp_p.t682 vdd.t2317 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X878 out_p.t1621 vp_p.t683 vdd.t2316 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X879 vdd.t2315 vp_p.t684 out_p.t1620 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X880 vdd.t2314 vp_p.t685 out_p.t1619 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X881 out_p.t1618 vp_p.t686 vdd.t2313 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X882 vdd.t2312 vp_p.t687 out_p.t1617 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X883 out_p.t1616 vp_p.t688 vdd.t2311 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X884 out_p.t1613 vp_p.t689 vdd.t2310 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X885 vdd.t2309 vp_p.t690 out_p.t1612 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X886 out_p.t1611 vp_p.t691 vdd.t2308 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X887 vdd.t2307 vp_p.t692 out_p.t1610 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X888 out_p.t1609 vp_p.t693 vdd.t2306 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X889 out_p.t1608 vp_p.t694 vdd.t2305 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X890 out_p.t1602 vp_p.t695 vdd.t2304 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X891 out_p.t1601 vp_p.t696 vdd.t2303 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X892 vdd.t2302 vp_p.t697 out_p.t1600 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X893 vdd.t2301 vp_p.t698 out_p.t1599 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X894 vdd.t2300 vp_p.t699 out_p.t1598 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X895 out_p.t1597 vp_p.t700 vdd.t2299 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X896 vdd.t2298 vp_p.t701 out_p.t1590 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X897 out_p.t1589 vp_p.t702 vdd.t2297 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X898 vdd.t2296 vp_p.t703 out_p.t1588 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X899 vdd.t2295 vp_p.t704 out_p.t1587 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X900 out_p.t1586 vp_p.t705 vdd.t2294 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X901 vdd.t2293 vp_p.t706 out_p.t1585 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X902 vdd.t2292 vp_p.t707 out_p.t1579 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X903 out_p.t1578 vp_p.t708 vdd.t2291 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X904 out_p.t1577 vp_p.t709 vdd.t2290 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X905 out_p.t3527 vp_n.t195 vss.t404 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X906 out_p.t1576 vp_p.t710 vdd.t2289 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X907 vdd.t2288 vp_p.t711 out_p.t1575 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X908 out_p.t1574 vp_p.t712 vdd.t2287 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X909 vdd.t2286 vp_p.t713 out_p.t1567 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X910 vdd.t2285 vp_p.t714 out_p.t1566 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X911 out_p.t1565 vp_p.t715 vdd.t2284 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X912 vdd.t2283 vp_p.t716 out_p.t1564 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X913 out_p.t1563 vp_p.t717 vdd.t2282 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X914 vdd.t2281 vp_p.t718 out_p.t1562 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X915 out_p.t355 vp_n.t196 vss.t403 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X916 out_p.t1556 vp_p.t719 vdd.t2280 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X917 vdd.t2279 vp_p.t720 out_p.t1555 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X918 vdd.t2278 vp_p.t721 out_p.t1554 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X919 vdd.t2277 vp_p.t722 out_p.t1553 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X920 out_p.t1552 vp_p.t723 vdd.t2276 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X921 out_p.t1551 vp_p.t724 vdd.t2275 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X922 vss.t402 vp_n.t197 out_p.t154 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X923 vdd.t2274 vp_p.t725 out_p.t1544 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X924 vdd.t2273 vp_p.t726 out_p.t1543 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X925 vdd.t2272 vp_p.t727 out_p.t1542 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X926 vdd.t2271 vp_p.t728 out_p.t1541 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X927 out_p.t1540 vp_p.t729 vdd.t2270 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X928 out_p.t1539 vp_p.t730 vdd.t2269 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X929 vdd.t2268 vp_p.t731 out_p.t1533 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X930 out_p.t1532 vp_p.t732 vdd.t2267 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X931 vdd.t2266 vp_p.t733 out_p.t1531 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X932 vdd.t2265 vp_p.t734 out_p.t1530 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X933 vdd.t2264 vp_p.t735 out_p.t1529 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X934 vdd.t2263 vp_p.t736 out_p.t1528 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X935 out_p.t1520 vp_p.t737 vdd.t2262 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X936 vdd.t2261 vp_p.t738 out_p.t1519 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X937 vdd.t2260 vp_p.t739 out_p.t1518 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X938 vdd.t2259 vp_p.t740 out_p.t1517 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X939 out_p.t1516 vp_p.t741 vdd.t2258 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X940 out_p.t1515 vp_p.t742 vdd.t2257 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X941 out_p.t1507 vp_p.t743 vdd.t2256 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X942 out_p.t1506 vp_p.t744 vdd.t2255 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X943 out_p.t1505 vp_p.t745 vdd.t2254 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X944 vdd.t2253 vp_p.t746 out_p.t1504 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X945 vdd.t2252 vp_p.t747 out_p.t1503 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X946 vdd.t2251 vp_p.t748 out_p.t1502 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X947 out_p.t1496 vp_p.t749 vdd.t2250 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X948 vdd.t2249 vp_p.t750 out_p.t1495 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X949 vdd.t2248 vp_p.t751 out_p.t1494 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X950 vdd.t2247 vp_p.t752 out_p.t1493 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X951 vdd.t2246 vp_p.t753 out_p.t1492 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X952 vdd.t2245 vp_p.t754 out_p.t1491 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X953 out_p.t1490 vp_p.t755 vdd.t2244 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X954 vdd.t2243 vp_p.t756 out_p.t1489 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X955 out_p.t1488 vp_p.t757 vdd.t2242 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X956 vdd.t2241 vp_p.t758 out_p.t1487 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X957 out_p.t1486 vp_p.t759 vdd.t2240 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X958 out_p.t1485 vp_p.t760 vdd.t2239 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X959 out_p.t1479 vp_p.t761 vdd.t2238 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X960 vdd.t2237 vp_p.t762 out_p.t1478 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X961 vdd.t2236 vp_p.t763 out_p.t1477 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X962 out_p.t1476 vp_p.t764 vdd.t2235 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X963 out_p.t1475 vp_p.t765 vdd.t2234 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X964 vdd.t2233 vp_p.t766 out_p.t1474 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X965 out_p.t1466 vp_p.t767 vdd.t2232 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X966 vdd.t2231 vp_p.t768 out_p.t1465 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X967 out_p.t1464 vp_p.t769 vdd.t2230 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X968 vdd.t2229 vp_p.t770 out_p.t1463 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X969 out_p.t1462 vp_p.t771 vdd.t2228 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X970 vdd.t2227 vp_p.t772 out_p.t1461 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X971 out_p.t1455 vp_p.t773 vdd.t2226 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X972 out_p.t1454 vp_p.t774 vdd.t2225 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X973 out_p.t1453 vp_p.t775 vdd.t2224 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X974 vdd.t2223 vp_p.t776 out_p.t1452 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X975 vdd.t2222 vp_p.t777 out_p.t1451 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X976 out_p.t1450 vp_p.t778 vdd.t2221 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X977 vdd.t2220 vp_p.t779 out_p.t1443 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X978 out_p.t1442 vp_p.t780 vdd.t2219 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X979 vdd.t2218 vp_p.t781 out_p.t1441 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X980 out_p.t1440 vp_p.t782 vdd.t2217 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X981 out_p.t1439 vp_p.t783 vdd.t2216 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X982 vdd.t2215 vp_p.t784 out_p.t1438 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X983 out_p.t1431 vp_p.t785 vdd.t2214 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X984 vdd.t2213 vp_p.t786 out_p.t1430 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X985 vdd.t2212 vp_p.t787 out_p.t1429 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X986 vdd.t2211 vp_p.t788 out_p.t1428 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X987 vdd.t2210 vp_p.t789 out_p.t1427 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X988 vdd.t2209 vp_p.t790 out_p.t1426 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X989 out_p.t1424 vp_p.t791 vdd.t2208 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X990 out_p.t1423 vp_p.t792 vdd.t2207 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X991 vdd.t2206 vp_p.t793 out_p.t1422 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X992 vdd.t2205 vp_p.t794 out_p.t1421 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X993 out_p.t1420 vp_p.t795 vdd.t2204 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X994 vdd.t2203 vp_p.t796 out_p.t1419 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X995 vdd.t2202 vp_p.t797 out_p.t1413 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X996 vdd.t2201 vp_p.t798 out_p.t1412 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X997 out_p.t1411 vp_p.t799 vdd.t2200 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X998 vdd.t2199 vp_p.t800 out_p.t1410 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X999 out_p.t1409 vp_p.t801 vdd.t2198 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1000 vdd.t2197 vp_p.t802 out_p.t1408 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1001 vdd.t2196 vp_p.t803 out_p.t1400 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1002 vdd.t2195 vp_p.t804 out_p.t1399 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1003 out_p.t1398 vp_p.t805 vdd.t2194 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1004 vdd.t2193 vp_p.t806 out_p.t1397 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1005 out_p.t1396 vp_p.t807 vdd.t2192 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1006 vdd.t2191 vp_p.t808 out_p.t1395 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1007 out_p.t1389 vp_p.t809 vdd.t2190 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1008 out_p.t1388 vp_p.t810 vdd.t2189 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1009 vdd.t2188 vp_p.t811 out_p.t1387 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1010 vdd.t2187 vp_p.t812 out_p.t1386 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1011 out_p.t1385 vp_p.t813 vdd.t2186 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1012 out_p.t1384 vp_p.t814 vdd.t2185 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1013 out_p.t1382 vp_p.t815 vdd.t2184 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1014 out_p.t1381 vp_p.t816 vdd.t2183 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1015 out_p.t1380 vp_p.t817 vdd.t2182 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1016 vdd.t2181 vp_p.t818 out_p.t1379 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1017 vdd.t2180 vp_p.t819 out_p.t1378 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1018 vdd.t2179 vp_p.t820 out_p.t1377 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1019 out_p.t1371 vp_p.t821 vdd.t2178 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1020 vdd.t2177 vp_p.t822 out_p.t1370 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1021 vdd.t2176 vp_p.t823 out_p.t1369 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1022 vdd.t2175 vp_p.t824 out_p.t1368 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1023 out_p.t1367 vp_p.t825 vdd.t2174 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1024 vdd.t2173 vp_p.t826 out_p.t1366 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1025 out_p.t2506 vp_p.t827 vdd.t2172 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1026 out_p.t2505 vp_p.t828 vdd.t2171 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1027 out_p.t2504 vp_p.t829 vdd.t2170 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1028 out_p.t2503 vp_p.t830 vdd.t2169 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1029 vdd.t2168 vp_p.t831 out_p.t2502 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1030 vdd.t2167 vp_p.t832 out_p.t2511 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1031 vdd.t2166 vp_p.t833 out_p.t2510 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1032 vdd.t2165 vp_p.t834 out_p.t2509 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1033 vdd.t2164 vp_p.t835 out_p.t2508 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1034 out_p.t2507 vp_p.t836 vdd.t2163 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1035 vdd.t2162 vp_p.t837 out_p.t1437 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1036 out_p.t1436 vp_p.t838 vdd.t2161 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1037 out_p.t1435 vp_p.t839 vdd.t2160 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1038 vdd.t2159 vp_p.t840 out_p.t1434 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1039 vdd.t2158 vp_p.t841 out_p.t1433 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1040 vdd.t2157 vp_p.t842 out_p.t2467 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1041 out_p.t2466 vp_p.t843 vdd.t2156 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1042 out_p.t2465 vp_p.t844 vdd.t2155 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1043 out_p.t2464 vp_p.t845 vdd.t2154 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1044 out_p.t2419 vp_p.t846 vdd.t2153 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1045 vdd.t2152 vp_p.t847 out_p.t2418 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1046 out_p.t2417 vp_p.t848 vdd.t2151 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1047 vdd.t2150 vp_p.t849 out_p.t2416 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1048 out_p.t2392 vp_p.t850 vdd.t2149 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1049 out_p.t2391 vp_p.t851 vdd.t2148 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1050 vdd.t2147 vp_p.t852 out_p.t2390 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1051 vdd.t2146 vp_p.t853 out_p.t2389 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1052 vdd.t2145 vp_p.t854 out_p.t2373 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1053 vdd.t2144 vp_p.t855 out_p.t2372 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1054 out_p.t2371 vp_p.t856 vdd.t2143 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1055 vdd.t2142 vp_p.t857 out_p.t2370 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1056 out_p.t2356 vp_p.t858 vdd.t2141 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1057 vdd.t2140 vp_p.t859 out_p.t2355 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1058 out_p.t2354 vp_p.t860 vdd.t2139 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1059 out_p.t2353 vp_p.t861 vdd.t2138 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1060 out_p.t2329 vp_p.t862 vdd.t2137 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1061 vdd.t2136 vp_p.t863 out_p.t2328 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1062 out_p.t2327 vp_p.t864 vdd.t2135 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1063 out_p.t2326 vp_p.t865 vdd.t2134 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1064 vdd.t2133 vp_p.t866 out_p.t2312 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1065 out_p.t2311 vp_p.t867 vdd.t2132 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1066 out_p.t2310 vp_p.t868 vdd.t2131 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1067 out_p.t2309 vp_p.t869 vdd.t2130 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1068 out_p.t2295 vp_p.t870 vdd.t2129 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1069 vdd.t2128 vp_p.t871 out_p.t2294 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1070 out_p.t2293 vp_p.t872 vdd.t2127 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1071 out_p.t2292 vp_p.t873 vdd.t2126 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1072 vdd.t2125 vp_p.t874 out_p.t2273 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1073 vdd.t2124 vp_p.t875 out_p.t2272 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1074 out_p.t2271 vp_p.t876 vdd.t2123 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1075 out_p.t2270 vp_p.t877 vdd.t2122 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1076 vdd.t2121 vp_p.t878 out_p.t2236 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1077 vdd.t2120 vp_p.t879 out_p.t2235 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1078 vdd.t2119 vp_p.t880 out_p.t2234 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1079 vdd.t2118 vp_p.t881 out_p.t2233 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1080 vdd.t2117 vp_p.t882 out_p.t2187 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1081 vdd.t2116 vp_p.t883 out_p.t2186 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1082 out_p.t2185 vp_p.t884 vdd.t2115 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1083 vdd.t2114 vp_p.t885 out_p.t2184 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1084 out_p.t2151 vp_p.t886 vdd.t2113 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1085 vdd.t2112 vp_p.t887 out_p.t2150 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1086 vdd.t2111 vp_p.t888 out_p.t2149 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1087 out_p.t2148 vp_p.t889 vdd.t2110 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1088 vdd.t2109 vp_p.t890 out_p.t2128 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1089 vdd.t2108 vp_p.t891 out_p.t2127 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1090 out_p.t2126 vp_p.t892 vdd.t2107 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1091 out_p.t2125 vp_p.t893 vdd.t2106 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1092 vdd.t2105 vp_p.t894 out_p.t2104 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1093 out_p.t2103 vp_p.t895 vdd.t2104 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1094 out_p.t2102 vp_p.t896 vdd.t2103 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1095 vdd.t2102 vp_p.t897 out_p.t2101 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1096 out_p.t2081 vp_p.t898 vdd.t2101 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1097 vss.t401 vp_n.t198 out_p.t152 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1098 vdd.t2100 vp_p.t899 out_p.t2080 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1099 vdd.t2099 vp_p.t900 out_p.t2079 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1100 vdd.t2098 vp_p.t901 out_p.t2078 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1101 out_p.t2058 vp_p.t902 vdd.t2097 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1102 vdd.t2096 vp_p.t903 out_p.t2057 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1103 vdd.t2095 vp_p.t904 out_p.t2056 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1104 vdd.t2094 vp_p.t905 out_p.t2055 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1105 out_p.t2035 vp_p.t906 vdd.t2093 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1106 vdd.t2092 vp_p.t907 out_p.t2034 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1107 vdd.t2091 vp_p.t908 out_p.t2033 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1108 vdd.t2090 vp_p.t909 out_p.t2032 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1109 out_p.t2012 vp_p.t910 vdd.t2089 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1110 vdd.t2088 vp_p.t911 out_p.t2011 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1111 out_p.t2010 vp_p.t912 vdd.t2087 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1112 vdd.t2086 vp_p.t913 out_p.t2009 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1113 vdd.t2085 vp_p.t914 out_p.t1989 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1114 vdd.t2084 vp_p.t915 out_p.t1988 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1115 vdd.t2083 vp_p.t916 out_p.t1987 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1116 vdd.t2082 vp_p.t917 out_p.t1986 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1117 vdd.t2081 vp_p.t918 out_p.t1966 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1118 out_p.t1965 vp_p.t919 vdd.t2080 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1119 vdd.t2079 vp_p.t920 out_p.t1964 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1120 out_p.t1963 vp_p.t921 vdd.t2078 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1121 vdd.t2077 vp_p.t922 out_p.t1930 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1122 out_p.t1929 vp_p.t923 vdd.t2076 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1123 out_p.t1928 vp_p.t924 vdd.t2075 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1124 vdd.t2074 vp_p.t925 out_p.t1927 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1125 vdd.t2073 vp_p.t926 out_p.t1907 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1126 vdd.t2072 vp_p.t927 out_p.t1906 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1127 out_p.t1905 vp_p.t928 vdd.t2071 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1128 vdd.t2070 vp_p.t929 out_p.t1904 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1129 out_p.t1884 vp_p.t930 vdd.t2069 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1130 out_p.t1883 vp_p.t931 vdd.t2068 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1131 vdd.t2067 vp_p.t932 out_p.t1882 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1132 vdd.t2066 vp_p.t933 out_p.t1881 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1133 out_p.t1861 vp_p.t934 vdd.t2065 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1134 vdd.t2064 vp_p.t935 out_p.t1860 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1135 vdd.t2063 vp_p.t936 out_p.t1859 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1136 vdd.t2062 vp_p.t937 out_p.t1858 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1137 out_p.t1825 vp_p.t938 vdd.t2061 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1138 out_p.t1824 vp_p.t939 vdd.t2060 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1139 out_p.t1823 vp_p.t940 vdd.t2059 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1140 out_p.t1822 vp_p.t941 vdd.t2058 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1141 out_p.t1802 vp_p.t942 vdd.t2057 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1142 out_p.t1801 vp_p.t943 vdd.t2056 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1143 vdd.t2055 vp_p.t944 out_p.t1800 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1144 vdd.t2054 vp_p.t945 out_p.t1799 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1145 out_p.t1778 vp_p.t946 vdd.t2053 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1146 out_p.t1777 vp_p.t947 vdd.t2052 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1147 out_p.t1776 vp_p.t948 vdd.t2051 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1148 out_p.t1775 vp_p.t949 vdd.t2050 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1149 vdd.t2049 vp_p.t950 out_p.t1755 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1150 out_p.t1754 vp_p.t951 vdd.t2048 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1151 out_p.t1753 vp_p.t952 vdd.t2047 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1152 out_p.t1752 vp_p.t953 vdd.t2046 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1153 vdd.t2045 vp_p.t954 out_p.t1719 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1154 vdd.t2044 vp_p.t955 out_p.t1718 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1155 out_p.t1717 vp_p.t956 vdd.t2043 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1156 vdd.t2042 vp_p.t957 out_p.t1716 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1157 vdd.t2041 vp_p.t958 out_p.t1696 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1158 out_p.t1695 vp_p.t959 vdd.t2040 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1159 out_p.t1694 vp_p.t960 vdd.t2039 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1160 vdd.t2038 vp_p.t961 out_p.t1693 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1161 vdd.t2037 vp_p.t962 out_p.t1673 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1162 vdd.t2036 vp_p.t963 out_p.t1672 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1163 out_p.t1671 vp_p.t964 vdd.t2035 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1164 vdd.t2034 vp_p.t965 out_p.t1670 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1165 out_p.t1649 vp_p.t966 vdd.t2033 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1166 vdd.t2032 vp_p.t967 out_p.t1648 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1167 out_p.t1647 vp_p.t968 vdd.t2031 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1168 vdd.t2030 vp_p.t969 out_p.t1646 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1169 vdd.t2029 vp_p.t970 out_p.t1626 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1170 out_p.t163 vp_n.t199 vss.t400 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1171 out_p.t1625 vp_p.t971 vdd.t2028 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1172 vdd.t2027 vp_p.t972 out_p.t1624 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1173 vdd.t2026 vp_p.t973 out_p.t1623 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1174 out_p.t1607 vp_p.t974 vdd.t2025 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1175 out_p.t1606 vp_p.t975 vdd.t2024 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1176 out_p.t1605 vp_p.t976 vdd.t2023 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1177 out_p.t1604 vp_p.t977 vdd.t2022 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1178 vdd.t2021 vp_p.t978 out_p.t1584 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1179 out_p.t1583 vp_p.t979 vdd.t2020 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1180 vdd.t2019 vp_p.t980 out_p.t1582 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1181 vdd.t2018 vp_p.t981 out_p.t1581 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1182 out_p.t1561 vp_p.t982 vdd.t2017 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1183 out_p.t1560 vp_p.t983 vdd.t2016 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1184 out_p.t1559 vp_p.t984 vdd.t2015 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1185 vdd.t2014 vp_p.t985 out_p.t1558 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1186 out_p.t1538 vp_p.t986 vdd.t2013 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1187 out_p.t1537 vp_p.t987 vdd.t2012 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1188 vdd.t2011 vp_p.t988 out_p.t1536 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1189 out_p.t1535 vp_p.t989 vdd.t2010 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1190 vdd.t2009 vp_p.t990 out_p.t1501 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1191 vdd.t2008 vp_p.t991 out_p.t1500 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1192 vdd.t2007 vp_p.t992 out_p.t1499 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1193 vdd.t2006 vp_p.t993 out_p.t1498 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1194 out_p.t1484 vp_p.t994 vdd.t2005 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1195 out_p.t1483 vp_p.t995 vdd.t2004 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1196 vdd.t2003 vp_p.t996 out_p.t1482 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1197 vdd.t2002 vp_p.t997 out_p.t1481 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1198 vdd.t2001 vp_p.t998 out_p.t1460 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1199 out_p.t1459 vp_p.t999 vdd.t2000 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1200 out_p.t1458 vp_p.t1000 vdd.t1999 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1201 out_p.t1457 vp_p.t1001 vdd.t1998 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1202 vdd.t1997 vp_p.t1002 out_p.t1418 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1203 vdd.t1996 vp_p.t1003 out_p.t1417 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1204 vdd.t1995 vp_p.t1004 out_p.t1416 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1205 vdd.t1994 vp_p.t1005 out_p.t1415 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1206 vdd.t1993 vp_p.t1006 out_p.t1394 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1207 out_p.t1393 vp_p.t1007 vdd.t1992 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1208 out_p.t1392 vp_p.t1008 vdd.t1991 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1209 out_p.t1391 vp_p.t1009 vdd.t1990 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1210 vdd.t1989 vp_p.t1010 out_p.t1376 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1211 vdd.t1988 vp_p.t1011 out_p.t1375 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1212 vdd.t1987 vp_p.t1012 out_p.t1374 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1213 vdd.t1986 vp_p.t1013 out_p.t1373 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1214 vdd.t1985 vp_p.t1014 out_p.t2345 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1215 out_p.t2344 vp_p.t1015 vdd.t1984 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1216 vdd.t1983 vp_p.t1016 out_p.t2343 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1217 vdd.t1982 vp_p.t1017 out_p.t1615 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1218 vss.t399 vp_n.t200 out_p.t2 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1219 out_p.t1614 vp_p.t1018 vdd.t1981 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1220 out_p.t2256 vp_p.t1019 vdd.t1980 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1221 vdd.t1979 vp_p.t1020 out_p.t1218 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1222 vdd.t1978 vp_p.t1021 out_p.t1219 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1223 out_p.t1203 vp_p.t1022 vdd.t1977 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1224 out_p.t1205 vp_p.t1023 vdd.t1976 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1225 vdd.t1975 vp_p.t1024 out_p.t1207 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1226 out_p.t1202 vp_p.t1025 vdd.t1974 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1227 out_p.t1206 vp_p.t1026 vdd.t1973 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1228 vdd.t1972 vp_p.t1027 out_p.t1201 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1229 vdd.t1971 vp_p.t1028 out_p.t1200 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1230 vdd.t1970 vp_p.t1029 out_p.t1199 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1231 vdd.t1969 vp_p.t1030 out_p.t1198 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1232 out_p.t2463 vp_p.t1031 vdd.t1968 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1233 out_p.t2415 vp_p.t1032 vdd.t1967 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1234 vdd.t1966 vp_p.t1033 out_p.t2388 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1235 vdd.t1965 vp_p.t1034 out_p.t1229 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1236 out_p.t1224 vp_p.t1035 vdd.t1964 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1237 vdd.t1963 vp_p.t1036 out_p.t2369 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1238 vdd.t1962 vp_p.t1037 out_p.t2352 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1239 out_p.t2342 vp_p.t1038 vdd.t1961 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1240 out_p.t2325 vp_p.t1039 vdd.t1960 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1241 out_p.t2308 vp_p.t1040 vdd.t1959 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1242 out_p.t1223 vp_p.t1041 vdd.t1958 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1243 out_p.t0 vp_n.t201 vss.t398 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1244 out_p.t2291 vp_p.t1042 vdd.t1957 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1245 vss.t397 vp_n.t202 out_p.t3485 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1246 vdd.t1956 vp_p.t1043 out_p.t2269 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1247 out_p.t2255 vp_p.t1044 vdd.t1955 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1248 vdd.t1954 vp_p.t1045 out_p.t2232 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1249 vss.t396 vp_n.t203 out_p.t3483 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1250 vdd.t1953 vp_p.t1046 out_p.t2219 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1251 vdd.t1952 vp_p.t1047 out_p.t1221 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1252 out_p.t1220 vp_p.t1048 vdd.t1951 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1253 out_p.t2206 vp_p.t1049 vdd.t1950 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1254 vdd.t1949 vp_p.t1050 out_p.t2183 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1255 out_p.t2170 vp_p.t1051 vdd.t1948 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1256 out_p.t2147 vp_p.t1052 vdd.t1947 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1257 out_p.t2111 vp_p.t1053 vdd.t1946 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1258 vdd.t1945 vp_p.t1054 out_p.t2124 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1259 vdd.t1944 vp_p.t1055 out_p.t1217 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1260 out_p.t2100 vp_p.t1056 vdd.t1943 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1261 vss.t395 vp_n.t204 out_p.t367 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1262 vdd.t1942 vp_p.t1057 out_p.t2077 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1263 out_p.t1216 vp_p.t1058 vdd.t1941 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1264 vdd.t1940 vp_p.t1059 out_p.t2054 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1265 out_p.t2031 vp_p.t1060 vdd.t1939 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1266 vdd.t1938 vp_p.t1061 out_p.t2008 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1267 vdd.t1937 vp_p.t1062 out_p.t1215 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1268 vdd.t1936 vp_p.t1063 out_p.t1985 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1269 vdd.t1935 vp_p.t1064 out_p.t1962 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1270 vdd.t1934 vp_p.t1065 out_p.t1949 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1271 out_p.t1211 vp_p.t1066 vdd.t1933 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1272 out_p.t1926 vp_p.t1067 vdd.t1932 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1273 vdd.t1931 vp_p.t1068 out_p.t1214 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1274 vdd.t1930 vp_p.t1069 out_p.t1903 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1275 out_p.t1213 vp_p.t1070 vdd.t1929 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1276 out_p.t1880 vp_p.t1071 vdd.t1928 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1277 out_p.t1857 vp_p.t1072 vdd.t1927 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1278 out_p.t1844 vp_p.t1073 vdd.t1926 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1279 vdd.t1925 vp_p.t1074 out_p.t1212 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1280 vdd.t1924 vp_p.t1075 out_p.t1821 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1281 vdd.t1923 vp_p.t1076 out_p.t1785 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1282 vss.t394 vp_n.t205 out_p.t3545 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1283 out_p.t1798 vp_p.t1077 vdd.t1922 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1284 out_p.t1210 vp_p.t1078 vdd.t1921 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1285 out_p.t1774 vp_p.t1079 vdd.t1920 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1286 vdd.t1919 vp_p.t1080 out_p.t1751 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1287 out_p.t1738 vp_p.t1081 vdd.t1918 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1288 out_p.t1715 vp_p.t1082 vdd.t1917 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1289 vdd.t1916 vp_p.t1083 out_p.t1656 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1290 out_p.t1692 vp_p.t1084 vdd.t1915 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1291 out_p.t364 vp_n.t206 vss.t393 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1292 out_p.t1208 vp_p.t1085 vdd.t1914 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1293 vdd.t1913 vp_p.t1086 out_p.t1209 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1294 vdd.t1912 vp_p.t1087 out_p.t1669 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1295 out_p.t1645 vp_p.t1088 vdd.t1911 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1296 vdd.t1910 vp_p.t1089 out_p.t1622 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1297 out_p.t1603 vp_p.t1090 vdd.t1909 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1298 vdd.t1908 vp_p.t1091 out_p.t1580 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1299 vdd.t1907 vp_p.t1092 out_p.t1557 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1300 vdd.t1906 vp_p.t1093 out_p.t1508 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1301 out_p.t1204 vp_p.t1094 vdd.t1905 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1302 out_p.t1534 vp_p.t1095 vdd.t1904 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1303 vss.t392 vp_n.t207 out_p.t3543 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1304 out_p.t1521 vp_p.t1096 vdd.t1903 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1305 vdd.t1902 vp_p.t1097 out_p.t1467 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1306 out_p.t1425 vp_p.t1098 vdd.t1901 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1307 out_p.t1497 vp_p.t1099 vdd.t1900 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1308 out_p.t1197 vp_p.t1100 vdd.t1899 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1309 vdd.t1898 vp_p.t1101 out_p.t1191 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1310 vdd.t1897 vp_p.t1102 out_p.t1192 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1311 vss.t391 vp_n.t208 out_p.t361 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1312 out_p.t1193 vp_p.t1103 vdd.t1896 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1313 vdd.t1895 vp_p.t1104 out_p.t1194 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1314 out_p.t1195 vp_p.t1105 vdd.t1894 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1315 vdd.t1893 vp_p.t1106 out_p.t1196 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1316 out_p.t1401 vp_p.t1107 vdd.t1892 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1317 out_p.t1480 vp_p.t1108 vdd.t1891 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1318 out_p.t186 vp_n.t209 vss.t390 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1319 vdd.t1890 vp_p.t1109 out_p.t1383 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1320 vdd.t1889 vp_p.t1110 out_p.t1456 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1321 out_p.t1432 vp_p.t1111 vdd.t1888 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1322 vss.t389 vp_n.t210 out_p.t358 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1323 vdd.t1887 vp_p.t1112 out_p.t1414 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1324 vdd.t1886 vp_p.t1113 out_p.t1390 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1325 out_p.t1372 vp_p.t1114 vdd.t1885 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1326 vdd.t1884 vp_p.t1115 out_p.t454 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1327 out_p.t455 vp_p.t1116 vdd.t1883 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1328 out_p.t446 vp_p.t1117 vdd.t1882 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1329 out_p.t447 vp_p.t1118 vdd.t1881 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1330 out_p.t184 vp_n.t211 vss.t388 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1331 out_p.t448 vp_p.t1119 vdd.t1880 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1332 vdd.t1879 vp_p.t1120 out_p.t445 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1333 vdd.t1878 vp_p.t1121 out_p.t444 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1334 vdd.t1877 vp_p.t1122 out_p.t450 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1335 vdd.t1876 vp_p.t1123 out_p.t443 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1336 out_p.t428 vp_p.t1124 vdd.t1875 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1337 vdd.t1874 vp_p.t1125 out_p.t442 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1338 vdd.t1873 vp_p.t1126 out_p.t431 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1339 vss.t387 vp_n.t212 out_p.t379 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1340 vdd.t1872 vp_p.t1127 out_p.t441 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1341 vdd.t1871 vp_p.t1128 out_p.t435 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1342 vdd.t1870 vp_p.t1129 out_p.t440 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1343 vdd.t1869 vp_p.t1130 out_p.t437 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1344 out_p.t438 vp_p.t1131 vdd.t1868 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1345 vdd.t1867 vp_p.t1132 out_p.t436 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1346 out_p.t429 vp_p.t1133 vdd.t1866 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1347 out_p.t3534 vp_n.t213 vss.t386 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1348 out_p.t430 vp_p.t1134 vdd.t1865 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1349 out_p.t432 vp_p.t1135 vdd.t1864 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1350 vdd.t1863 vp_p.t1136 out_p.t433 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1351 vdd.t1862 vp_p.t1137 out_p.t434 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1352 vdd.t1861 vp_p.t1138 out_p.t3427 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1353 out_p.t3426 vp_p.t1139 vdd.t1860 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1354 out_p.t3425 vp_p.t1140 vdd.t1859 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1355 out_p.t3424 vp_p.t1141 vdd.t1858 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1356 out_p.t3423 vp_p.t1142 vdd.t1857 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1357 out_p.t376 vp_n.t214 vss.t385 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1358 vdd.t1856 vp_p.t1143 out_p.t3422 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1359 vdd.t1855 vp_p.t1144 out_p.t3421 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1360 vdd.t1854 vp_p.t1145 out_p.t3420 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1361 out_p.t3419 vp_p.t1146 vdd.t1853 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1362 out_p.t3418 vp_p.t1147 vdd.t1852 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1363 out_p.t3417 vp_p.t1148 vdd.t1851 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1364 vdd.t1850 vp_p.t1149 out_p.t3416 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1365 vdd.t1849 vp_p.t1150 out_p.t3415 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1366 vdd.t1848 vp_p.t1151 out_p.t3414 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1367 out_p.t3413 vp_p.t1152 vdd.t1847 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1368 vss.t384 vp_n.t215 out_p.t3531 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1369 out_p.t3412 vp_p.t1153 vdd.t1846 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1370 out_p.t3411 vp_p.t1154 vdd.t1845 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1371 vdd.t1844 vp_p.t1155 out_p.t3410 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1372 vdd.t1843 vp_p.t1156 out_p.t3409 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1373 out_p.t3408 vp_p.t1157 vdd.t1842 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1374 out_p.t3407 vp_p.t1158 vdd.t1841 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1375 vdd.t1840 vp_p.t1159 out_p.t3406 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1376 vdd.t1839 vp_p.t1160 out_p.t3405 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1377 vss.t383 vp_n.t216 out_p.t373 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1378 vss.t382 vp_n.t217 out_p.t3540 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1379 out_p.t3404 vp_p.t1161 vdd.t1838 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1380 out_p.t3403 vp_p.t1162 vdd.t1837 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1381 out_p.t3402 vp_p.t1163 vdd.t1836 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1382 vdd.t1835 vp_p.t1164 out_p.t3401 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1383 vdd.t1834 vp_p.t1165 out_p.t3400 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1384 out_p.t370 vp_n.t218 vss.t381 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1385 vdd.t1833 vp_p.t1166 out_p.t3399 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1386 vdd.t1832 vp_p.t1167 out_p.t3398 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1387 out_p.t3538 vp_n.t219 vss.t380 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1388 out_p.t391 vp_n.t220 vss.t379 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1389 vdd.t1831 vp_p.t1168 out_p.t3397 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1390 vdd.t1830 vp_p.t1169 out_p.t3396 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1391 out_p.t3395 vp_p.t1170 vdd.t1829 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1392 vdd.t1828 vp_p.t1171 out_p.t3394 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1393 out_p.t3393 vp_p.t1172 vdd.t1827 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1394 out_p.t3392 vp_p.t1173 vdd.t1826 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1395 out_p.t3391 vp_p.t1174 vdd.t1825 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1396 out_p.t3390 vp_p.t1175 vdd.t1824 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1397 vss.t378 vp_n.t221 out_p.t3549 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1398 out_p.t3389 vp_p.t1176 vdd.t1823 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1399 out_p.t3388 vp_p.t1177 vdd.t1822 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1400 vss.t377 vp_n.t222 out_p.t388 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1401 vdd.t1821 vp_p.t1178 out_p.t3387 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1402 out_p.t3386 vp_p.t1179 vdd.t1820 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1403 out_p.t3385 vp_p.t1180 vdd.t1819 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1404 out_p.t3384 vp_p.t1181 vdd.t1818 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1405 out_p.t3547 vp_n.t223 vss.t376 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1406 vdd.t1817 vp_p.t1182 out_p.t3383 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1407 vdd.t1816 vp_p.t1183 out_p.t3382 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1408 out_p.t385 vp_n.t224 vss.t375 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1409 out_p.t3381 vp_p.t1184 vdd.t1815 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1410 vdd.t1814 vp_p.t1185 out_p.t3380 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1411 vdd.t1813 vp_p.t1186 out_p.t3379 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1412 out_p.t3378 vp_p.t1187 vdd.t1812 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1413 vss.t374 vp_n.t225 out_p.t3555 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1414 vdd.t1811 vp_p.t1188 out_p.t3377 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1415 vdd.t1810 vp_p.t1189 out_p.t3376 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1416 out_p.t3375 vp_p.t1190 vdd.t1809 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1417 vdd.t1808 vp_p.t1191 out_p.t3374 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1418 vdd.t1807 vp_p.t1192 out_p.t3373 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1419 out_p.t3372 vp_p.t1193 vdd.t1806 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1420 vdd.t1805 vp_p.t1194 out_p.t3371 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1421 out_p.t3370 vp_p.t1195 vdd.t1804 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1422 vdd.t1803 vp_p.t1196 out_p.t3369 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1423 out_p.t3368 vp_p.t1197 vdd.t1802 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1424 out_p.t3367 vp_p.t1198 vdd.t1801 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1425 out_p.t3366 vp_p.t1199 vdd.t1800 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1426 vss.t373 vp_n.t226 out_p.t382 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1427 vss.t372 vp_n.t227 out_p.t3553 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1428 vdd.t1799 vp_p.t1200 out_p.t3365 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1429 out_p.t3364 vp_p.t1201 vdd.t1798 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1430 vss.t371 vp_n.t228 out_p.t403 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1431 vdd.t1797 vp_p.t1202 out_p.t3363 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1432 vdd.t1796 vp_p.t1203 out_p.t3362 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1433 out_p.t3361 vp_p.t1204 vdd.t1795 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1434 vdd.t1794 vp_p.t1205 out_p.t3360 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1435 vdd.t1793 vp_p.t1206 out_p.t3359 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1436 out_p.t3358 vp_p.t1207 vdd.t1792 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1437 vdd.t1791 vp_p.t1208 out_p.t3357 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1438 out_p.t3356 vp_p.t1209 vdd.t1790 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1439 out_p.t3473 vp_n.t229 vss.t370 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1440 out_p.t3355 vp_p.t1210 vdd.t1789 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1441 vdd.t1788 vp_p.t1211 out_p.t3354 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1442 out_p.t3353 vp_p.t1212 vdd.t1787 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1443 out_p.t3352 vp_p.t1213 vdd.t1786 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1444 out_p.t3351 vp_p.t1214 vdd.t1785 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1445 out_p.t400 vp_n.t230 vss.t369 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1446 vss.t368 vp_n.t231 out_p.t3457 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1447 out_p.t3350 vp_p.t1215 vdd.t1784 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1448 vss.t367 vp_n.t232 out_p.t397 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1449 out_p.t420 vp_n.t233 vss.t366 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1450 out_p.t3349 vp_p.t1216 vdd.t1783 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1451 vdd.t1782 vp_p.t1217 out_p.t3348 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1452 vdd.t1781 vp_p.t1218 out_p.t3347 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1453 vss.t365 vp_n.t234 out_p.t394 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1454 vss.t364 vp_n.t235 out_p.t418 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1455 out_p.t3346 vp_p.t1219 vdd.t1780 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1456 out_p.t3345 vp_p.t1220 vdd.t1779 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1457 out_p.t3344 vp_p.t1221 vdd.t1778 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1458 vdd.t1777 vp_p.t1222 out_p.t3343 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1459 vdd.t1776 vp_p.t1223 out_p.t3342 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1460 out_p.t407 vp_n.t236 vss.t363 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1461 vdd.t1775 vp_p.t1224 out_p.t3341 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1462 out_p.t3340 vp_p.t1225 vdd.t1774 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1463 out_p.t3496 vp_n.t237 vss.t362 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1464 out_p.t3339 vp_p.t1226 vdd.t1773 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1465 vss.t361 vp_n.t238 out_p.t346 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1466 vdd.t1772 vp_p.t1227 out_p.t3338 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1467 out_p.t3337 vp_p.t1228 vdd.t1771 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1468 vss.t360 vp_n.t239 out_p.t406 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1469 out_p.t3336 vp_p.t1229 vdd.t1770 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1470 vdd.t1769 vp_p.t1230 out_p.t3335 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1471 out_p.t68 vp_n.t240 vss.t359 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1472 vss.t358 vp_n.t241 out_p.t349 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1473 out_p.t3334 vp_p.t1231 vdd.t1768 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1474 out_p.t3333 vp_p.t1232 vdd.t1767 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1475 out_p.t3332 vp_p.t1233 vdd.t1766 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1476 vss.t357 vp_n.t242 out_p.t3475 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1477 out_p.t405 vp_n.t243 vss.t356 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1478 out_p.t3462 vp_n.t244 vss.t355 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1479 vss.t354 vp_n.t245 out_p.t266 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1480 vdd.t1765 vp_p.t1234 out_p.t3331 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1481 out_p.t3330 vp_p.t1235 vdd.t1764 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1482 vss.t353 vp_n.t246 out_p.t409 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1483 vdd.t1763 vp_p.t1236 out_p.t3329 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1484 vdd.t1762 vp_p.t1237 out_p.t3328 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1485 out_p.t3327 vp_p.t1238 vdd.t1761 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1486 out_p.t3326 vp_p.t1239 vdd.t1760 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1487 out_p.t3325 vp_p.t1240 vdd.t1759 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1488 out_p.t262 vp_n.t247 vss.t352 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1489 vdd.t1758 vp_p.t1241 out_p.t3324 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1490 out_p.t246 vp_n.t248 vss.t351 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1491 vdd.t1757 vp_p.t1242 out_p.t3323 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1492 vdd.t1756 vp_p.t1243 out_p.t3322 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1493 out_p.t3321 vp_p.t1244 vdd.t1755 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1494 out_p.t3320 vp_p.t1245 vdd.t1754 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1495 out_p.t3319 vp_p.t1246 vdd.t1753 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1496 vdd.t1752 vp_p.t1247 out_p.t3318 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1497 vdd.t1751 vp_p.t1248 out_p.t3317 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1498 vss.t350 vp_n.t249 out_p.t3571 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1499 vdd.t1750 vp_p.t1249 out_p.t3316 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1500 vss.t349 vp_n.t250 out_p.t408 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1501 out_p.t3315 vp_p.t1250 vdd.t1749 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1502 out_p.t3314 vp_p.t1251 vdd.t1748 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1503 out_p.t3313 vp_p.t1252 vdd.t1747 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1504 out_p.t3312 vp_p.t1253 vdd.t1746 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1505 out_p.t3311 vp_p.t1254 vdd.t1745 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1506 vss.t348 vp_n.t251 out_p.t3569 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1507 vdd.t1744 vp_p.t1255 out_p.t3310 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1508 out_p.t3309 vp_p.t1256 vdd.t1743 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1509 vss.t347 vp_n.t252 out_p.t174 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1510 out_p.t413 vp_n.t253 vss.t346 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1511 vss.t345 vp_n.t254 out_p.t3598 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1512 out_p.t3308 vp_p.t1257 vdd.t1742 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1513 vdd.t1741 vp_p.t1258 out_p.t3307 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1514 vdd.t1740 vp_p.t1259 out_p.t3306 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1515 vdd.t1739 vp_p.t1260 out_p.t3305 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1516 out_p.t3304 vp_p.t1261 vdd.t1738 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1517 vdd.t1737 vp_p.t1262 out_p.t3303 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1518 out_p.t412 vp_n.t255 vss.t344 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1519 vdd.t1736 vp_p.t1263 out_p.t3302 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1520 vdd.t1735 vp_p.t1264 out_p.t3301 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1521 out_p.t3596 vp_n.t256 vss.t343 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1522 out_p.t3300 vp_p.t1265 vdd.t1734 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1523 out_p.t3299 vp_p.t1266 vdd.t1733 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1524 out_p.t411 vp_n.t257 vss.t342 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1525 vdd.t1732 vp_p.t1267 out_p.t3298 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1526 out_p.t3297 vp_p.t1268 vdd.t1731 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1527 vdd.t1730 vp_p.t1269 out_p.t3296 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1528 vdd.t1729 vp_p.t1270 out_p.t3295 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1529 out_p.t3464 vp_n.t258 vss.t341 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1530 vss.t340 vp_n.t259 out_p.t410 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1531 vdd.t1728 vp_p.t1271 out_p.t3294 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1532 out_p.t3293 vp_p.t1272 vdd.t1727 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1533 vdd.t1726 vp_p.t1273 out_p.t3292 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1534 vss.t339 vp_n.t260 out_p.t181 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1535 vdd.t1725 vp_p.t1274 out_p.t3291 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1536 out_p.t3290 vp_p.t1275 vdd.t1724 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1537 vss.t338 vp_n.t261 out_p.t417 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1538 out_p.t3289 vp_p.t1276 vdd.t1723 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1539 out_p.t3288 vp_p.t1277 vdd.t1722 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1540 vdd.t1721 vp_p.t1278 out_p.t3287 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1541 out_p.t347 vp_n.t262 vss.t337 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1542 vdd.t1720 vp_p.t1279 out_p.t3286 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1543 out_p.t3285 vp_p.t1280 vdd.t1719 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1544 vss.t336 vp_n.t263 out_p.t179 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1545 vss.t335 vp_n.t264 out_p.t416 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1546 vdd.t1718 vp_p.t1281 out_p.t3284 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1547 out_p.t3283 vp_p.t1282 vdd.t1717 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1548 out_p.t3282 vp_p.t1283 vdd.t1716 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1549 out_p.t3281 vp_p.t1284 vdd.t1715 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1550 vdd.t1714 vp_p.t1285 out_p.t3280 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1551 vdd.t1713 vp_p.t1286 out_p.t3279 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1552 vss.t334 vp_n.t265 out_p.t415 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1553 out_p.t3278 vp_p.t1287 vdd.t1712 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1554 vss.t333 vp_n.t266 out_p.t176 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1555 out_p.t414 vp_n.t267 vss.t332 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1556 vdd.t1711 vp_p.t1288 out_p.t3277 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1557 vdd.t1710 vp_p.t1289 out_p.t3276 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1558 vss.t331 vp_n.t268 out_p.t3453 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1559 out_p.t3517 vp_n.t269 vss.t330 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1560 vdd.t1709 vp_p.t1290 out_p.t3275 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1561 out_p.t3589 vp_n.t270 vss.t329 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1562 out_p.t3274 vp_p.t1291 vdd.t1708 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1563 out_p.t336 vp_n.t271 vss.t328 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1564 vdd.t1707 vp_p.t1292 out_p.t3273 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1565 vdd.t1706 vp_p.t1293 out_p.t3272 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1566 out_p.t329 vp_n.t272 vss.t327 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1567 vdd.t1705 vp_p.t1294 out_p.t3271 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1568 out_p.t335 vp_n.t273 vss.t326 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1569 vdd.t1704 vp_p.t1295 out_p.t3270 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1570 vdd.t1703 vp_p.t1296 out_p.t3269 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1571 vss.t325 vp_n.t274 out_p.t343 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1572 vdd.t1702 vp_p.t1297 out_p.t3268 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1573 vss.t324 vp_n.t275 out_p.t338 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1574 out_p.t3267 vp_p.t1298 vdd.t1701 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1575 out_p.t3266 vp_p.t1299 vdd.t1700 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1576 out_p.t3514 vp_n.t276 vss.t323 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1577 vdd.t1699 vp_p.t1300 out_p.t3265 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1578 out_p.t3264 vp_p.t1301 vdd.t1698 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1579 vss.t322 vp_n.t277 out_p.t3519 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1580 vss.t321 vp_n.t278 out_p.t3504 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1581 vdd.t1697 vp_p.t1302 out_p.t3263 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1582 vdd.t1696 vp_p.t1303 out_p.t3262 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1583 vdd.t1695 vp_p.t1304 out_p.t3261 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1584 vdd.t1694 vp_p.t1305 out_p.t3260 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1585 vdd.t1693 vp_p.t1306 out_p.t3259 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1586 vss.t320 vp_n.t279 out_p.t3498 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1587 vdd.t1692 vp_p.t1307 out_p.t3258 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1588 vdd.t1691 vp_p.t1308 out_p.t3257 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1589 out_p.t3256 vp_p.t1309 vdd.t1690 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1590 out_p.t3512 vp_n.t280 vss.t319 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1591 vdd.t1689 vp_p.t1310 out_p.t3255 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1592 vdd.t1688 vp_p.t1311 out_p.t3254 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1593 vdd.t1687 vp_p.t1312 out_p.t3253 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1594 vss.t318 vp_n.t281 out_p.t3520 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1595 vdd.t1686 vp_p.t1313 out_p.t3252 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1596 vdd.t1685 vp_p.t1314 out_p.t3251 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1597 out_p.t3250 vp_p.t1315 vdd.t1684 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1598 out_p.t3249 vp_p.t1316 vdd.t1683 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1599 out_p.t3248 vp_p.t1317 vdd.t1682 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1600 vdd.t1681 vp_p.t1318 out_p.t3247 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1601 vdd.t1680 vp_p.t1319 out_p.t3246 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1602 out_p.t188 vp_n.t282 vss.t317 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1603 vss.t316 vp_n.t283 out_p.t404 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1604 out_p.t3566 vp_n.t284 vss.t315 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1605 out_p.t3245 vp_p.t1320 vdd.t1679 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1606 out_p.t3244 vp_p.t1321 vdd.t1678 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1607 vdd.t1677 vp_p.t1322 out_p.t3243 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1608 out_p.t3242 vp_p.t1323 vdd.t1676 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1609 vdd.t1675 vp_p.t1324 out_p.t3241 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1610 vdd.t1674 vp_p.t1325 out_p.t3240 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1611 out_p.t3239 vp_p.t1326 vdd.t1673 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1612 vdd.t1672 vp_p.t1327 out_p.t3238 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1613 vdd.t1671 vp_p.t1328 out_p.t3237 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1614 out_p.t3236 vp_p.t1329 vdd.t1670 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1615 out_p.t402 vp_n.t285 vss.t314 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1616 out_p.t3235 vp_p.t1330 vdd.t1669 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1617 vdd.t1668 vp_p.t1331 out_p.t3234 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1618 out_p.t3233 vp_p.t1332 vdd.t1667 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1619 vss.t313 vp_n.t286 out_p.t3565 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1620 vss.t312 vp_n.t287 out_p.t5 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1621 vdd.t1666 vp_p.t1333 out_p.t3232 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1622 out_p.t3231 vp_p.t1334 vdd.t1665 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1623 out_p.t3230 vp_p.t1335 vdd.t1664 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1624 vdd.t1663 vp_p.t1336 out_p.t3229 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1625 vdd.t1662 vp_p.t1337 out_p.t3228 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1626 out_p.t3227 vp_p.t1338 vdd.t1661 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1627 vdd.t1660 vp_p.t1339 out_p.t3226 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1628 vss.t311 vp_n.t288 out_p.t401 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1629 vdd.t1659 vp_p.t1340 out_p.t3225 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1630 out_p.t224 vp_n.t289 vss.t310 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1631 vdd.t1658 vp_p.t1341 out_p.t3224 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1632 vss.t309 vp_n.t290 out_p.t3590 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1633 out_p.t308 vp_n.t291 vss.t308 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1634 out_p.t3223 vp_p.t1342 vdd.t1657 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1635 vdd.t1656 vp_p.t1343 out_p.t3222 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1636 vdd.t1655 vp_p.t1344 out_p.t3221 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1637 vdd.t1654 vp_p.t1345 out_p.t3220 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1638 out_p.t3219 vp_p.t1346 vdd.t1653 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1639 vdd.t1652 vp_p.t1347 out_p.t3218 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1640 vss.t307 vp_n.t292 out_p.t309 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1641 out_p.t399 vp_n.t293 vss.t306 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1642 vdd.t1651 vp_p.t1348 out_p.t3217 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1643 vdd.t1650 vp_p.t1349 out_p.t3216 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1644 out_p.t6 vp_n.t294 vss.t305 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1645 out_p.t3215 vp_p.t1350 vdd.t1649 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1646 vdd.t1648 vp_p.t1351 out_p.t3214 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1647 vdd.t1647 vp_p.t1352 out_p.t3213 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1648 vdd.t1646 vp_p.t1353 out_p.t3212 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1649 out_p.t172 vp_n.t295 vss.t304 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1650 vss.t303 vp_n.t296 out_p.t398 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1651 out_p.t3211 vp_p.t1354 vdd.t1645 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1652 vdd.t1644 vp_p.t1355 out_p.t3210 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1653 vss.t302 vp_n.t297 out_p.t3588 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1654 out_p.t306 vp_n.t298 vss.t301 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1655 out_p.t3209 vp_p.t1356 vdd.t1643 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1656 vdd.t1642 vp_p.t1357 out_p.t3208 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1657 out_p.t307 vp_n.t299 vss.t300 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1658 vss.t299 vp_n.t300 out_p.t396 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1659 out_p.t3207 vp_p.t1358 vdd.t1641 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1660 out_p.t3206 vp_p.t1359 vdd.t1640 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1661 out_p.t173 vp_n.t301 vss.t298 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1662 vss.t297 vp_n.t302 out_p.t169 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1663 vdd.t1639 vp_p.t1360 out_p.t3205 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1664 vdd.t1638 vp_p.t1361 out_p.t3204 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1665 vdd.t1637 vp_p.t1362 out_p.t3203 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1666 out_p.t395 vp_n.t303 vss.t296 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1667 vdd.t1636 vp_p.t1363 out_p.t3202 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1668 vdd.t1635 vp_p.t1364 out_p.t3201 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1669 vss.t295 vp_n.t304 out_p.t223 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1670 vdd.t1634 vp_p.t1365 out_p.t3200 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1671 out_p.t3199 vp_p.t1366 vdd.t1633 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1672 vdd.t1632 vp_p.t1367 out_p.t3198 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1673 out_p.t3582 vp_n.t305 vss.t294 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1674 out_p.t303 vp_n.t306 vss.t293 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1675 vdd.t1631 vp_p.t1368 out_p.t3197 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1676 out_p.t3196 vp_p.t1369 vdd.t1630 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1677 vdd.t1629 vp_p.t1370 out_p.t3195 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1678 vss.t292 vp_n.t307 out_p.t304 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1679 out_p.t3194 vp_p.t1371 vdd.t1628 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1680 vdd.t1627 vp_p.t1372 out_p.t3193 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1681 out_p.t3192 vp_p.t1373 vdd.t1626 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1682 vdd.t1625 vp_p.t1374 out_p.t3191 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1683 out_p.t3190 vp_p.t1375 vdd.t1624 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1684 out_p.t3189 vp_p.t1376 vdd.t1623 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1685 vdd.t1622 vp_p.t1377 out_p.t3188 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1686 out_p.t3187 vp_p.t1378 vdd.t1621 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1687 out_p.t3186 vp_p.t1379 vdd.t1620 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1688 out_p.t3185 vp_p.t1380 vdd.t1619 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1689 vdd.t1618 vp_p.t1381 out_p.t3184 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1690 out_p.t3183 vp_p.t1382 vdd.t1617 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1691 vdd.t1616 vp_p.t1383 out_p.t3182 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1692 out_p.t3181 vp_p.t1384 vdd.t1615 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1693 out_p.t393 vp_n.t308 vss.t291 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1694 out_p.t3180 vp_p.t1385 vdd.t1614 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1695 out_p.t170 vp_n.t309 vss.t290 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1696 out_p.t3179 vp_p.t1386 vdd.t1613 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1697 vdd.t1612 vp_p.t1387 out_p.t3178 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1698 vdd.t1611 vp_p.t1388 out_p.t3177 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1699 vss.t289 vp_n.t310 out_p.t167 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1700 vdd.t1610 vp_p.t1389 out_p.t3176 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1701 out_p.t3175 vp_p.t1390 vdd.t1609 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1702 out_p.t3174 vp_p.t1391 vdd.t1608 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1703 out_p.t3173 vp_p.t1392 vdd.t1607 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1704 vdd.t1606 vp_p.t1393 out_p.t3172 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1705 vdd.t1605 vp_p.t1394 out_p.t3171 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1706 out_p.t392 vp_n.t311 vss.t288 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1707 vss.t287 vp_n.t312 out_p.t3581 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1708 out_p.t3170 vp_p.t1395 vdd.t1604 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1709 vdd.t1603 vp_p.t1396 out_p.t3169 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1710 out_p.t3168 vp_p.t1397 vdd.t1602 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1711 out_p.t3167 vp_p.t1398 vdd.t1601 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1712 vdd.t1600 vp_p.t1399 out_p.t3166 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1713 out_p.t301 vp_n.t313 vss.t286 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1714 out_p.t3165 vp_p.t1400 vdd.t1599 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1715 vdd.t1598 vp_p.t1401 out_p.t3164 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1716 vss.t285 vp_n.t314 out_p.t302 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1717 out_p.t3163 vp_p.t1402 vdd.t1597 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1718 out_p.t390 vp_n.t315 vss.t284 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1719 vss.t283 vp_n.t316 out_p.t168 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1720 vdd.t1596 vp_p.t1403 out_p.t3162 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1721 out_p.t161 vp_n.t317 vss.t282 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1722 out_p.t389 vp_n.t318 vss.t281 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1723 out_p.t222 vp_n.t319 vss.t280 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1724 vdd.t1595 vp_p.t1404 out_p.t3161 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1725 vdd.t1594 vp_p.t1405 out_p.t3160 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1726 out_p.t3580 vp_n.t320 vss.t279 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1727 vss.t278 vp_n.t321 out_p.t299 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1728 vdd.t1593 vp_p.t1406 out_p.t3159 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1729 out_p.t3158 vp_p.t1407 vdd.t1592 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1730 vdd.t1591 vp_p.t1408 out_p.t3157 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1731 vss.t277 vp_n.t322 out_p.t300 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1732 out_p.t387 vp_n.t323 vss.t276 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1733 out_p.t3156 vp_p.t1409 vdd.t1590 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1734 vdd.t1589 vp_p.t1410 out_p.t3155 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1735 out_p.t3154 vp_p.t1411 vdd.t1588 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1736 vss.t275 vp_n.t324 out_p.t162 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1737 out_p.t3153 vp_p.t1412 vdd.t1587 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1738 out_p.t160 vp_n.t325 vss.t274 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1739 out_p.t3152 vp_p.t1413 vdd.t1586 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1740 vss.t273 vp_n.t326 out_p.t386 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1741 out_p.t221 vp_n.t327 vss.t272 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1742 out_p.t3151 vp_p.t1414 vdd.t1585 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1743 out_p.t3150 vp_p.t1415 vdd.t1584 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1744 vdd.t1583 vp_p.t1416 out_p.t3149 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1745 vss.t271 vp_n.t328 out_p.t3447 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1746 vdd.t1582 vp_p.t1417 out_p.t3148 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1747 vdd.t1581 vp_p.t1418 out_p.t3147 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1748 vdd.t1580 vp_p.t1419 out_p.t3146 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1749 out_p.t296 vp_n.t329 vss.t270 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1750 out_p.t297 vp_n.t330 vss.t269 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1751 out_p.t3145 vp_p.t1420 vdd.t1579 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1752 out_p.t3144 vp_p.t1421 vdd.t1578 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1753 vdd.t1577 vp_p.t1422 out_p.t3143 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1754 vdd.t1576 vp_p.t1423 out_p.t3142 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1755 vdd.t1575 vp_p.t1424 out_p.t3141 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1756 vdd.t1574 vp_p.t1425 out_p.t3140 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1757 out_p.t384 vp_n.t331 vss.t268 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1758 vdd.t1573 vp_p.t1426 out_p.t3139 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1759 vss.t267 vp_n.t332 out_p.t159 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1760 vdd.t1572 vp_p.t1427 out_p.t3138 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1761 out_p.t3137 vp_p.t1428 vdd.t1571 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1762 vss.t266 vp_n.t333 out_p.t383 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1763 out_p.t3136 vp_p.t1429 vdd.t1570 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1764 vss.t265 vp_n.t334 out_p.t220 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1765 vdd.t1569 vp_p.t1430 out_p.t3135 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1766 vdd.t1568 vp_p.t1431 out_p.t3134 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1767 out_p.t3133 vp_p.t1432 vdd.t1567 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1768 out_p.t3132 vp_p.t1433 vdd.t1566 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1769 out_p.t3446 vp_n.t335 vss.t264 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1770 vdd.t1565 vp_p.t1434 out_p.t3131 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1771 vss.t263 vp_n.t336 out_p.t295 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1772 out_p.t3130 vp_p.t1435 vdd.t1564 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1773 out_p.t3129 vp_p.t1436 vdd.t1563 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1774 vdd.t1562 vp_p.t1437 out_p.t3128 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1775 vdd.t1561 vp_p.t1438 out_p.t3127 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1776 out_p.t3126 vp_p.t1439 vdd.t1560 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1777 out_p.t3125 vp_p.t1440 vdd.t1559 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1778 vss.t262 vp_n.t337 out_p.t381 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1779 out_p.t3124 vp_p.t1441 vdd.t1558 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1780 out_p.t3123 vp_p.t1442 vdd.t1557 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1781 vdd.t1556 vp_p.t1443 out_p.t3122 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1782 out_p.t3121 vp_p.t1444 vdd.t1555 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1783 out_p.t33 vp_n.t338 vss.t261 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1784 vdd.t1554 vp_p.t1445 out_p.t3120 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1785 vdd.t1553 vp_p.t1446 out_p.t3119 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1786 out_p.t3118 vp_p.t1447 vdd.t1552 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1787 vdd.t1551 vp_p.t1448 out_p.t3117 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1788 out_p.t34 vp_n.t339 vss.t260 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1789 out_p.t293 vp_n.t340 vss.t259 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1790 out_p.t3116 vp_p.t1449 vdd.t1550 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1791 vdd.t1549 vp_p.t1450 out_p.t3115 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1792 out_p.t3114 vp_p.t1451 vdd.t1548 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1793 out_p.t3113 vp_p.t1452 vdd.t1547 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1794 vdd.t1546 vp_p.t1453 out_p.t3112 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1795 vdd.t1545 vp_p.t1454 out_p.t3111 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1796 vss.t258 vp_n.t341 out_p.t380 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1797 vdd.t1544 vp_p.t1455 out_p.t3110 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1798 out_p.t3109 vp_p.t1456 vdd.t1543 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1799 vdd.t1542 vp_p.t1457 out_p.t3108 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1800 out_p.t3107 vp_p.t1458 vdd.t1541 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1801 out_p.t3106 vp_p.t1459 vdd.t1540 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1802 out_p.t3105 vp_p.t1460 vdd.t1539 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1803 vss.t257 vp_n.t342 out_p.t3478 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1804 out_p.t292 vp_n.t343 vss.t256 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1805 vss.t255 vp_n.t344 out_p.t378 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1806 vdd.t1538 vp_p.t1461 out_p.t3104 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1807 out_p.t35 vp_n.t345 vss.t254 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1808 out_p.t3103 vp_p.t1462 vdd.t1537 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1809 out_p.t3102 vp_p.t1463 vdd.t1536 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1810 vdd.t1535 vp_p.t1464 out_p.t3101 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1811 vdd.t1534 vp_p.t1465 out_p.t3100 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1812 out_p.t3099 vp_p.t1466 vdd.t1533 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1813 vdd.t1532 vp_p.t1467 out_p.t3098 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1814 vss.t253 vp_n.t346 out_p.t37 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1815 out_p.t3097 vp_p.t1468 vdd.t1531 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1816 vdd.t1530 vp_p.t1469 out_p.t3096 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1817 vss.t252 vp_n.t347 out_p.t377 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1818 out_p.t3095 vp_p.t1470 vdd.t1529 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1819 out_p.t219 vp_n.t348 vss.t251 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1820 out_p.t3094 vp_p.t1471 vdd.t1528 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1821 vdd.t1527 vp_p.t1472 out_p.t3093 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1822 vdd.t1526 vp_p.t1473 out_p.t3092 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1823 vdd.t1525 vp_p.t1474 out_p.t3091 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1824 out_p.t3477 vp_n.t349 vss.t250 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1825 vdd.t1524 vp_p.t1475 out_p.t3090 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1826 vdd.t1523 vp_p.t1476 out_p.t3089 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1827 vdd.t1522 vp_p.t1477 out_p.t3088 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1828 out_p.t3087 vp_p.t1478 vdd.t1521 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1829 out_p.t3086 vp_p.t1479 vdd.t1520 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1830 vss.t249 vp_n.t350 out_p.t291 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1831 vdd.t1519 vp_p.t1480 out_p.t3085 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1832 vdd.t1518 vp_p.t1481 out_p.t3084 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1833 vss.t248 vp_n.t351 out_p.t375 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1834 vdd.t1517 vp_p.t1482 out_p.t3083 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1835 out_p.t3082 vp_p.t1483 vdd.t1516 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1836 vdd.t1515 vp_p.t1484 out_p.t3081 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1837 vdd.t1514 vp_p.t1485 out_p.t3080 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1838 out_p.t38 vp_n.t352 vss.t247 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1839 vdd.t1513 vp_p.t1486 out_p.t3079 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1840 out_p.t3078 vp_p.t1487 vdd.t1512 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1841 out_p.t3077 vp_p.t1488 vdd.t1511 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1842 out_p.t3076 vp_p.t1489 vdd.t1510 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1843 vdd.t1509 vp_p.t1490 out_p.t3075 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1844 vdd.t1508 vp_p.t1491 out_p.t3074 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1845 vdd.t1507 vp_p.t1492 out_p.t3073 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1846 vdd.t1506 vp_p.t1493 out_p.t3072 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1847 out_p.t3071 vp_p.t1494 vdd.t1505 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1848 out_p.t3070 vp_p.t1495 vdd.t1504 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1849 out_p.t3069 vp_p.t1496 vdd.t1503 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1850 out_p.t3068 vp_p.t1497 vdd.t1502 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1851 out_p.t40 vp_n.t353 vss.t246 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1852 vdd.t1501 vp_p.t1498 out_p.t3067 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1853 out_p.t374 vp_n.t354 vss.t245 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1854 vdd.t1500 vp_p.t1499 out_p.t3066 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1855 out_p.t3065 vp_p.t1500 vdd.t1499 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1856 out_p.t3064 vp_p.t1501 vdd.t1498 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1857 out_p.t3063 vp_p.t1502 vdd.t1497 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1858 vdd.t1496 vp_p.t1503 out_p.t3062 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1859 out_p.t3061 vp_p.t1504 vdd.t1495 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1860 out_p.t3060 vp_p.t1505 vdd.t1494 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1861 vss.t244 vp_n.t355 out_p.t3439 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1862 vdd.t1493 vp_p.t1506 out_p.t3059 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1863 vdd.t1492 vp_p.t1507 out_p.t3058 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1864 out_p.t289 vp_n.t356 vss.t243 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1865 out_p.t3057 vp_p.t1508 vdd.t1491 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1866 out_p.t3056 vp_p.t1509 vdd.t1490 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1867 out_p.t3055 vp_p.t1510 vdd.t1489 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1868 vdd.t1488 vp_p.t1511 out_p.t3054 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1869 vdd.t1487 vp_p.t1512 out_p.t3053 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1870 out_p.t3052 vp_p.t1513 vdd.t1486 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1871 vdd.t1485 vp_p.t1514 out_p.t3051 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1872 out_p.t3050 vp_p.t1515 vdd.t1484 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1873 vdd.t1483 vp_p.t1516 out_p.t3049 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1874 vss.t242 vp_n.t357 out_p.t372 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1875 out_p.t41 vp_n.t358 vss.t241 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1876 vdd.t1482 vp_p.t1517 out_p.t3048 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1877 out_p.t3047 vp_p.t1518 vdd.t1481 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1878 out_p.t3046 vp_p.t1519 vdd.t1480 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1879 vss.t240 vp_n.t359 out_p.t43 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1880 out_p.t371 vp_n.t360 vss.t239 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1881 vdd.t1479 vp_p.t1520 out_p.t3045 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1882 vdd.t1478 vp_p.t1521 out_p.t3044 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1883 out_p.t218 vp_n.t361 vss.t238 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1884 out_p.t3043 vp_p.t1522 vdd.t1477 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1885 vdd.t1476 vp_p.t1523 out_p.t3042 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1886 out_p.t3041 vp_p.t1524 vdd.t1475 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1887 out_p.t3040 vp_p.t1525 vdd.t1474 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1888 out_p.t3039 vp_p.t1526 vdd.t1473 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1889 vdd.t1472 vp_p.t1527 out_p.t3038 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1890 vdd.t1471 vp_p.t1528 out_p.t3037 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1891 vdd.t1470 vp_p.t1529 out_p.t3036 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1892 out_p.t3035 vp_p.t1530 vdd.t1469 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1893 vdd.t1468 vp_p.t1531 out_p.t3034 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1894 vss.t237 vp_n.t362 out_p.t3438 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1895 out_p.t3033 vp_p.t1532 vdd.t1467 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1896 out_p.t3032 vp_p.t1533 vdd.t1466 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1897 out_p.t3031 vp_p.t1534 vdd.t1465 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1898 out_p.t286 vp_n.t363 vss.t236 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1899 vss.t235 vp_n.t364 out_p.t287 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1900 out_p.t3030 vp_p.t1535 vdd.t1464 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1901 out_p.t3029 vp_p.t1536 vdd.t1463 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1902 vdd.t1462 vp_p.t1537 out_p.t3028 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1903 out_p.t369 vp_n.t365 vss.t234 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1904 out_p.t3027 vp_p.t1538 vdd.t1461 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1905 out_p.t3026 vp_p.t1539 vdd.t1460 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1906 vdd.t1459 vp_p.t1540 out_p.t3025 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1907 out_p.t44 vp_n.t366 vss.t233 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1908 out_p.t3024 vp_p.t1541 vdd.t1458 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1909 vdd.t1457 vp_p.t1542 out_p.t3023 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1910 out_p.t3022 vp_p.t1543 vdd.t1456 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1911 vdd.t1455 vp_p.t1544 out_p.t3021 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1912 out_p.t3020 vp_p.t1545 vdd.t1454 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1913 out_p.t46 vp_n.t367 vss.t232 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1914 vss.t231 vp_n.t368 out_p.t368 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1915 vdd.t1453 vp_p.t1546 out_p.t3019 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1916 out_p.t3018 vp_p.t1547 vdd.t1452 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1917 out_p.t3017 vp_p.t1548 vdd.t1451 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1918 out_p.t3016 vp_p.t1549 vdd.t1450 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1919 vdd.t1449 vp_p.t1550 out_p.t3015 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1920 vss.t230 vp_n.t369 out_p.t217 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1921 out_p.t3014 vp_p.t1551 vdd.t1448 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1922 vdd.t1447 vp_p.t1552 out_p.t3013 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1923 vdd.t1446 vp_p.t1553 out_p.t3012 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1924 out_p.t3011 vp_p.t1554 vdd.t1445 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1925 out_p.t3010 vp_p.t1555 vdd.t1444 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1926 vdd.t1443 vp_p.t1556 out_p.t3009 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1927 vdd.t1442 vp_p.t1557 out_p.t3008 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1928 vdd.t1441 vp_p.t1558 out_p.t3007 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1929 vdd.t1440 vp_p.t1559 out_p.t3006 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1930 vdd.t1439 vp_p.t1560 out_p.t3005 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1931 vdd.t1438 vp_p.t1561 out_p.t3004 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1932 out_p.t3003 vp_p.t1562 vdd.t1437 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1933 vdd.t1436 vp_p.t1563 out_p.t3002 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1934 out_p.t3437 vp_n.t370 vss.t229 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1935 out_p.t283 vp_n.t371 vss.t228 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1936 vdd.t1435 vp_p.t1564 out_p.t3001 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1937 out_p.t3000 vp_p.t1565 vdd.t1434 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1938 vdd.t1433 vp_p.t1566 out_p.t2999 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1939 vdd.t1432 vp_p.t1567 out_p.t2998 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1940 out_p.t2997 vp_p.t1568 vdd.t1431 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1941 out_p.t2996 vp_p.t1569 vdd.t1430 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1942 out_p.t2995 vp_p.t1570 vdd.t1429 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1943 vdd.t1428 vp_p.t1571 out_p.t2994 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1944 out_p.t284 vp_n.t372 vss.t227 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1945 vdd.t1427 vp_p.t1572 out_p.t2993 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1946 vdd.t1426 vp_p.t1573 out_p.t2992 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1947 out_p.t2991 vp_p.t1574 vdd.t1425 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1948 vdd.t1424 vp_p.t1575 out_p.t2990 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1949 vdd.t1423 vp_p.t1576 out_p.t2989 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1950 vss.t226 vp_n.t373 out_p.t366 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1951 vdd.t1422 vp_p.t1577 out_p.t2988 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1952 vdd.t1421 vp_p.t1578 out_p.t2987 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1953 out_p.t2986 vp_p.t1579 vdd.t1420 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1954 vdd.t1419 vp_p.t1580 out_p.t2985 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1955 vdd.t1418 vp_p.t1581 out_p.t2984 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1956 vss.t225 vp_n.t374 out_p.t47 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1957 out_p.t49 vp_n.t375 vss.t224 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1958 out_p.t2983 vp_p.t1582 vdd.t1417 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1959 out_p.t2982 vp_p.t1583 vdd.t1416 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1960 out_p.t2981 vp_p.t1584 vdd.t1415 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1961 vss.t223 vp_n.t376 out_p.t365 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1962 out_p.t2980 vp_p.t1585 vdd.t1414 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1963 vdd.t1413 vp_p.t1586 out_p.t2979 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1964 out_p.t2978 vp_p.t1587 vdd.t1412 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1965 out_p.t216 vp_n.t377 vss.t222 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1966 out_p.t2977 vp_p.t1588 vdd.t1411 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1967 vdd.t1410 vp_p.t1589 out_p.t2976 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1968 out_p.t2975 vp_p.t1590 vdd.t1409 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1969 vdd.t1408 vp_p.t1591 out_p.t2974 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1970 vss.t221 vp_n.t378 out_p.t3436 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1971 out_p.t2973 vp_p.t1592 vdd.t1407 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1972 out_p.t280 vp_n.t379 vss.t220 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1973 vdd.t1406 vp_p.t1593 out_p.t2972 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1974 vdd.t1405 vp_p.t1594 out_p.t2971 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1975 vss.t219 vp_n.t380 out_p.t281 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1976 vdd.t1404 vp_p.t1595 out_p.t2970 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1977 out_p.t363 vp_n.t381 vss.t218 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1978 vdd.t1403 vp_p.t1596 out_p.t2969 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1979 out_p.t2968 vp_p.t1597 vdd.t1402 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1980 vss.t217 vp_n.t382 out_p.t50 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1981 out_p.t2967 vp_p.t1598 vdd.t1401 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1982 vdd.t1400 vp_p.t1599 out_p.t2966 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1983 out_p.t2965 vp_p.t1600 vdd.t1399 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1984 vdd.t1398 vp_p.t1601 out_p.t2964 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1985 vss.t216 vp_n.t383 out_p.t52 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1986 out_p.t362 vp_n.t384 vss.t215 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1987 vdd.t1397 vp_p.t1602 out_p.t2963 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1988 vdd.t1396 vp_p.t1603 out_p.t2962 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1989 out_p.t2961 vp_p.t1604 vdd.t1395 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1990 vdd.t1394 vp_p.t1605 out_p.t2960 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1991 vdd.t1393 vp_p.t1606 out_p.t2959 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1992 vss.t214 vp_n.t385 out_p.t215 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1993 vdd.t1392 vp_p.t1607 out_p.t2958 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1994 out_p.t2957 vp_p.t1608 vdd.t1391 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1995 vdd.t1390 vp_p.t1609 out_p.t2956 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1996 vdd.t1389 vp_p.t1610 out_p.t2955 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1997 out_p.t2954 vp_p.t1611 vdd.t1388 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1998 out_p.t3584 vp_n.t386 vss.t213 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1999 out_p.t2953 vp_p.t1612 vdd.t1387 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2000 out_p.t2952 vp_p.t1613 vdd.t1386 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2001 out_p.t2951 vp_p.t1614 vdd.t1385 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2002 out_p.t2950 vp_p.t1615 vdd.t1384 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2003 out_p.t2949 vp_p.t1616 vdd.t1383 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2004 out_p.t2948 vp_p.t1617 vdd.t1382 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2005 out_p.t2947 vp_p.t1618 vdd.t1381 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2006 vdd.t1380 vp_p.t1619 out_p.t2946 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2007 vdd.t1379 vp_p.t1620 out_p.t2945 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2008 out_p.t2944 vp_p.t1621 vdd.t1378 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2009 out_p.t276 vp_n.t387 vss.t212 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2010 out_p.t2943 vp_p.t1622 vdd.t1377 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2011 out_p.t2942 vp_p.t1623 vdd.t1376 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2012 out_p.t2941 vp_p.t1624 vdd.t1375 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2013 vdd.t1374 vp_p.t1625 out_p.t2940 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2014 vdd.t1373 vp_p.t1626 out_p.t2939 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2015 vss.t211 vp_n.t388 out_p.t277 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2016 out_p.t2938 vp_p.t1627 vdd.t1372 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2017 out_p.t2937 vp_p.t1628 vdd.t1371 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2018 out_p.t2936 vp_p.t1629 vdd.t1370 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2019 vdd.t1369 vp_p.t1630 out_p.t2935 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2020 out_p.t2934 vp_p.t1631 vdd.t1368 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2021 vss.t210 vp_n.t389 out_p.t360 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2022 vdd.t1367 vp_p.t1632 out_p.t2933 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2023 out_p.t2932 vp_p.t1633 vdd.t1366 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2024 out_p.t53 vp_n.t390 vss.t209 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2025 vdd.t1365 vp_p.t1634 out_p.t2931 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2026 vdd.t1364 vp_p.t1635 out_p.t2930 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2027 out_p.t55 vp_n.t391 vss.t208 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2028 vdd.t1363 vp_p.t1636 out_p.t2929 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2029 out_p.t2928 vp_p.t1637 vdd.t1362 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2030 vdd.t1361 vp_p.t1638 out_p.t2927 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2031 vdd.t1360 vp_p.t1639 out_p.t2926 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2032 vss.t207 vp_n.t392 out_p.t359 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2033 out_p.t2925 vp_p.t1640 vdd.t1359 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2034 vss.t206 vp_n.t393 out_p.t214 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2035 out_p.t2924 vp_p.t1641 vdd.t1358 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2036 out_p.t2923 vp_p.t1642 vdd.t1357 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2037 vdd.t1356 vp_p.t1643 out_p.t2922 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2038 out_p.t2921 vp_p.t1644 vdd.t1355 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2039 vdd.t1354 vp_p.t1645 out_p.t2920 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2040 out_p.t2919 vp_p.t1646 vdd.t1353 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2041 out_p.t2918 vp_p.t1647 vdd.t1352 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2042 out_p.t2917 vp_p.t1648 vdd.t1351 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2043 vdd.t1350 vp_p.t1649 out_p.t2916 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2044 out_p.t3583 vp_n.t394 vss.t205 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2045 vdd.t1349 vp_p.t1650 out_p.t2915 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2046 vdd.t1348 vp_p.t1651 out_p.t2914 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2047 out_p.t2913 vp_p.t1652 vdd.t1347 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2048 out_p.t2912 vp_p.t1653 vdd.t1346 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2049 out_p.t2911 vp_p.t1654 vdd.t1345 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2050 out_p.t2910 vp_p.t1655 vdd.t1344 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2051 out_p.t2909 vp_p.t1656 vdd.t1343 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2052 vdd.t1342 vp_p.t1657 out_p.t2908 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2053 out_p.t2907 vp_p.t1658 vdd.t1341 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2054 vss.t204 vp_n.t395 out_p.t274 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2055 vdd.t1340 vp_p.t1659 out_p.t2906 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2056 vdd.t1339 vp_p.t1660 out_p.t2905 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2057 vdd.t1338 vp_p.t1661 out_p.t2904 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2058 out_p.t2903 vp_p.t1662 vdd.t1337 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2059 vdd.t1336 vp_p.t1663 out_p.t2902 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2060 out_p.t2901 vp_p.t1664 vdd.t1335 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2061 out_p.t2900 vp_p.t1665 vdd.t1334 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2062 vdd.t1333 vp_p.t1666 out_p.t2899 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2063 vdd.t1332 vp_p.t1667 out_p.t2898 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2064 out_p.t2897 vp_p.t1668 vdd.t1331 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2065 vdd.t1330 vp_p.t1669 out_p.t2896 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2066 out_p.t2895 vp_p.t1670 vdd.t1329 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2067 out_p.t2894 vp_p.t1671 vdd.t1328 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2068 out_p.t2893 vp_p.t1672 vdd.t1327 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2069 out_p.t2892 vp_p.t1673 vdd.t1326 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2070 out_p.t2891 vp_p.t1674 vdd.t1325 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2071 out_p.t2890 vp_p.t1675 vdd.t1324 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2072 vdd.t1323 vp_p.t1676 out_p.t2889 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2073 vdd.t1322 vp_p.t1677 out_p.t2888 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2074 vdd.t1321 vp_p.t1678 out_p.t2887 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2075 vdd.t1320 vp_p.t1679 out_p.t2886 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2076 out_p.t2885 vp_p.t1680 vdd.t1319 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2077 vdd.t1318 vp_p.t1681 out_p.t2884 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2078 out_p.t2883 vp_p.t1682 vdd.t1317 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2079 out_p.t2882 vp_p.t1683 vdd.t1316 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2080 out_p.t2881 vp_p.t1684 vdd.t1315 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2081 vdd.t1314 vp_p.t1685 out_p.t2880 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2082 out_p.t2879 vp_p.t1686 vdd.t1313 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2083 vdd.t1312 vp_p.t1687 out_p.t2878 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2084 out_p.t2877 vp_p.t1688 vdd.t1311 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2085 vdd.t1310 vp_p.t1689 out_p.t2876 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2086 out_p.t2875 vp_p.t1690 vdd.t1309 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2087 out_p.t2874 vp_p.t1691 vdd.t1308 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2088 vdd.t1307 vp_p.t1692 out_p.t2873 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2089 vdd.t1306 vp_p.t1693 out_p.t2872 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2090 out_p.t2871 vp_p.t1694 vdd.t1305 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2091 vss.t203 vp_n.t396 out_p.t357 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2092 vdd.t1304 vp_p.t1695 out_p.t2870 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2093 out_p.t2869 vp_p.t1696 vdd.t1303 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2094 out_p.t2868 vp_p.t1697 vdd.t1302 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2095 out_p.t2867 vp_p.t1698 vdd.t1301 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2096 vdd.t1300 vp_p.t1699 out_p.t2866 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2097 vdd.t1299 vp_p.t1700 out_p.t2865 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2098 out_p.t2864 vp_p.t1701 vdd.t1298 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2099 vdd.t1297 vp_p.t1702 out_p.t2863 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2100 out_p.t56 vp_n.t397 vss.t202 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2101 vdd.t1296 vp_p.t1703 out_p.t2862 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2102 out_p.t2861 vp_p.t1704 vdd.t1295 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2103 vdd.t1294 vp_p.t1705 out_p.t2860 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2104 out_p.t2859 vp_p.t1706 vdd.t1293 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2105 out_p.t2858 vp_p.t1707 vdd.t1292 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2106 vdd.t1291 vp_p.t1708 out_p.t2857 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2107 out_p.t2856 vp_p.t1709 vdd.t1290 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2108 vdd.t1289 vp_p.t1710 out_p.t2855 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2109 out_p.t2854 vp_p.t1711 vdd.t1288 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2110 out_p.t2853 vp_p.t1712 vdd.t1287 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2111 vdd.t1286 vp_p.t1713 out_p.t2852 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2112 out_p.t2851 vp_p.t1714 vdd.t1285 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2113 out_p.t2850 vp_p.t1715 vdd.t1284 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2114 vdd.t1283 vp_p.t1716 out_p.t2849 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2115 vdd.t1282 vp_p.t1717 out_p.t2848 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2116 out_p.t2847 vp_p.t1718 vdd.t1281 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2117 out_p.t2846 vp_p.t1719 vdd.t1280 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2118 out_p.t58 vp_n.t398 vss.t201 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2119 out_p.t2845 vp_p.t1720 vdd.t1279 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2120 vdd.t1278 vp_p.t1721 out_p.t2844 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2121 out_p.t2843 vp_p.t1722 vdd.t1277 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2122 out_p.t2842 vp_p.t1723 vdd.t1276 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2123 vdd.t1275 vp_p.t1724 out_p.t2841 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2124 out_p.t2840 vp_p.t1725 vdd.t1274 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2125 out_p.t2839 vp_p.t1726 vdd.t1273 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2126 vdd.t1272 vp_p.t1727 out_p.t2838 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2127 vdd.t1271 vp_p.t1728 out_p.t2837 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2128 out_p.t2836 vp_p.t1729 vdd.t1270 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2129 vdd.t1269 vp_p.t1730 out_p.t2835 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2130 out_p.t2834 vp_p.t1731 vdd.t1268 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2131 vdd.t1267 vp_p.t1732 out_p.t2833 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2132 vdd.t1266 vp_p.t1733 out_p.t2832 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2133 vdd.t1265 vp_p.t1734 out_p.t2831 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2134 vdd.t1264 vp_p.t1735 out_p.t2830 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2135 vdd.t1263 vp_p.t1736 out_p.t2829 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2136 out_p.t2828 vp_p.t1737 vdd.t1262 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2137 vdd.t1261 vp_p.t1738 out_p.t2827 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2138 vdd.t1260 vp_p.t1739 out_p.t2826 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2139 vdd.t1259 vp_p.t1740 out_p.t2825 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2140 out_p.t2824 vp_p.t1741 vdd.t1258 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2141 vdd.t1257 vp_p.t1742 out_p.t2823 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2142 out_p.t2822 vp_p.t1743 vdd.t1256 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2143 vdd.t1255 vp_p.t1744 out_p.t2821 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2144 out_p.t2820 vp_p.t1745 vdd.t1254 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2145 out_p.t2819 vp_p.t1746 vdd.t1253 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2146 out_p.t2818 vp_p.t1747 vdd.t1252 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2147 out_p.t2817 vp_p.t1748 vdd.t1251 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2148 out_p.t2816 vp_p.t1749 vdd.t1250 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2149 vdd.t1249 vp_p.t1750 out_p.t2815 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2150 vdd.t1248 vp_p.t1751 out_p.t2814 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2151 out_p.t2813 vp_p.t1752 vdd.t1247 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2152 out_p.t2812 vp_p.t1753 vdd.t1246 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2153 out_p.t2811 vp_p.t1754 vdd.t1245 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2154 out_p.t2810 vp_p.t1755 vdd.t1244 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2155 vss.t200 vp_n.t399 out_p.t272 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2156 out_p.t2809 vp_p.t1756 vdd.t1243 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2157 out_p.t2808 vp_p.t1757 vdd.t1242 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2158 out_p.t2807 vp_p.t1758 vdd.t1241 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2159 out_p.t2806 vp_p.t1759 vdd.t1240 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2160 vdd.t1239 vp_p.t1760 out_p.t2805 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2161 vdd.t1238 vp_p.t1761 out_p.t2804 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2162 out_p.t2803 vp_p.t1762 vdd.t1237 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2163 vdd.t1236 vp_p.t1763 out_p.t2802 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2164 vdd.t1235 vp_p.t1764 out_p.t2801 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2165 out_p.t2800 vp_p.t1765 vdd.t1234 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2166 out_p.t2799 vp_p.t1766 vdd.t1233 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2167 vdd.t1232 vp_p.t1767 out_p.t2798 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2168 vdd.t1231 vp_p.t1768 out_p.t2797 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2169 out_p.t2796 vp_p.t1769 vdd.t1230 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2170 vdd.t1229 vp_p.t1770 out_p.t2795 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2171 out_p.t2794 vp_p.t1771 vdd.t1228 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2172 vdd.t1227 vp_p.t1772 out_p.t2793 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2173 out_p.t2792 vp_p.t1773 vdd.t1226 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2174 out_p.t2791 vp_p.t1774 vdd.t1225 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2175 vdd.t1224 vp_p.t1775 out_p.t2790 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2176 out_p.t2789 vp_p.t1776 vdd.t1223 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2177 out_p.t2788 vp_p.t1777 vdd.t1222 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2178 vdd.t1221 vp_p.t1778 out_p.t2787 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2179 out_p.t2786 vp_p.t1779 vdd.t1220 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2180 out_p.t2785 vp_p.t1780 vdd.t1219 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2181 vdd.t1218 vp_p.t1781 out_p.t2784 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2182 vdd.t1217 vp_p.t1782 out_p.t2783 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2183 vdd.t1216 vp_p.t1783 out_p.t2782 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2184 out_p.t2781 vp_p.t1784 vdd.t1215 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2185 out_p.t2780 vp_p.t1785 vdd.t1214 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2186 out_p.t2779 vp_p.t1786 vdd.t1213 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2187 out_p.t2778 vp_p.t1787 vdd.t1212 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2188 out_p.t2777 vp_p.t1788 vdd.t1211 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2189 out_p.t2776 vp_p.t1789 vdd.t1210 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2190 out_p.t2775 vp_p.t1790 vdd.t1209 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2191 out_p.t2774 vp_p.t1791 vdd.t1208 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2192 vdd.t1207 vp_p.t1792 out_p.t2773 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2193 out_p.t2772 vp_p.t1793 vdd.t1206 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2194 vdd.t1205 vp_p.t1794 out_p.t2771 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2195 out_p.t2770 vp_p.t1795 vdd.t1204 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2196 out_p.t2769 vp_p.t1796 vdd.t1203 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2197 vdd.t1202 vp_p.t1797 out_p.t2768 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2198 out_p.t2767 vp_p.t1798 vdd.t1201 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2199 out_p.t2766 vp_p.t1799 vdd.t1200 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2200 out_p.t2765 vp_p.t1800 vdd.t1199 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2201 out_p.t2764 vp_p.t1801 vdd.t1198 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2202 vdd.t1197 vp_p.t1802 out_p.t2763 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2203 vdd.t1196 vp_p.t1803 out_p.t2762 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2204 out_p.t2761 vp_p.t1804 vdd.t1195 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2205 out_p.t2760 vp_p.t1805 vdd.t1194 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2206 out_p.t2759 vp_p.t1806 vdd.t1193 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2207 out_p.t2758 vp_p.t1807 vdd.t1192 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2208 out_p.t2757 vp_p.t1808 vdd.t1191 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2209 out_p.t2756 vp_p.t1809 vdd.t1190 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2210 out_p.t2755 vp_p.t1810 vdd.t1189 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2211 out_p.t2754 vp_p.t1811 vdd.t1188 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2212 vdd.t1187 vp_p.t1812 out_p.t2753 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2213 out_p.t2752 vp_p.t1813 vdd.t1186 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2214 out_p.t2751 vp_p.t1814 vdd.t1185 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2215 vdd.t1184 vp_p.t1815 out_p.t2750 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2216 vdd.t1183 vp_p.t1816 out_p.t2749 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2217 vdd.t1182 vp_p.t1817 out_p.t2748 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2218 vdd.t1181 vp_p.t1818 out_p.t2747 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2219 out_p.t2746 vp_p.t1819 vdd.t1180 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2220 vdd.t1179 vp_p.t1820 out_p.t2745 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2221 vdd.t1178 vp_p.t1821 out_p.t2744 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2222 out_p.t2743 vp_p.t1822 vdd.t1177 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2223 vdd.t1176 vp_p.t1823 out_p.t2742 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2224 out_p.t2741 vp_p.t1824 vdd.t1175 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2225 vdd.t1174 vp_p.t1825 out_p.t2740 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2226 out_p.t2739 vp_p.t1826 vdd.t1173 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2227 out_p.t2738 vp_p.t1827 vdd.t1172 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2228 vdd.t1171 vp_p.t1828 out_p.t2737 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2229 out_p.t2736 vp_p.t1829 vdd.t1170 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2230 out_p.t2735 vp_p.t1830 vdd.t1169 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2231 vdd.t1168 vp_p.t1831 out_p.t2734 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2232 out_p.t2733 vp_p.t1832 vdd.t1167 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2233 out_p.t2732 vp_p.t1833 vdd.t1166 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2234 out_p.t2731 vp_p.t1834 vdd.t1165 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2235 vdd.t1164 vp_p.t1835 out_p.t2730 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2236 out_p.t2729 vp_p.t1836 vdd.t1163 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2237 out_p.t2728 vp_p.t1837 vdd.t1162 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2238 out_p.t2727 vp_p.t1838 vdd.t1161 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2239 out_p.t2726 vp_p.t1839 vdd.t1160 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2240 vdd.t1159 vp_p.t1840 out_p.t2725 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2241 vdd.t1158 vp_p.t1841 out_p.t2724 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2242 out_p.t2723 vp_p.t1842 vdd.t1157 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2243 out_p.t2722 vp_p.t1843 vdd.t1156 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2244 vdd.t1155 vp_p.t1844 out_p.t2721 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2245 out_p.t2720 vp_p.t1845 vdd.t1154 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2246 out_p.t2719 vp_p.t1846 vdd.t1153 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2247 vdd.t1152 vp_p.t1847 out_p.t2718 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2248 out_p.t2717 vp_p.t1848 vdd.t1151 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2249 vdd.t1150 vp_p.t1849 out_p.t2716 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2250 vdd.t1149 vp_p.t1850 out_p.t2715 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2251 vdd.t1148 vp_p.t1851 out_p.t2714 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2252 out_p.t2713 vp_p.t1852 vdd.t1147 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2253 vdd.t1146 vp_p.t1853 out_p.t2712 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2254 out_p.t2711 vp_p.t1854 vdd.t1145 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2255 out_p.t2710 vp_p.t1855 vdd.t1144 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2256 out_p.t2709 vp_p.t1856 vdd.t1143 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2257 out_p.t2708 vp_p.t1857 vdd.t1142 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2258 out_p.t2707 vp_p.t1858 vdd.t1141 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2259 out_p.t2706 vp_p.t1859 vdd.t1140 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2260 out_p.t2705 vp_p.t1860 vdd.t1139 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2261 out_p.t2704 vp_p.t1861 vdd.t1138 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2262 vdd.t1137 vp_p.t1862 out_p.t2703 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2263 out_p.t2702 vp_p.t1863 vdd.t1136 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2264 vdd.t1135 vp_p.t1864 out_p.t2701 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2265 out_p.t2700 vp_p.t1865 vdd.t1134 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2266 vdd.t1133 vp_p.t1866 out_p.t2699 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2267 vdd.t1132 vp_p.t1867 out_p.t2698 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2268 out_p.t2697 vp_p.t1868 vdd.t1131 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2269 out_p.t2696 vp_p.t1869 vdd.t1130 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2270 vdd.t1129 vp_p.t1870 out_p.t2695 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2271 vdd.t1128 vp_p.t1871 out_p.t2694 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2272 out_p.t2693 vp_p.t1872 vdd.t1127 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2273 vdd.t1126 vp_p.t1873 out_p.t2692 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2274 vdd.t1125 vp_p.t1874 out_p.t2691 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2275 out_p.t2690 vp_p.t1875 vdd.t1124 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2276 out_p.t2689 vp_p.t1876 vdd.t1123 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2277 out_p.t2688 vp_p.t1877 vdd.t1122 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2278 out_p.t2687 vp_p.t1878 vdd.t1121 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2279 out_p.t2686 vp_p.t1879 vdd.t1120 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2280 out_p.t2685 vp_p.t1880 vdd.t1119 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2281 vdd.t1118 vp_p.t1881 out_p.t2684 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2282 out_p.t2683 vp_p.t1882 vdd.t1117 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2283 vdd.t1116 vp_p.t1883 out_p.t2682 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2284 out_p.t356 vp_n.t400 vss.t199 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2285 vdd.t1115 vp_p.t1884 out_p.t2681 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2286 out_p.t2680 vp_p.t1885 vdd.t1114 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2287 vdd.t1113 vp_p.t1886 out_p.t2679 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2288 out_p.t2678 vp_p.t1887 vdd.t1112 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2289 out_p.t2677 vp_p.t1888 vdd.t1111 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2290 vdd.t1110 vp_p.t1889 out_p.t2676 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2291 vdd.t1109 vp_p.t1890 out_p.t2675 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2292 vdd.t1108 vp_p.t1891 out_p.t2674 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2293 out_p.t2673 vp_p.t1892 vdd.t1107 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2294 out_p.t2672 vp_p.t1893 vdd.t1106 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2295 out_p.t2671 vp_p.t1894 vdd.t1105 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2296 vdd.t1104 vp_p.t1895 out_p.t2670 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2297 vdd.t1103 vp_p.t1896 out_p.t2669 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2298 vdd.t1102 vp_p.t1897 out_p.t2668 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2299 vdd.t1101 vp_p.t1898 out_p.t2667 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2300 vdd.t1100 vp_p.t1899 out_p.t2666 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2301 out_p.t2665 vp_p.t1900 vdd.t1099 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2302 vdd.t1098 vp_p.t1901 out_p.t2664 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2303 out_p.t2663 vp_p.t1902 vdd.t1097 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2304 vdd.t1096 vp_p.t1903 out_p.t2662 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2305 out_p.t2661 vp_p.t1904 vdd.t1095 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2306 out_p.t2660 vp_p.t1905 vdd.t1094 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2307 vdd.t1093 vp_p.t1906 out_p.t2659 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2308 out_p.t2658 vp_p.t1907 vdd.t1092 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2309 vdd.t1091 vp_p.t1908 out_p.t2657 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2310 vdd.t1090 vp_p.t1909 out_p.t2656 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2311 out_p.t2655 vp_p.t1910 vdd.t1089 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2312 out_p.t2654 vp_p.t1911 vdd.t1088 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2313 out_p.t2653 vp_p.t1912 vdd.t1087 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2314 vdd.t1086 vp_p.t1913 out_p.t2652 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2315 out_p.t2651 vp_p.t1914 vdd.t1085 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2316 out_p.t2650 vp_p.t1915 vdd.t1084 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2317 out_p.t2649 vp_p.t1916 vdd.t1083 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2318 vdd.t1082 vp_p.t1917 out_p.t2648 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2319 out_p.t2647 vp_p.t1918 vdd.t1081 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2320 out_p.t2646 vp_p.t1919 vdd.t1080 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2321 vdd.t1079 vp_p.t1920 out_p.t2645 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2322 out_p.t2644 vp_p.t1921 vdd.t1078 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2323 vdd.t1077 vp_p.t1922 out_p.t2643 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2324 out_p.t2642 vp_p.t1923 vdd.t1076 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2325 out_p.t2641 vp_p.t1924 vdd.t1075 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2326 vdd.t1074 vp_p.t1925 out_p.t2640 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2327 vdd.t1073 vp_p.t1926 out_p.t2639 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2328 out_p.t2638 vp_p.t1927 vdd.t1072 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2329 out_p.t2637 vp_p.t1928 vdd.t1071 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2330 vdd.t1070 vp_p.t1929 out_p.t2636 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2331 vdd.t1069 vp_p.t1930 out_p.t2635 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2332 vdd.t1068 vp_p.t1931 out_p.t2634 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2333 out_p.t2633 vp_p.t1932 vdd.t1067 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2334 vdd.t1066 vp_p.t1933 out_p.t2632 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2335 out_p.t2631 vp_p.t1934 vdd.t1065 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2336 vdd.t1064 vp_p.t1935 out_p.t2630 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2337 vdd.t1063 vp_p.t1936 out_p.t2629 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2338 vdd.t1062 vp_p.t1937 out_p.t2628 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2339 vdd.t1061 vp_p.t1938 out_p.t2627 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2340 out_p.t2626 vp_p.t1939 vdd.t1060 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2341 out_p.t2625 vp_p.t1940 vdd.t1059 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2342 out_p.t2624 vp_p.t1941 vdd.t1058 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2343 vdd.t1057 vp_p.t1942 out_p.t2623 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2344 vdd.t1056 vp_p.t1943 out_p.t2622 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2345 vdd.t1055 vp_p.t1944 out_p.t2621 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2346 out_p.t2620 vp_p.t1945 vdd.t1054 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2347 vdd.t1053 vp_p.t1946 out_p.t2619 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2348 vdd.t1052 vp_p.t1947 out_p.t2618 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2349 vdd.t1051 vp_p.t1948 out_p.t2617 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2350 out_p.t2616 vp_p.t1949 vdd.t1050 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2351 vdd.t1049 vp_p.t1950 out_p.t2615 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2352 out_p.t2614 vp_p.t1951 vdd.t1048 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2353 vdd.t1047 vp_p.t1952 out_p.t2613 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2354 vdd.t1046 vp_p.t1953 out_p.t2612 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2355 out_p.t2611 vp_p.t1954 vdd.t1045 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2356 vdd.t1044 vp_p.t1955 out_p.t2610 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2357 vdd.t1043 vp_p.t1956 out_p.t2609 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2358 vdd.t1042 vp_p.t1957 out_p.t2608 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2359 out_p.t2607 vp_p.t1958 vdd.t1041 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2360 vdd.t1040 vp_p.t1959 out_p.t2606 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2361 vdd.t1039 vp_p.t1960 out_p.t2605 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2362 out_p.t2604 vp_p.t1961 vdd.t1038 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2363 out_p.t2603 vp_p.t1962 vdd.t1037 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2364 out_p.t2602 vp_p.t1963 vdd.t1036 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2365 out_p.t2601 vp_p.t1964 vdd.t1035 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2366 vss.t198 vp_n.t401 out_p.t213 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2367 vdd.t1034 vp_p.t1965 out_p.t2600 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2368 vdd.t1033 vp_p.t1966 out_p.t2599 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2369 out_p.t2598 vp_p.t1967 vdd.t1032 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2370 vdd.t1031 vp_p.t1968 out_p.t2597 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2371 out_p.t2596 vp_p.t1969 vdd.t1030 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2372 vdd.t1029 vp_p.t1970 out_p.t2595 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2373 out_p.t2594 vp_p.t1971 vdd.t1028 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2374 vdd.t1027 vp_p.t1972 out_p.t2593 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2375 vdd.t1026 vp_p.t1973 out_p.t2592 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2376 out_p.t2591 vp_p.t1974 vdd.t1025 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2377 vdd.t1024 vp_p.t1975 out_p.t2590 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2378 vdd.t1023 vp_p.t1976 out_p.t2589 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2379 vdd.t1022 vp_p.t1977 out_p.t2588 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2380 vdd.t1021 vp_p.t1978 out_p.t2587 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2381 vdd.t1020 vp_p.t1979 out_p.t2586 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2382 vdd.t1019 vp_p.t1980 out_p.t2585 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2383 vdd.t1018 vp_p.t1981 out_p.t2584 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2384 out_p.t2583 vp_p.t1982 vdd.t1017 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2385 out_p.t2582 vp_p.t1983 vdd.t1016 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2386 out_p.t2581 vp_p.t1984 vdd.t1015 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2387 vdd.t1014 vp_p.t1985 out_p.t2580 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2388 vdd.t1013 vp_p.t1986 out_p.t2579 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2389 vdd.t1012 vp_p.t1987 out_p.t2578 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2390 out_p.t2577 vp_p.t1988 vdd.t1011 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2391 vdd.t1010 vp_p.t1989 out_p.t2576 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2392 out_p.t2575 vp_p.t1990 vdd.t1009 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2393 out_p.t2574 vp_p.t1991 vdd.t1008 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2394 vdd.t1007 vp_p.t1992 out_p.t2573 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2395 out_p.t2572 vp_p.t1993 vdd.t1006 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2396 vdd.t1005 vp_p.t1994 out_p.t2571 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2397 vdd.t1004 vp_p.t1995 out_p.t2570 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2398 out_p.t2569 vp_p.t1996 vdd.t1003 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2399 out_p.t2568 vp_p.t1997 vdd.t1002 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2400 vdd.t1001 vp_p.t1998 out_p.t2567 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2401 out_p.t2566 vp_p.t1999 vdd.t1000 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2402 out_p.t2565 vp_p.t2000 vdd.t999 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2403 out_p.t2564 vp_p.t2001 vdd.t998 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2404 vdd.t997 vp_p.t2002 out_p.t2563 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2405 vdd.t996 vp_p.t2003 out_p.t2562 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2406 out_p.t2561 vp_p.t2004 vdd.t995 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2407 vdd.t994 vp_p.t2005 out_p.t2560 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2408 out_p.t2559 vp_p.t2006 vdd.t993 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2409 vdd.t992 vp_p.t2007 out_p.t2558 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2410 vdd.t991 vp_p.t2008 out_p.t2557 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2411 out_p.t2556 vp_p.t2009 vdd.t990 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2412 out_p.t2555 vp_p.t2010 vdd.t989 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2413 vdd.t988 vp_p.t2011 out_p.t2554 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2414 out_p.t2553 vp_p.t2012 vdd.t987 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2415 vdd.t986 vp_p.t2013 out_p.t2552 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2416 out_p.t2551 vp_p.t2014 vdd.t985 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2417 vdd.t984 vp_p.t2015 out_p.t2550 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2418 out_p.t2549 vp_p.t2016 vdd.t983 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2419 out_p.t2548 vp_p.t2017 vdd.t982 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2420 vdd.t981 vp_p.t2018 out_p.t2547 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2421 out_p.t2546 vp_p.t2019 vdd.t980 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2422 vdd.t979 vp_p.t2020 out_p.t2545 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2423 out_p.t2544 vp_p.t2021 vdd.t978 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2424 out_p.t2543 vp_p.t2022 vdd.t977 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2425 out_p.t2542 vp_p.t2023 vdd.t976 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2426 vdd.t975 vp_p.t2024 out_p.t2541 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2427 vdd.t974 vp_p.t2025 out_p.t2540 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2428 out_p.t2539 vp_p.t2026 vdd.t973 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2429 vdd.t972 vp_p.t2027 out_p.t2538 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2430 out_p.t2537 vp_p.t2028 vdd.t971 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2431 vdd.t970 vp_p.t2029 out_p.t2536 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2432 vdd.t969 vp_p.t2030 out_p.t2535 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2433 vdd.t968 vp_p.t2031 out_p.t2534 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2434 out_p.t2533 vp_p.t2032 vdd.t967 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2435 vdd.t966 vp_p.t2033 out_p.t2532 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2436 out_p.t3480 vp_n.t402 vss.t197 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2437 out_p.t2531 vp_p.t2034 vdd.t965 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2438 vdd.t964 vp_p.t2035 out_p.t2530 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2439 vdd.t963 vp_p.t2036 out_p.t2529 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2440 vdd.t962 vp_p.t2037 out_p.t2528 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2441 vdd.t961 vp_p.t2038 out_p.t2527 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2442 out_p.t2526 vp_p.t2039 vdd.t960 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2443 vss.t196 vp_n.t403 out_p.t271 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2444 out_p.t2525 vp_p.t2040 vdd.t959 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2445 vdd.t958 vp_p.t2041 out_p.t2524 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2446 vdd.t957 vp_p.t2042 out_p.t2523 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2447 vdd.t956 vp_p.t2043 out_p.t2522 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2448 vdd.t955 vp_p.t2044 out_p.t2521 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2449 out_p.t2520 vp_p.t2045 vdd.t954 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2450 out_p.t2519 vp_p.t2046 vdd.t953 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2451 out_p.t2518 vp_p.t2047 vdd.t952 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2452 vdd.t951 vp_p.t2048 out_p.t1190 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2453 out_p.t1189 vp_p.t2049 vdd.t950 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2454 vdd.t949 vp_p.t2050 out_p.t1188 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2455 vdd.t948 vp_p.t2051 out_p.t1187 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2456 out_p.t1186 vp_p.t2052 vdd.t947 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2457 vdd.t946 vp_p.t2053 out_p.t1185 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2458 out_p.t1184 vp_p.t2054 vdd.t945 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2459 vdd.t944 vp_p.t2055 out_p.t1183 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2460 vdd.t943 vp_p.t2056 out_p.t1182 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2461 out_p.t1181 vp_p.t2057 vdd.t942 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2462 out_p.t1180 vp_p.t2058 vdd.t941 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2463 out_p.t1179 vp_p.t2059 vdd.t940 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2464 out_p.t1178 vp_p.t2060 vdd.t939 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2465 vdd.t938 vp_p.t2061 out_p.t1177 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2466 out_p.t1176 vp_p.t2062 vdd.t937 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2467 vdd.t936 vp_p.t2063 out_p.t1175 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2468 out_p.t1174 vp_p.t2064 vdd.t935 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2469 out_p.t1173 vp_p.t2065 vdd.t934 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2470 out_p.t1172 vp_p.t2066 vdd.t933 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2471 out_p.t1171 vp_p.t2067 vdd.t932 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2472 vdd.t931 vp_p.t2068 out_p.t1170 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2473 out_p.t354 vp_n.t404 vss.t195 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2474 vdd.t930 vp_p.t2069 out_p.t1169 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2475 vdd.t929 vp_p.t2070 out_p.t1168 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2476 out_p.t155 vp_n.t405 vss.t194 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2477 vdd.t928 vp_p.t2071 out_p.t1167 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2478 out_p.t1166 vp_p.t2072 vdd.t927 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2479 vdd.t926 vp_p.t2073 out_p.t1165 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2480 vdd.t925 vp_p.t2074 out_p.t1164 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2481 vdd.t924 vp_p.t2075 out_p.t1163 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2482 out_p.t1162 vp_p.t2076 vdd.t923 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2483 out_p.t1161 vp_p.t2077 vdd.t922 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2484 vdd.t921 vp_p.t2078 out_p.t1160 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2485 out_p.t1159 vp_p.t2079 vdd.t920 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2486 out_p.t1158 vp_p.t2080 vdd.t919 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2487 vss.t193 vp_n.t406 out_p.t59 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2488 out_p.t1157 vp_p.t2081 vdd.t918 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2489 out_p.t1156 vp_p.t2082 vdd.t917 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2490 vdd.t916 vp_p.t2083 out_p.t1155 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2491 vdd.t915 vp_p.t2084 out_p.t1154 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2492 out_p.t1153 vp_p.t2085 vdd.t914 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2493 vdd.t913 vp_p.t2086 out_p.t1152 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2494 out_p.t1151 vp_p.t2087 vdd.t912 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2495 out_p.t61 vp_n.t407 vss.t192 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2496 vdd.t911 vp_p.t2088 out_p.t1150 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2497 out_p.t1149 vp_p.t2089 vdd.t910 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2498 out_p.t212 vp_n.t408 vss.t191 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2499 vdd.t909 vp_p.t2090 out_p.t1148 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2500 out_p.t1147 vp_p.t2091 vdd.t908 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2501 vdd.t907 vp_p.t2092 out_p.t1146 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2502 vdd.t906 vp_p.t2093 out_p.t1145 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2503 vdd.t905 vp_p.t2094 out_p.t1144 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2504 out_p.t1143 vp_p.t2095 vdd.t904 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2505 vdd.t903 vp_p.t2096 out_p.t1142 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2506 out_p.t1141 vp_p.t2097 vdd.t902 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2507 out_p.t1140 vp_p.t2098 vdd.t901 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2508 vdd.t900 vp_p.t2099 out_p.t1139 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2509 out_p.t1138 vp_p.t2100 vdd.t899 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2510 vss.t190 vp_n.t409 out_p.t3479 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2511 out_p.t1137 vp_p.t2101 vdd.t898 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2512 vdd.t897 vp_p.t2102 out_p.t1136 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2513 out_p.t1135 vp_p.t2103 vdd.t896 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2514 out_p.t269 vp_n.t410 vss.t189 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2515 out_p.t1134 vp_p.t2104 vdd.t895 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2516 vdd.t894 vp_p.t2105 out_p.t1133 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2517 out_p.t1132 vp_p.t2106 vdd.t893 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2518 vdd.t892 vp_p.t2107 out_p.t1131 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2519 out_p.t62 vp_n.t411 vss.t188 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2520 vdd.t891 vp_p.t2108 out_p.t1130 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2521 vdd.t890 vp_p.t2109 out_p.t1129 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2522 vdd.t889 vp_p.t2110 out_p.t1128 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2523 vdd.t888 vp_p.t2111 out_p.t1127 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2524 out_p.t1126 vp_p.t2112 vdd.t887 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2525 vdd.t886 vp_p.t2113 out_p.t1125 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2526 out_p.t1124 vp_p.t2114 vdd.t885 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2527 out_p.t1123 vp_p.t2115 vdd.t884 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2528 out_p.t1122 vp_p.t2116 vdd.t883 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2529 vdd.t882 vp_p.t2117 out_p.t1121 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2530 vdd.t881 vp_p.t2118 out_p.t1120 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2531 vdd.t880 vp_p.t2119 out_p.t1119 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2532 vss.t187 vp_n.t412 out_p.t211 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2533 out_p.t1118 vp_p.t2120 vdd.t879 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2534 out_p.t1117 vp_p.t2121 vdd.t878 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2535 out_p.t1116 vp_p.t2122 vdd.t877 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2536 vdd.t876 vp_p.t2123 out_p.t1115 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2537 vdd.t875 vp_p.t2124 out_p.t1114 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2538 vdd.t874 vp_p.t2125 out_p.t1113 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2539 out_p.t1112 vp_p.t2126 vdd.t873 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2540 vdd.t872 vp_p.t2127 out_p.t1111 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2541 vdd.t871 vp_p.t2128 out_p.t1110 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2542 out_p.t3441 vp_n.t413 vss.t186 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2543 out_p.t1109 vp_p.t2129 vdd.t870 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2544 vdd.t869 vp_p.t2130 out_p.t1108 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2545 vdd.t868 vp_p.t2131 out_p.t1107 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2546 vdd.t867 vp_p.t2132 out_p.t1106 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2547 out_p.t1105 vp_p.t2133 vdd.t866 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2548 out_p.t1104 vp_p.t2134 vdd.t865 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2549 vdd.t864 vp_p.t2135 out_p.t1103 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2550 out_p.t1102 vp_p.t2136 vdd.t863 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2551 vss.t185 vp_n.t414 out_p.t64 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2552 vdd.t862 vp_p.t2137 out_p.t1101 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2553 vdd.t861 vp_p.t2138 out_p.t1100 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2554 out_p.t1099 vp_p.t2139 vdd.t860 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2555 vss.t184 vp_n.t415 out_p.t66 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2556 vss.t183 vp_n.t416 out_p.t65 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2557 out_p.t1098 vp_p.t2140 vdd.t859 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2558 vdd.t858 vp_p.t2141 out_p.t1097 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2559 out_p.t1096 vp_p.t2142 vdd.t857 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2560 vdd.t856 vp_p.t2143 out_p.t1095 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2561 vdd.t855 vp_p.t2144 out_p.t1094 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2562 vdd.t854 vp_p.t2145 out_p.t1093 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2563 out_p.t1092 vp_p.t2146 vdd.t853 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2564 out_p.t1091 vp_p.t2147 vdd.t852 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2565 out_p.t1090 vp_p.t2148 vdd.t851 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2566 vdd.t850 vp_p.t2149 out_p.t1089 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2567 vdd.t849 vp_p.t2150 out_p.t1088 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2568 out_p.t1087 vp_p.t2151 vdd.t848 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2569 out_p.t210 vp_n.t417 vss.t182 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2570 out_p.t1086 vp_p.t2152 vdd.t847 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2571 vdd.t846 vp_p.t2153 out_p.t1085 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2572 vdd.t845 vp_p.t2154 out_p.t1084 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2573 vdd.t844 vp_p.t2155 out_p.t1083 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2574 vdd.t843 vp_p.t2156 out_p.t1082 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2575 out_p.t1081 vp_p.t2157 vdd.t842 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2576 vss.t181 vp_n.t418 out_p.t3440 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2577 out_p.t1080 vp_p.t2158 vdd.t841 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2578 vss.t180 vp_n.t419 out_p.t67 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2579 out_p.t1079 vp_p.t2159 vdd.t840 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2580 out_p.t209 vp_n.t420 vss.t179 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2581 out_p.t1078 vp_p.t2160 vdd.t839 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2582 vdd.t838 vp_p.t2161 out_p.t1077 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2583 vss.t178 vp_n.t421 out_p.t3592 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2584 vdd.t837 vp_p.t2162 out_p.t1076 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2585 out_p.t1075 vp_p.t2163 vdd.t836 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2586 out_p.t1074 vp_p.t2164 vdd.t835 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2587 vdd.t834 vp_p.t2165 out_p.t1073 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2588 out_p.t1072 vp_p.t2166 vdd.t833 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2589 out_p.t70 vp_n.t422 vss.t177 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2590 out_p.t1071 vp_p.t2167 vdd.t832 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2591 vdd.t831 vp_p.t2168 out_p.t1070 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2592 vdd.t830 vp_p.t2169 out_p.t1069 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2593 vss.t176 vp_n.t423 out_p.t72 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2594 out_p.t1068 vp_p.t2170 vdd.t829 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2595 vdd.t828 vp_p.t2171 out_p.t1067 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2596 out_p.t1066 vp_p.t2172 vdd.t827 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2597 vdd.t826 vp_p.t2173 out_p.t1065 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2598 out_p.t1064 vp_p.t2174 vdd.t825 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2599 vss.t175 vp_n.t424 out_p.t208 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2600 out_p.t1063 vp_p.t2175 vdd.t824 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2601 out_p.t1062 vp_p.t2176 vdd.t823 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2602 out_p.t1061 vp_p.t2177 vdd.t822 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2603 vdd.t821 vp_p.t2178 out_p.t1060 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2604 out_p.t1059 vp_p.t2179 vdd.t820 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2605 vdd.t819 vp_p.t2180 out_p.t1058 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2606 out_p.t3591 vp_n.t425 vss.t174 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2607 out_p.t1057 vp_p.t2181 vdd.t818 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2608 vdd.t817 vp_p.t2182 out_p.t1056 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2609 vdd.t816 vp_p.t2183 out_p.t1055 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2610 vdd.t815 vp_p.t2184 out_p.t1054 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2611 out_p.t1053 vp_p.t2185 vdd.t814 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2612 out_p.t73 vp_n.t426 vss.t173 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2613 vdd.t813 vp_p.t2186 out_p.t1052 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2614 out_p.t74 vp_n.t427 vss.t172 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2615 out_p.t207 vp_n.t428 vss.t171 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2616 vdd.t812 vp_p.t2187 out_p.t1051 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2617 vdd.t811 vp_p.t2188 out_p.t1050 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2618 out_p.t3449 vp_n.t429 vss.t170 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2619 out_p.t75 vp_n.t430 vss.t169 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2620 out_p.t1049 vp_p.t2189 vdd.t810 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2621 vdd.t809 vp_p.t2190 out_p.t1048 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2622 vss.t168 vp_n.t431 out_p.t76 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2623 out_p.t206 vp_n.t432 vss.t167 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2624 out_p.t1047 vp_p.t2191 vdd.t808 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2625 vdd.t807 vp_p.t2192 out_p.t1046 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2626 vdd.t806 vp_p.t2193 out_p.t1045 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2627 out_p.t3448 vp_n.t433 vss.t166 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2628 vss.t165 vp_n.t434 out_p.t77 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2629 vdd.t805 vp_p.t2194 out_p.t1044 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2630 out_p.t1043 vp_p.t2195 vdd.t804 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2631 out_p.t79 vp_n.t435 vss.t164 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2632 vss.t163 vp_n.t436 out_p.t205 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2633 out_p.t1042 vp_p.t2196 vdd.t803 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2634 out_p.t1041 vp_p.t2197 vdd.t802 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2635 vdd.t801 vp_p.t2198 out_p.t1040 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2636 out_p.t3482 vp_n.t437 vss.t162 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2637 out_p.t1039 vp_p.t2199 vdd.t800 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2638 vdd.t799 vp_p.t2200 out_p.t1038 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2639 out_p.t80 vp_n.t438 vss.t161 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2640 vdd.t798 vp_p.t2201 out_p.t1037 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2641 out_p.t1036 vp_p.t2202 vdd.t797 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2642 out_p.t204 vp_n.t439 vss.t160 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2643 out_p.t1035 vp_p.t2203 vdd.t796 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2644 out_p.t1034 vp_p.t2204 vdd.t795 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2645 vss.t159 vp_n.t440 out_p.t3481 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2646 out_p.t1033 vp_p.t2205 vdd.t794 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2647 vss.t158 vp_n.t441 out_p.t81 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2648 out_p.t203 vp_n.t442 vss.t157 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2649 vdd.t793 vp_p.t2206 out_p.t1032 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2650 vdd.t792 vp_p.t2207 out_p.t1031 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2651 vdd.t791 vp_p.t2208 out_p.t1030 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2652 vdd.t790 vp_p.t2209 out_p.t1029 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2653 out_p.t1028 vp_p.t2210 vdd.t789 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2654 vdd.t788 vp_p.t2211 out_p.t1027 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2655 out_p.t82 vp_n.t443 vss.t156 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2656 out_p.t1026 vp_p.t2212 vdd.t787 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2657 out_p.t1025 vp_p.t2213 vdd.t786 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2658 out_p.t1024 vp_p.t2214 vdd.t785 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2659 out_p.t1023 vp_p.t2215 vdd.t784 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2660 out_p.t1022 vp_p.t2216 vdd.t783 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2661 vdd.t782 vp_p.t2217 out_p.t1021 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2662 vdd.t781 vp_p.t2218 out_p.t1020 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2663 vdd.t780 vp_p.t2219 out_p.t1019 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2664 out_p.t1018 vp_p.t2220 vdd.t779 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2665 out_p.t84 vp_n.t444 vss.t155 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2666 out_p.t1017 vp_p.t2221 vdd.t778 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2667 out_p.t1016 vp_p.t2222 vdd.t777 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2668 vdd.t776 vp_p.t2223 out_p.t1015 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2669 vdd.t775 vp_p.t2224 out_p.t1014 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2670 vdd.t774 vp_p.t2225 out_p.t1013 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2671 out_p.t3443 vp_n.t445 vss.t154 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2672 out_p.t85 vp_n.t446 vss.t153 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2673 out_p.t1012 vp_p.t2226 vdd.t773 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2674 vdd.t772 vp_p.t2227 out_p.t1011 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2675 vss.t152 vp_n.t447 out_p.t86 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2676 vdd.t771 vp_p.t2228 out_p.t1010 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2677 vdd.t770 vp_p.t2229 out_p.t1009 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2678 out_p.t3442 vp_n.t448 vss.t151 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2679 out_p.t1008 vp_p.t2230 vdd.t769 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2680 vss.t150 vp_n.t449 out_p.t87 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2681 vdd.t768 vp_p.t2231 out_p.t1007 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2682 out_p.t1006 vp_p.t2232 vdd.t767 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2683 vdd.t766 vp_p.t2233 out_p.t1005 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2684 out_p.t1004 vp_p.t2234 vdd.t765 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2685 vdd.t764 vp_p.t2235 out_p.t1003 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2686 out_p.t89 vp_n.t450 vss.t149 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2687 vss.t148 vp_n.t451 out_p.t3594 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2688 vdd.t763 vp_p.t2236 out_p.t1002 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2689 out_p.t1001 vp_p.t2237 vdd.t762 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2690 out_p.t90 vp_n.t452 vss.t147 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2691 out_p.t1000 vp_p.t2238 vdd.t761 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2692 vss.t146 vp_n.t453 out_p.t202 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2693 out_p.t3593 vp_n.t454 vss.t145 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2694 vdd.t760 vp_p.t2239 out_p.t999 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2695 vdd.t759 vp_p.t2240 out_p.t998 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2696 vdd.t758 vp_p.t2241 out_p.t997 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2697 vdd.t757 vp_p.t2242 out_p.t996 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2698 vss.t144 vp_n.t455 out_p.t92 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2699 vdd.t756 vp_p.t2243 out_p.t995 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2700 vdd.t755 vp_p.t2244 out_p.t994 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2701 out_p.t94 vp_n.t456 vss.t143 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2702 vss.t142 vp_n.t457 out_p.t201 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2703 vdd.t754 vp_p.t2245 out_p.t993 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2704 out_p.t3586 vp_n.t458 vss.t141 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2705 out_p.t992 vp_p.t2246 vdd.t753 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2706 vdd.t752 vp_p.t2247 out_p.t991 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2707 vss.t140 vp_n.t459 out_p.t95 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2708 out_p.t990 vp_p.t2248 vdd.t751 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2709 out_p.t989 vp_p.t2249 vdd.t750 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2710 vss.t139 vp_n.t460 out_p.t200 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2711 out_p.t3585 vp_n.t461 vss.t138 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2712 vss.t137 vp_n.t462 out_p.t97 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2713 vdd.t749 vp_p.t2250 out_p.t988 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2714 out_p.t987 vp_p.t2251 vdd.t748 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2715 vdd.t747 vp_p.t2252 out_p.t986 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2716 vdd.t746 vp_p.t2253 out_p.t985 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2717 out_p.t984 vp_p.t2254 vdd.t745 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2718 out_p.t99 vp_n.t463 vss.t136 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2719 vdd.t744 vp_p.t2255 out_p.t983 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2720 vdd.t743 vp_p.t2256 out_p.t982 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2721 out_p.t981 vp_p.t2257 vdd.t742 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2722 out_p.t980 vp_p.t2258 vdd.t741 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2723 out_p.t199 vp_n.t464 vss.t135 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2724 out_p.t3452 vp_n.t465 vss.t134 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2725 out_p.t979 vp_p.t2259 vdd.t740 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2726 out_p.t978 vp_p.t2260 vdd.t739 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2727 vss.t133 vp_n.t466 out_p.t100 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2728 out_p.t977 vp_p.t2261 vdd.t738 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2729 vdd.t737 vp_p.t2262 out_p.t976 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2730 vss.t132 vp_n.t467 out_p.t198 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2731 out_p.t975 vp_p.t2263 vdd.t736 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2732 out_p.t3451 vp_n.t468 vss.t131 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2733 vdd.t735 vp_p.t2264 out_p.t974 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2734 vdd.t734 vp_p.t2265 out_p.t973 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2735 out_p.t102 vp_n.t469 vss.t130 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2736 out_p.t972 vp_p.t2266 vdd.t733 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2737 vss.t129 vp_n.t470 out_p.t104 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2738 out_p.t971 vp_p.t2267 vdd.t732 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2739 vdd.t731 vp_p.t2268 out_p.t970 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2740 out_p.t969 vp_p.t2269 vdd.t730 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2741 out_p.t968 vp_p.t2270 vdd.t729 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2742 vss.t128 vp_n.t471 out_p.t191 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2743 vdd.t728 vp_p.t2271 out_p.t967 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2744 vdd.t727 vp_p.t2272 out_p.t966 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2745 vdd.t726 vp_p.t2273 out_p.t965 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2746 out_p.t964 vp_p.t2274 vdd.t725 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2747 out_p.t963 vp_p.t2275 vdd.t724 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2748 out_p.t105 vp_n.t472 vss.t127 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2749 vss.t126 vp_n.t473 out_p.t106 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2750 out_p.t197 vp_n.t474 vss.t125 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2751 out_p.t962 vp_p.t2276 vdd.t723 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2752 vdd.t722 vp_p.t2277 out_p.t961 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2753 out_p.t960 vp_p.t2278 vdd.t721 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2754 out_p.t959 vp_p.t2279 vdd.t720 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2755 out_p.t958 vp_p.t2280 vdd.t719 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2756 out_p.t957 vp_p.t2281 vdd.t718 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2757 vdd.t717 vp_p.t2282 out_p.t956 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2758 out_p.t955 vp_p.t2283 vdd.t716 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2759 vdd.t715 vp_p.t2284 out_p.t954 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2760 vss.t124 vp_n.t475 out_p.t190 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2761 out_p.t108 vp_n.t476 vss.t123 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2762 out_p.t953 vp_p.t2285 vdd.t714 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2763 vdd.t713 vp_p.t2286 out_p.t952 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2764 vdd.t712 vp_p.t2287 out_p.t951 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2765 vdd.t711 vp_p.t2288 out_p.t950 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2766 out_p.t949 vp_p.t2289 vdd.t710 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2767 out_p.t948 vp_p.t2290 vdd.t709 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2768 out_p.t110 vp_n.t477 vss.t122 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2769 vdd.t708 vp_p.t2291 out_p.t947 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2770 out_p.t196 vp_n.t478 vss.t121 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2771 vss.t120 vp_n.t479 out_p.t3576 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2772 vdd.t707 vp_p.t2292 out_p.t946 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2773 vss.t119 vp_n.t480 out_p.t111 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2774 out_p.t945 vp_p.t2293 vdd.t706 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2775 out_p.t944 vp_p.t2294 vdd.t705 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2776 vdd.t704 vp_p.t2295 out_p.t943 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2777 vdd.t703 vp_p.t2296 out_p.t942 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2778 vdd.t702 vp_p.t2297 out_p.t941 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2779 vdd.t701 vp_p.t2298 out_p.t940 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2780 vss.t118 vp_n.t481 out_p.t112 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2781 out_p.t195 vp_n.t482 vss.t117 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2782 out_p.t939 vp_p.t2299 vdd.t700 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2783 vss.t116 vp_n.t483 out_p.t3575 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2784 out_p.t938 vp_p.t2300 vdd.t699 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2785 vdd.t698 vp_p.t2301 out_p.t937 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2786 vdd.t697 vp_p.t2302 out_p.t936 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2787 out_p.t113 vp_n.t484 vss.t115 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2788 out_p.t935 vp_p.t2303 vdd.t696 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2789 out_p.t934 vp_p.t2304 vdd.t695 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2790 vdd.t694 vp_p.t2305 out_p.t933 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2791 vdd.t693 vp_p.t2306 out_p.t932 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2792 out_p.t931 vp_p.t2307 vdd.t692 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2793 out_p.t930 vp_p.t2308 vdd.t691 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2794 out_p.t115 vp_n.t485 vss.t114 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2795 vdd.t690 vp_p.t2309 out_p.t929 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2796 vss.t113 vp_n.t486 out_p.t194 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2797 out_p.t928 vp_p.t2310 vdd.t689 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2798 out_p.t927 vp_p.t2311 vdd.t688 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2799 out_p.t926 vp_p.t2312 vdd.t687 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2800 out_p.t3435 vp_n.t487 vss.t112 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2801 out_p.t116 vp_n.t488 vss.t111 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2802 vdd.t686 vp_p.t2313 out_p.t925 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2803 vss.t110 vp_n.t489 out_p.t117 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2804 vdd.t685 vp_p.t2314 out_p.t924 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2805 vdd.t684 vp_p.t2315 out_p.t923 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2806 vdd.t683 vp_p.t2316 out_p.t922 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2807 out_p.t427 vp_n.t490 vss.t109 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2808 vdd.t682 vp_p.t2317 out_p.t921 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2809 out_p.t920 vp_p.t2318 vdd.t681 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2810 out_p.t118 vp_n.t491 vss.t108 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2811 vdd.t680 vp_p.t2319 out_p.t919 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2812 out_p.t918 vp_p.t2320 vdd.t679 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2813 vss.t107 vp_n.t492 out_p.t127 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2814 out_p.t426 vp_n.t493 vss.t106 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2815 out_p.t917 vp_p.t2321 vdd.t678 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2816 out_p.t916 vp_p.t2322 vdd.t677 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2817 vdd.t676 vp_p.t2323 out_p.t915 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2818 out_p.t914 vp_p.t2324 vdd.t675 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2819 vdd.t674 vp_p.t2325 out_p.t913 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2820 vss.t105 vp_n.t494 out_p.t128 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2821 out_p.t912 vp_p.t2326 vdd.t673 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2822 out_p.t119 vp_n.t495 vss.t104 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2823 vss.t103 vp_n.t496 out_p.t3558 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2824 vdd.t672 vp_p.t2327 out_p.t911 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2825 out_p.t910 vp_p.t2328 vdd.t671 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2826 out_p.t909 vp_p.t2329 vdd.t670 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2827 vdd.t669 vp_p.t2330 out_p.t908 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2828 out_p.t907 vp_p.t2331 vdd.t668 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2829 out_p.t906 vp_p.t2332 vdd.t667 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2830 vdd.t666 vp_p.t2333 out_p.t905 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2831 out_p.t904 vp_p.t2334 vdd.t665 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2832 vdd.t664 vp_p.t2335 out_p.t903 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2833 out_p.t902 vp_p.t2336 vdd.t663 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2834 out_p.t901 vp_p.t2337 vdd.t662 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2835 vdd.t661 vp_p.t2338 out_p.t900 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2836 vdd.t660 vp_p.t2339 out_p.t899 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2837 out_p.t120 vp_n.t497 vss.t102 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2838 out_p.t898 vp_p.t2340 vdd.t659 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2839 out_p.t897 vp_p.t2341 vdd.t658 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2840 out_p.t896 vp_p.t2342 vdd.t657 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2841 out_p.t895 vp_p.t2343 vdd.t656 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2842 out_p.t894 vp_p.t2344 vdd.t655 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2843 out_p.t129 vp_n.t498 vss.t101 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2844 out_p.t193 vp_n.t499 vss.t100 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2845 vdd.t654 vp_p.t2345 out_p.t893 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2846 vdd.t653 vp_p.t2346 out_p.t892 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2847 vss.t99 vp_n.t500 out_p.t3557 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2848 out_p.t891 vp_p.t2347 vdd.t652 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2849 vdd.t651 vp_p.t2348 out_p.t890 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2850 out_p.t130 vp_n.t501 vss.t98 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2851 vdd.t650 vp_p.t2349 out_p.t889 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2852 out_p.t888 vp_p.t2350 vdd.t649 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2853 out_p.t887 vp_p.t2351 vdd.t648 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2854 out_p.t886 vp_p.t2352 vdd.t647 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2855 vss.t97 vp_n.t502 out_p.t122 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2856 vdd.t646 vp_p.t2353 out_p.t885 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2857 out_p.t884 vp_p.t2354 vdd.t645 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2858 out_p.t78 vp_n.t503 vss.t96 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2859 out_p.t883 vp_p.t2355 vdd.t644 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2860 out_p.t882 vp_p.t2356 vdd.t643 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2861 vdd.t642 vp_p.t2357 out_p.t881 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2862 vdd.t641 vp_p.t2358 out_p.t880 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2863 out_p.t879 vp_p.t2359 vdd.t640 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2864 vdd.t639 vp_p.t2360 out_p.t878 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2865 out_p.t877 vp_p.t2361 vdd.t638 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2866 vdd.t637 vp_p.t2362 out_p.t876 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2867 out_p.t875 vp_p.t2363 vdd.t636 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2868 vss.t95 vp_n.t504 out_p.t3560 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2869 out_p.t874 vp_p.t2364 vdd.t635 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2870 vdd.t634 vp_p.t2365 out_p.t873 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2871 vdd.t633 vp_p.t2366 out_p.t872 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2872 out_p.t123 vp_n.t505 vss.t94 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2873 out_p.t150 vp_n.t506 vss.t93 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2874 out_p.t871 vp_p.t2367 vdd.t632 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2875 out_p.t192 vp_n.t507 vss.t92 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2876 vss.t91 vp_n.t508 out_p.t3559 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2877 out_p.t151 vp_n.t509 vss.t90 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2878 vdd.t631 vp_p.t2368 out_p.t870 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2879 out_p.t869 vp_p.t2369 vdd.t630 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2880 vss.t89 vp_n.t510 out_p.t141 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2881 vdd.t629 vp_p.t2370 out_p.t868 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2882 out_p.t867 vp_p.t2371 vdd.t628 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2883 out_p.t3429 vp_n.t511 vss.t88 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2884 vss.t87 vp_n.t512 out_p.t142 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2885 out_p.t866 vp_p.t2372 vdd.t627 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2886 vdd.t626 vp_p.t2373 out_p.t865 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2887 out_p.t864 vp_p.t2374 vdd.t625 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2888 out_p.t138 vp_n.t513 vss.t86 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2889 vdd.t624 vp_p.t2375 out_p.t863 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2890 out_p.t862 vp_p.t2376 vdd.t623 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2891 out_p.t32 vp_n.t514 vss.t85 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2892 vdd.t622 vp_p.t2377 out_p.t861 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2893 out_p.t860 vp_p.t2378 vdd.t621 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2894 out_p.t3428 vp_n.t515 vss.t84 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2895 vss.t83 vp_n.t516 out_p.t139 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2896 vdd.t620 vp_p.t2379 out_p.t859 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2897 vss.t82 vp_n.t517 out_p.t132 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2898 out_p.t858 vp_p.t2380 vdd.t619 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2899 out_p.t31 vp_n.t518 vss.t81 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2900 vdd.t618 vp_p.t2381 out_p.t857 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2901 out_p.t856 vp_p.t2382 vdd.t617 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2902 out_p.t3563 vp_n.t519 vss.t80 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2903 vss.t79 vp_n.t520 out_p.t133 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2904 out_p.t855 vp_p.t2383 vdd.t616 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2905 out_p.t854 vp_p.t2384 vdd.t615 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2906 vss.t78 vp_n.t521 out_p.t125 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2907 vdd.t614 vp_p.t2385 out_p.t853 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2908 vdd.t613 vp_p.t2386 out_p.t852 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2909 vdd.t612 vp_p.t2387 out_p.t851 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2910 vdd.t611 vp_p.t2388 out_p.t850 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2911 out_p.t849 vp_p.t2389 vdd.t610 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2912 vdd.t609 vp_p.t2390 out_p.t848 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2913 out_p.t847 vp_p.t2391 vdd.t608 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2914 out_p.t30 vp_n.t522 vss.t77 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2915 vdd.t607 vp_p.t2392 out_p.t846 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2916 out_p.t3562 vp_n.t523 vss.t76 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2917 out_p.t845 vp_p.t2393 vdd.t606 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2918 out_p.t844 vp_p.t2394 vdd.t605 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2919 out_p.t843 vp_p.t2395 vdd.t604 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2920 vss.t75 vp_n.t524 out_p.t126 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2921 out_p.t135 vp_n.t525 vss.t74 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2922 out_p.t842 vp_p.t2396 vdd.t603 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2923 out_p.t841 vp_p.t2397 vdd.t602 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2924 out_p.t840 vp_p.t2398 vdd.t601 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2925 out_p.t839 vp_p.t2399 vdd.t600 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2926 vdd.t599 vp_p.t2400 out_p.t838 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2927 out_p.t837 vp_p.t2401 vdd.t598 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2928 out_p.t29 vp_n.t526 vss.t73 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2929 out_p.t836 vp_p.t2402 vdd.t597 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2930 vss.t72 vp_n.t527 out_p.t3430 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2931 vss.t71 vp_n.t528 out_p.t136 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2932 out_p.t835 vp_p.t2403 vdd.t596 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2933 vdd.t595 vp_p.t2404 out_p.t834 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2934 out_p.t833 vp_p.t2405 vdd.t594 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2935 vss.t70 vp_n.t529 out_p.t145 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2936 out_p.t832 vp_p.t2406 vdd.t593 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2937 out_p.t28 vp_n.t530 vss.t69 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2938 vss.t68 vp_n.t531 out_p.t3432 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2939 vdd.t592 vp_p.t2407 out_p.t831 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2940 out_p.t830 vp_p.t2408 vdd.t591 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2941 out_p.t829 vp_p.t2409 vdd.t590 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2942 vdd.t589 vp_p.t2410 out_p.t828 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2943 vdd.t588 vp_p.t2411 out_p.t827 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2944 vdd.t587 vp_p.t2412 out_p.t826 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2945 vdd.t586 vp_p.t2413 out_p.t825 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2946 vdd.t585 vp_p.t2414 out_p.t824 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2947 out_p.t823 vp_p.t2415 vdd.t584 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2948 out_p.t146 vp_n.t532 vss.t67 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2949 out_p.t822 vp_p.t2416 vdd.t583 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2950 vdd.t582 vp_p.t2417 out_p.t821 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2951 out_p.t820 vp_p.t2418 vdd.t581 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2952 out_p.t819 vp_p.t2419 vdd.t580 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2953 vss.t66 vp_n.t533 out_p.t148 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2954 out_p.t27 vp_n.t534 vss.t65 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2955 vdd.t579 vp_p.t2420 out_p.t818 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2956 vdd.t578 vp_p.t2421 out_p.t817 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2957 vss.t64 vp_n.t535 out_p.t3431 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2958 out_p.t816 vp_p.t2422 vdd.t577 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2959 out_p.t182 vp_n.t536 vss.t63 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2960 out_p.t26 vp_n.t537 vss.t62 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2961 vdd.t576 vp_p.t2423 out_p.t815 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2962 vdd.t575 vp_p.t2424 out_p.t814 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2963 out_p.t813 vp_p.t2425 vdd.t574 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2964 out_p.t3434 vp_n.t538 vss.t61 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2965 out_p.t812 vp_p.t2426 vdd.t573 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2966 vss.t60 vp_n.t539 out_p.t7 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2967 out_p.t811 vp_p.t2427 vdd.t572 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2968 vdd.t571 vp_p.t2428 out_p.t810 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2969 vdd.t570 vp_p.t2429 out_p.t809 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2970 vdd.t569 vp_p.t2430 out_p.t808 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2971 out_p.t9 vp_n.t540 vss.t59 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2972 vss.t58 vp_n.t541 out_p.t25 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2973 vss.t57 vp_n.t542 out_p.t3433 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2974 out_p.t807 vp_p.t2431 vdd.t568 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2975 out_p.t806 vp_p.t2432 vdd.t567 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2976 vdd.t566 vp_p.t2433 out_p.t805 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2977 out_p.t804 vp_p.t2434 vdd.t565 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2978 vdd.t564 vp_p.t2435 out_p.t803 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2979 vdd.t563 vp_p.t2436 out_p.t802 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2980 vdd.t562 vp_p.t2437 out_p.t801 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2981 out_p.t800 vp_p.t2438 vdd.t561 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2982 vdd.t560 vp_p.t2439 out_p.t799 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2983 out_p.t798 vp_p.t2440 vdd.t559 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2984 out_p.t797 vp_p.t2441 vdd.t558 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2985 out_p.t796 vp_p.t2442 vdd.t557 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2986 out_p.t3445 vp_n.t543 vss.t56 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2987 vdd.t556 vp_p.t2443 out_p.t795 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2988 vss.t55 vp_n.t544 out_p.t10 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2989 out_p.t794 vp_p.t2444 vdd.t555 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2990 out_p.t793 vp_p.t2445 vdd.t554 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2991 out_p.t792 vp_p.t2446 vdd.t553 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2992 vss.t54 vp_n.t545 out_p.t24 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2993 vdd.t552 vp_p.t2447 out_p.t791 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2994 out_p.t3574 vp_n.t546 vss.t53 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2995 out_p.t790 vp_p.t2448 vdd.t551 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2996 out_p.t12 vp_n.t547 vss.t52 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2997 out_p.t789 vp_p.t2449 vdd.t550 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2998 out_p.t788 vp_p.t2450 vdd.t549 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2999 out_p.t787 vp_p.t2451 vdd.t548 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3000 out_p.t786 vp_p.t2452 vdd.t547 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3001 vdd.t546 vp_p.t2453 out_p.t785 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3002 out_p.t784 vp_p.t2454 vdd.t545 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3003 vdd.t544 vp_p.t2455 out_p.t783 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3004 out_p.t782 vp_p.t2456 vdd.t543 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3005 vdd.t542 vp_p.t2457 out_p.t781 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3006 out_p.t780 vp_p.t2458 vdd.t541 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3007 out_p.t779 vp_p.t2459 vdd.t540 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3008 vdd.t539 vp_p.t2460 out_p.t778 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3009 vdd.t538 vp_p.t2461 out_p.t777 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3010 vdd.t537 vp_p.t2462 out_p.t776 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3011 vdd.t536 vp_p.t2463 out_p.t775 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3012 vdd.t535 vp_p.t2464 out_p.t774 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3013 out_p.t773 vp_p.t2465 vdd.t534 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3014 out_p.t772 vp_p.t2466 vdd.t533 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3015 out_p.t14 vp_n.t548 vss.t51 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3016 vdd.t532 vp_p.t2467 out_p.t771 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3017 vdd.t531 vp_p.t2468 out_p.t770 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3018 vdd.t530 vp_p.t2469 out_p.t769 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3019 out_p.t768 vp_p.t2470 vdd.t529 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3020 out_p.t767 vp_p.t2471 vdd.t528 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3021 vdd.t527 vp_p.t2472 out_p.t766 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3022 out_p.t765 vp_p.t2473 vdd.t526 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3023 vdd.t525 vp_p.t2474 out_p.t764 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3024 vss.t50 vp_n.t549 out_p.t23 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3025 out_p.t3573 vp_n.t550 vss.t49 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3026 vss.t48 vp_n.t551 out_p.t15 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3027 out_p.t16 vp_n.t552 vss.t47 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3028 out_p.t763 vp_p.t2475 vdd.t524 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3029 out_p.t22 vp_n.t553 vss.t46 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3030 vdd.t523 vp_p.t2476 out_p.t762 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3031 vss.t45 vp_n.t554 out_p.t3587 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3032 out_p.t17 vp_n.t555 vss.t44 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3033 vdd.t522 vp_p.t2477 out_p.t761 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3034 out_p.t760 vp_p.t2478 vdd.t521 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3035 vdd.t520 vp_p.t2479 out_p.t759 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3036 vdd.t519 vp_p.t2480 out_p.t758 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3037 vdd.t518 vp_p.t2481 out_p.t757 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3038 vdd.t517 vp_p.t2482 out_p.t756 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3039 vss.t43 vp_n.t556 out_p.t18 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3040 vdd.t516 vp_p.t2483 out_p.t755 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3041 vdd.t515 vp_p.t2484 out_p.t754 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3042 vdd.t514 vp_p.t2485 out_p.t753 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3043 vdd.t513 vp_p.t2486 out_p.t752 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3044 vdd.t512 vp_p.t2487 out_p.t751 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3045 out_p.t750 vp_p.t2488 vdd.t511 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3046 out_p.t749 vp_p.t2489 vdd.t510 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3047 vdd.t509 vp_p.t2490 out_p.t748 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3048 vdd.t508 vp_p.t2491 out_p.t747 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3049 vdd.t507 vp_p.t2492 out_p.t746 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3050 out_p.t21 vp_n.t557 vss.t42 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3051 out_p.t745 vp_p.t2493 vdd.t506 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3052 vss.t41 vp_n.t558 out_p.t19 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3053 out_p.t744 vp_p.t2494 vdd.t505 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3054 out_p.t743 vp_p.t2495 vdd.t504 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3055 out_p.t742 vp_p.t2496 vdd.t503 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3056 out_p.t741 vp_p.t2497 vdd.t502 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3057 vdd.t501 vp_p.t2498 out_p.t740 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3058 vss.t40 vp_n.t559 out_p.t20 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3059 out_p.t739 vp_p.t2499 vdd.t500 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3060 vdd.t499 vp_p.t2500 out_p.t738 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3061 vdd.t498 vp_p.t2501 out_p.t737 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3062 out_p.t424 vp_n.t560 vss.t39 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3063 vss.t38 vp_n.t561 out_p.t143 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3064 vdd.t497 vp_p.t2502 out_p.t736 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3065 out_p.t735 vp_p.t2503 vdd.t496 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3066 out_p.t3471 vp_n.t562 vss.t37 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3067 vdd.t495 vp_p.t2504 out_p.t734 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3068 vdd.t494 vp_p.t2505 out_p.t733 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3069 out_p.t732 vp_p.t2506 vdd.t493 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3070 out_p.t731 vp_p.t2507 vdd.t492 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3071 out_p.t730 vp_p.t2508 vdd.t491 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3072 vdd.t490 vp_p.t2509 out_p.t729 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3073 out_p.t728 vp_p.t2510 vdd.t489 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3074 vdd.t488 vp_p.t2511 out_p.t727 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3075 vdd.t487 vp_p.t2512 out_p.t726 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3076 vdd.t486 vp_p.t2513 out_p.t725 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3077 vdd.t485 vp_p.t2514 out_p.t724 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3078 out_p.t723 vp_p.t2515 vdd.t484 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3079 out_p.t722 vp_p.t2516 vdd.t483 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3080 out_p.t3577 vp_n.t563 vss.t36 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3081 out_p.t721 vp_p.t2517 vdd.t482 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3082 vdd.t481 vp_p.t2518 out_p.t720 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3083 vdd.t480 vp_p.t2519 out_p.t719 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3084 out_p.t718 vp_p.t2520 vdd.t479 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3085 vdd.t478 vp_p.t2521 out_p.t717 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3086 vdd.t477 vp_p.t2522 out_p.t716 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3087 out_p.t715 vp_p.t2523 vdd.t476 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3088 out_p.t714 vp_p.t2524 vdd.t475 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3089 vss.t35 vp_n.t564 out_p.t3536 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3090 vdd.t474 vp_p.t2525 out_p.t713 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3091 out_p.t712 vp_p.t2526 vdd.t473 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3092 vdd.t472 vp_p.t2527 out_p.t711 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3093 vss.t34 vp_n.t565 out_p.t4 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3094 vdd.t471 vp_p.t2528 out_p.t710 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3095 vdd.t470 vp_p.t2529 out_p.t709 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3096 out_p.t708 vp_p.t2530 vdd.t469 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3097 out_p.t707 vp_p.t2531 vdd.t468 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3098 vdd.t467 vp_p.t2532 out_p.t706 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3099 vdd.t466 vp_p.t2533 out_p.t705 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3100 vdd.t465 vp_p.t2534 out_p.t704 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3101 out_p.t3579 vp_n.t566 vss.t33 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3102 vdd.t464 vp_p.t2535 out_p.t703 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3103 out_p.t3551 vp_n.t567 vss.t32 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3104 out_p.t702 vp_p.t2536 vdd.t463 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3105 vss.t31 vp_n.t568 out_p.t423 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3106 vdd.t462 vp_p.t2537 out_p.t701 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3107 vdd.t461 vp_p.t2538 out_p.t700 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3108 vdd.t460 vp_p.t2539 out_p.t699 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3109 vss.t30 vp_n.t569 out_p.t425 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3110 vdd.t459 vp_p.t2540 out_p.t698 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3111 vdd.t458 vp_p.t2541 out_p.t697 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3112 vdd.t457 vp_p.t2542 out_p.t696 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3113 out_p.t695 vp_p.t2543 vdd.t456 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3114 out_p.t694 vp_p.t2544 vdd.t455 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3115 vss.t29 vp_n.t570 out_p.t3465 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3116 out_p.t3511 vp_n.t571 vss.t28 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3117 vdd.t454 vp_p.t2545 out_p.t693 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3118 vdd.t453 vp_p.t2546 out_p.t692 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3119 vdd.t452 vp_p.t2547 out_p.t691 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3120 vdd.t451 vp_p.t2548 out_p.t690 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3121 out_p.t689 vp_p.t2549 vdd.t450 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3122 out_p.t3450 vp_n.t572 vss.t27 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3123 vss.t26 vp_n.t573 out_p.t305 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3124 vss.t25 vp_n.t574 out_p.t278 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3125 out_p.t688 vp_p.t2550 vdd.t449 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3126 vdd.t448 vp_p.t2551 out_p.t687 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3127 out_p.t316 vp_n.t575 vss.t24 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3128 out_p.t686 vp_p.t2552 vdd.t447 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3129 out_p.t3469 vp_n.t576 vss.t23 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3130 vss.t22 vp_n.t577 out_p.t3470 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3131 vdd.t446 vp_p.t2553 out_p.t685 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3132 vdd.t445 vp_p.t2554 out_p.t684 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3133 out_p.t683 vp_p.t2555 vdd.t444 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3134 vdd.t443 vp_p.t2556 out_p.t682 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3135 vdd.t442 vp_p.t2557 out_p.t681 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3136 out_p.t680 vp_p.t2558 vdd.t441 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3137 out_p.t679 vp_p.t2559 vdd.t440 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3138 vdd.t439 vp_p.t2560 out_p.t678 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3139 vss.t21 vp_n.t578 out_p.t3466 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3140 out_p.t677 vp_p.t2561 vdd.t438 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3141 vdd.t437 vp_p.t2562 out_p.t676 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3142 out_p.t675 vp_p.t2563 vdd.t436 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3143 out_p.t674 vp_p.t2564 vdd.t435 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3144 out_p.t673 vp_p.t2565 vdd.t434 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3145 out_p.t672 vp_p.t2566 vdd.t433 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3146 vss.t20 vp_n.t579 out_p.t3501 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3147 out_p.t3502 vp_n.t580 vss.t19 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3148 out_p.t671 vp_p.t2567 vdd.t432 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3149 vdd.t431 vp_p.t2568 out_p.t670 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3150 vdd.t430 vp_p.t2569 out_p.t669 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3151 out_p.t668 vp_p.t2570 vdd.t429 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3152 out_p.t667 vp_p.t2571 vdd.t428 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3153 vdd.t427 vp_p.t2572 out_p.t666 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3154 out_p.t665 vp_p.t2573 vdd.t426 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3155 vdd.t425 vp_p.t2574 out_p.t664 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3156 out_p.t663 vp_p.t2575 vdd.t424 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3157 vdd.t423 vp_p.t2576 out_p.t662 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3158 out_p.t3518 vp_n.t581 vss.t18 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3159 vdd.t422 vp_p.t2577 out_p.t661 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3160 vdd.t421 vp_p.t2578 out_p.t660 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3161 out_p.t659 vp_p.t2579 vdd.t420 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3162 vdd.t419 vp_p.t2580 out_p.t658 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3163 out_p.t657 vp_p.t2581 vdd.t418 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3164 out_p.t656 vp_p.t2582 vdd.t417 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3165 out_p.t655 vp_p.t2583 vdd.t416 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3166 vdd.t415 vp_p.t2584 out_p.t654 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3167 out_p.t3513 vp_n.t582 vss.t17 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3168 vss.t16 vp_n.t583 out_p.t3507 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3169 vdd.t414 vp_p.t2585 out_p.t653 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3170 vdd.t413 vp_p.t2586 out_p.t652 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3171 vdd.t412 vp_p.t2587 out_p.t651 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3172 vdd.t411 vp_p.t2588 out_p.t650 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3173 vdd.t410 vp_p.t2589 out_p.t649 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3174 vdd.t409 vp_p.t2590 out_p.t648 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3175 vdd.t408 vp_p.t2591 out_p.t647 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3176 out_p.t319 vp_n.t584 vss.t15 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3177 out_p.t646 vp_p.t2592 vdd.t407 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3178 vdd.t406 vp_p.t2593 out_p.t645 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3179 vdd.t405 vp_p.t2594 out_p.t644 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3180 vss.t14 vp_n.t585 out_p.t318 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3181 vss.t13 vp_n.t586 out_p.t3489 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3182 out_p.t643 vp_p.t2595 vdd.t404 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3183 vdd.t403 vp_p.t2596 out_p.t642 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3184 out_p.t641 vp_p.t2597 vdd.t402 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3185 out_p.t317 vp_n.t587 vss.t12 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3186 vdd.t401 vp_p.t2598 out_p.t640 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3187 vdd.t400 vp_p.t2599 out_p.t639 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3188 vdd.t399 vp_p.t2600 out_p.t638 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3189 out_p.t637 vp_p.t2601 vdd.t398 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3190 out_p.t314 vp_n.t588 vss.t11 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3191 vdd.t397 vp_p.t2602 out_p.t636 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3192 out_p.t635 vp_p.t2603 vdd.t396 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3193 vdd.t395 vp_p.t2604 out_p.t634 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3194 vdd.t394 vp_p.t2605 out_p.t633 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3195 vdd.t393 vp_p.t2606 out_p.t632 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3196 out_p.t631 vp_p.t2607 vdd.t392 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3197 vss.t10 vp_n.t589 out_p.t315 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3198 out_p.t630 vp_p.t2608 vdd.t391 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3199 vdd.t390 vp_p.t2609 out_p.t629 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3200 vdd.t389 vp_p.t2610 out_p.t628 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3201 vss.t9 vp_n.t590 out_p.t298 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3202 out_p.t627 vp_p.t2611 vdd.t388 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3203 vdd.t387 vp_p.t2612 out_p.t626 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3204 out_p.t3532 vp_n.t591 vss.t8 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3205 out_p.t625 vp_p.t2613 vdd.t386 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3206 vdd.t385 vp_p.t2614 out_p.t624 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3207 vdd.t384 vp_p.t2615 out_p.t623 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3208 out_p.t622 vp_p.t2616 vdd.t383 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3209 out_p.t621 vp_p.t2617 vdd.t382 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3210 vss.t7 vp_n.t592 out_p.t225 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3211 out_p.t620 vp_p.t2618 vdd.t381 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3212 out_p.t619 vp_p.t2619 vdd.t380 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3213 out_p.t618 vp_p.t2620 vdd.t379 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3214 out_p.t617 vp_p.t2621 vdd.t378 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3215 vdd.t377 vp_p.t2622 out_p.t616 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3216 out_p.t615 vp_p.t2623 vdd.t376 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3217 out_p.t614 vp_p.t2624 vdd.t375 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3218 out_p.t613 vp_p.t2625 vdd.t374 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3219 out_p.t612 vp_p.t2626 vdd.t373 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3220 vdd.t372 vp_p.t2627 out_p.t611 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3221 vdd.t371 vp_p.t2628 out_p.t610 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3222 vdd.t370 vp_p.t2629 out_p.t609 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3223 vdd.t369 vp_p.t2630 out_p.t608 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3224 out_p.t607 vp_p.t2631 vdd.t368 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3225 out_p.t606 vp_p.t2632 vdd.t367 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3226 out_p.t605 vp_p.t2633 vdd.t366 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3227 vdd.t365 vp_p.t2634 out_p.t604 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3228 vdd.t364 vp_p.t2635 out_p.t603 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3229 out_p.t602 vp_p.t2636 vdd.t363 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3230 vdd.t362 vp_p.t2637 out_p.t601 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3231 out_p.t600 vp_p.t2638 vdd.t361 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3232 vdd.t360 vp_p.t2639 out_p.t599 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3233 vdd.t359 vp_p.t2640 out_p.t598 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3234 out_p.t597 vp_p.t2641 vdd.t358 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3235 vdd.t357 vp_p.t2642 out_p.t596 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3236 out_p.t595 vp_p.t2643 vdd.t356 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3237 vdd.t355 vp_p.t2644 out_p.t594 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3238 out_p.t593 vp_p.t2645 vdd.t354 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3239 vdd.t353 vp_p.t2646 out_p.t592 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3240 vdd.t352 vp_p.t2647 out_p.t591 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3241 vss.t6 vp_n.t593 out_p.t234 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3242 out_p.t590 vp_p.t2648 vdd.t351 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3243 out_p.t589 vp_p.t2649 vdd.t350 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3244 vss.t5 vp_n.t594 out_p.t241 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3245 vdd.t349 vp_p.t2650 out_p.t588 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3246 out_p.t587 vp_p.t2651 vdd.t348 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3247 out_p.t586 vp_p.t2652 vdd.t347 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3248 vdd.t346 vp_p.t2653 out_p.t585 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3249 vdd.t345 vp_p.t2654 out_p.t584 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3250 out_p.t583 vp_p.t2655 vdd.t344 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3251 out_p.t582 vp_p.t2656 vdd.t343 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3252 out_p.t581 vp_p.t2657 vdd.t342 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3253 vdd.t341 vp_p.t2658 out_p.t580 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3254 vdd.t340 vp_p.t2659 out_p.t579 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3255 vdd.t339 vp_p.t2660 out_p.t578 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3256 vdd.t338 vp_p.t2661 out_p.t577 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3257 vss.t4 vp_n.t595 out_p.t245 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3258 out_p.t576 vp_p.t2662 vdd.t337 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3259 out_p.t575 vp_p.t2663 vdd.t336 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3260 out_p.t574 vp_p.t2664 vdd.t335 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3261 out_p.t573 vp_p.t2665 vdd.t334 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3262 vdd.t333 vp_p.t2666 out_p.t572 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3263 out_p.t248 vp_n.t596 vss.t3 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3264 out_p.t571 vp_p.t2667 vdd.t332 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3265 out_p.t570 vp_p.t2668 vdd.t331 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3266 vdd.t330 vp_p.t2669 out_p.t569 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3267 vdd.t329 vp_p.t2670 out_p.t568 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3268 vss.t2 vp_n.t597 out_p.t252 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3269 vdd.t328 vp_p.t2671 out_p.t567 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3270 vdd.t327 vp_p.t2672 out_p.t566 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3271 out_p.t565 vp_p.t2673 vdd.t326 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3272 vdd.t325 vp_p.t2674 out_p.t564 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3273 vdd.t324 vp_p.t2675 out_p.t563 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3274 vdd.t323 vp_p.t2676 out_p.t562 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3275 out_p.t561 vp_p.t2677 vdd.t322 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3276 out_p.t560 vp_p.t2678 vdd.t321 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3277 vdd.t320 vp_p.t2679 out_p.t559 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3278 vdd.t319 vp_p.t2680 out_p.t558 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3279 out_p.t557 vp_p.t2681 vdd.t318 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3280 vdd.t317 vp_p.t2682 out_p.t556 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3281 vdd.t316 vp_p.t2683 out_p.t555 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3282 vdd.t315 vp_p.t2684 out_p.t554 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3283 out_p.t553 vp_p.t2685 vdd.t314 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3284 vdd.t313 vp_p.t2686 out_p.t552 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3285 out_p.t551 vp_p.t2687 vdd.t312 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3286 vdd.t311 vp_p.t2688 out_p.t550 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3287 vdd.t310 vp_p.t2689 out_p.t549 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3288 vdd.t309 vp_p.t2690 out_p.t548 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3289 out_p.t547 vp_p.t2691 vdd.t308 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3290 vdd.t307 vp_p.t2692 out_p.t546 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3291 out_p.t545 vp_p.t2693 vdd.t306 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3292 vdd.t305 vp_p.t2694 out_p.t544 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3293 out_p.t543 vp_p.t2695 vdd.t304 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3294 vdd.t303 vp_p.t2696 out_p.t542 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3295 out_p.t541 vp_p.t2697 vdd.t302 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3296 out_p.t540 vp_p.t2698 vdd.t301 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3297 vdd.t300 vp_p.t2699 out_p.t539 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3298 vdd.t299 vp_p.t2700 out_p.t538 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3299 out_p.t537 vp_p.t2701 vdd.t298 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3300 out_p.t536 vp_p.t2702 vdd.t297 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3301 vdd.t296 vp_p.t2703 out_p.t535 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3302 vdd.t295 vp_p.t2704 out_p.t534 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3303 out_p.t533 vp_p.t2705 vdd.t294 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3304 out_p.t532 vp_p.t2706 vdd.t293 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3305 out_p.t531 vp_p.t2707 vdd.t292 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3306 vdd.t291 vp_p.t2708 out_p.t530 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3307 out_p.t529 vp_p.t2709 vdd.t290 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3308 vdd.t289 vp_p.t2710 out_p.t528 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3309 vdd.t288 vp_p.t2711 out_p.t527 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3310 out_p.t526 vp_p.t2712 vdd.t287 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3311 out_p.t525 vp_p.t2713 vdd.t286 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3312 out_p.t524 vp_p.t2714 vdd.t285 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3313 out_p.t254 vp_n.t598 vss.t1 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3314 vdd.t284 vp_p.t2715 out_p.t523 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3315 vdd.t283 vp_p.t2716 out_p.t522 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3316 vdd.t282 vp_p.t2717 out_p.t521 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3317 vdd.t281 vp_p.t2718 out_p.t520 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3318 vdd.t280 vp_p.t2719 out_p.t519 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3319 vdd.t279 vp_p.t2720 out_p.t518 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3320 vss.t0 vp_n.t599 out_p.t259 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3321 vdd.t278 vp_p.t2721 out_p.t517 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3322 vdd.t277 vp_p.t2722 out_p.t516 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3323 vdd.t276 vp_p.t2723 out_p.t515 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3324 vdd.t275 vp_p.t2724 out_p.t514 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3325 vdd.t274 vp_p.t2725 out_p.t513 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3326 out_p.t512 vp_p.t2726 vdd.t273 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3327 out_p.t511 vp_p.t2727 vdd.t272 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3328 out_p.t510 vp_p.t2728 vdd.t271 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3329 vdd.t270 vp_p.t2729 out_p.t509 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3330 vdd.t269 vp_p.t2730 out_p.t508 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3331 out_p.t507 vp_p.t2731 vdd.t268 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3332 vdd.t267 vp_p.t2732 out_p.t506 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3333 out_p.t505 vp_p.t2733 vdd.t266 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3334 out_p.t504 vp_p.t2734 vdd.t265 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3335 vdd.t264 vp_p.t2735 out_p.t503 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3336 out_p.t502 vp_p.t2736 vdd.t263 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3337 vdd.t262 vp_p.t2737 out_p.t501 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3338 out_p.t500 vp_p.t2738 vdd.t261 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3339 out_p.t499 vp_p.t2739 vdd.t260 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3340 vdd.t259 vp_p.t2740 out_p.t498 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3341 out_p.t497 vp_p.t2741 vdd.t258 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3342 out_p.t496 vp_p.t2742 vdd.t257 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3343 out_p.t495 vp_p.t2743 vdd.t256 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3344 out_p.t494 vp_p.t2744 vdd.t255 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3345 vdd.t254 vp_p.t2745 out_p.t493 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3346 out_p.t492 vp_p.t2746 vdd.t253 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3347 out_p.t491 vp_p.t2747 vdd.t252 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3348 vdd.t251 vp_p.t2748 out_p.t490 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3349 out_p.t489 vp_p.t2749 vdd.t250 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3350 vdd.t249 vp_p.t2750 out_p.t488 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3351 vdd.t248 vp_p.t2751 out_p.t487 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3352 out_p.t486 vp_p.t2752 vdd.t247 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3353 vdd.t246 vp_p.t2753 out_p.t485 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3354 vdd.t245 vp_p.t2754 out_p.t484 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3355 vdd.t244 vp_p.t2755 out_p.t483 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3356 vdd.t243 vp_p.t2756 out_p.t482 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3357 out_p.t481 vp_p.t2757 vdd.t242 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3358 out_p.t480 vp_p.t2758 vdd.t241 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3359 out_p.t479 vp_p.t2759 vdd.t240 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3360 vdd.t239 vp_p.t2760 out_p.t478 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3361 out_p.t477 vp_p.t2761 vdd.t238 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3362 vdd.t237 vp_p.t2762 out_p.t476 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3363 vdd.t236 vp_p.t2763 out_p.t475 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3364 vdd.t235 vp_p.t2764 out_p.t474 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3365 out_p.t473 vp_p.t2765 vdd.t234 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3366 vdd.t233 vp_p.t2766 out_p.t472 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3367 out_p.t471 vp_p.t2767 vdd.t232 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3368 vdd.t231 vp_p.t2768 out_p.t470 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3369 out_p.t469 vp_p.t2769 vdd.t230 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3370 vdd.t229 vp_p.t2770 out_p.t468 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3371 vdd.t228 vp_p.t2771 out_p.t467 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3372 vdd.t227 vp_p.t2772 out_p.t466 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3373 vdd.t226 vp_p.t2773 out_p.t465 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3374 vdd.t225 vp_p.t2774 out_p.t464 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3375 vdd.t224 vp_p.t2775 out_p.t463 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3376 out_p.t462 vp_p.t2776 vdd.t223 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3377 out_p.t461 vp_p.t2777 vdd.t222 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3378 vdd.t221 vp_p.t2778 out_p.t460 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3379 vdd.t220 vp_p.t2779 out_p.t459 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3380 out_p.t458 vp_p.t2780 vdd.t219 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3381 vdd.t218 vp_p.t2781 out_p.t2501 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3382 vdd.t217 vp_p.t2782 out_p.t2500 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3383 vdd.t216 vp_p.t2783 out_p.t2499 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3384 out_p.t2498 vp_p.t2784 vdd.t215 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3385 out_p.t2497 vp_p.t2785 vdd.t214 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3386 vdd.t213 vp_p.t2786 out_p.t2496 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3387 out_p.t1346 vp_p.t2787 vdd.t212 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3388 vdd.t211 vp_p.t2788 out_p.t1345 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3389 out_p.t1344 vp_p.t2789 vdd.t210 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3390 vdd.t209 vp_p.t2790 out_p.t1343 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3391 out_p.t1342 vp_p.t2791 vdd.t208 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3392 vdd.t207 vp_p.t2792 out_p.t1341 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3393 vdd.t206 vp_p.t2793 out_p.t1351 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3394 out_p.t1350 vp_p.t2794 vdd.t205 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3395 out_p.t1349 vp_p.t2795 vdd.t204 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3396 vdd.t203 vp_p.t2796 out_p.t1348 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3397 vdd.t202 vp_p.t2797 out_p.t1267 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3398 out_p.t1266 vp_p.t2798 vdd.t201 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3399 out_p.t1265 vp_p.t2799 vdd.t200 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3400 vdd.t199 vp_p.t2800 out_p.t1264 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3401 out_p.t2495 vp_p.t2801 vdd.t198 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3402 out_p.t2494 vp_p.t2802 vdd.t197 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3403 vdd.t196 vp_p.t2803 out_p.t2493 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3404 out_p.t2491 vp_p.t2804 vdd.t195 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3405 out_p.t2490 vp_p.t2805 vdd.t194 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3406 vdd.t193 vp_p.t2806 out_p.t2489 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3407 vdd.t192 vp_p.t2807 out_p.t2454 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3408 out_p.t2453 vp_p.t2808 vdd.t191 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3409 out_p.t2452 vp_p.t2809 vdd.t190 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3410 out_p.t1256 vp_p.t2810 vdd.t189 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3411 out_p.t1255 vp_p.t2811 vdd.t188 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3412 vdd.t187 vp_p.t2812 out_p.t1318 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3413 vdd.t186 vp_p.t2813 out_p.t1317 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3414 out_p.t1313 vp_p.t2814 vdd.t185 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3415 out_p.t1312 vp_p.t2815 vdd.t184 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3416 out_p.t1305 vp_p.t2816 vdd.t183 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3417 vdd.t182 vp_p.t2817 out_p.t1304 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3418 vdd.t181 vp_p.t2818 out_p.t2449 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3419 out_p.t2448 vp_p.t2819 vdd.t180 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3420 out_p.t2483 vp_p.t2820 vdd.t179 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3421 vdd.t178 vp_p.t2821 out_p.t2482 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3422 vdd.t177 vp_p.t2822 out_p.t2481 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3423 vdd.t176 vp_p.t2823 out_p.t2480 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3424 vdd.t175 vp_p.t2824 out_p.t2479 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3425 out_p.t2478 vp_p.t2825 vdd.t174 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3426 out_p.t2517 vp_p.t2826 vdd.t173 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3427 out_p.t2516 vp_p.t2827 vdd.t172 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3428 out_p.t1253 vp_p.t2828 vdd.t171 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3429 out_p.t1252 vp_p.t2829 vdd.t170 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3430 vdd.t169 vp_p.t2830 out_p.t1339 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3431 vdd.t168 vp_p.t2831 out_p.t1338 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3432 out_p.t1331 vp_p.t2832 vdd.t167 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3433 out_p.t1330 vp_p.t2833 vdd.t166 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3434 out_p.t1356 vp_p.t2834 vdd.t165 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3435 vdd.t164 vp_p.t2835 out_p.t1355 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3436 vdd.t163 vp_p.t2836 out_p.t1353 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3437 out_p.t1352 vp_p.t2837 vdd.t162 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3438 out_p.t1359 vp_p.t2838 vdd.t161 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3439 out_p.t1358 vp_p.t2839 vdd.t160 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3440 vdd.t159 vp_p.t2840 out_p.t2487 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3441 vdd.t158 vp_p.t2841 out_p.t2486 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3442 vdd.t157 vp_p.t2842 out_p.t1242 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3443 out_p.t1241 vp_p.t2843 vdd.t156 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3444 vdd.t155 vp_p.t2844 out_p.t1235 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3445 vdd.t154 vp_p.t2845 out_p.t1234 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3446 vdd.t153 vp_p.t2846 out_p.t1263 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3447 vdd.t152 vp_p.t2847 out_p.t1262 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3448 vdd.t151 vp_p.t2848 out_p.t1246 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3449 out_p.t1245 vp_p.t2849 vdd.t150 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3450 vdd.t149 vp_p.t2850 out_p.t1244 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3451 out_p.t1243 vp_p.t2851 vdd.t148 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3452 vdd.t147 vp_p.t2852 out_p.t1269 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3453 vdd.t146 vp_p.t2853 out_p.t1268 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3454 out_p.t1334 vp_p.t2854 vdd.t145 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3455 vdd.t144 vp_p.t2855 out_p.t1333 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3456 vdd.t143 vp_p.t2856 out_p.t1274 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3457 out_p.t1273 vp_p.t2857 vdd.t142 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3458 vdd.t141 vp_p.t2858 out_p.t1328 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3459 vdd.t140 vp_p.t2859 out_p.t1327 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3460 vdd.t139 vp_p.t2860 out_p.t1323 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3461 out_p.t1322 vp_p.t2861 vdd.t138 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3462 vdd.t137 vp_p.t2862 out_p.t1282 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3463 vdd.t136 vp_p.t2863 out_p.t1281 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3464 out_p.t1285 vp_p.t2864 vdd.t135 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3465 out_p.t1284 vp_p.t2865 vdd.t134 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3466 out_p.t1289 vp_p.t2866 vdd.t133 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3467 out_p.t1288 vp_p.t2867 vdd.t132 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3468 out_p.t1293 vp_p.t2868 vdd.t131 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3469 out_p.t1292 vp_p.t2869 vdd.t130 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3470 out_p.t2515 vp_p.t2870 vdd.t129 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3471 vdd.t128 vp_p.t2871 out_p.t1237 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3472 out_p.t1257 vp_p.t2872 vdd.t127 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3473 out_p.t1251 vp_p.t2873 vdd.t126 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3474 vdd.t125 vp_p.t2874 out_p.t1336 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3475 out_p.t1320 vp_p.t2875 vdd.t124 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3476 out_p.t1319 vp_p.t2876 vdd.t123 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3477 out_p.t1315 vp_p.t2877 vdd.t122 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3478 out_p.t1310 vp_p.t2878 vdd.t121 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3479 vdd.t120 vp_p.t2879 out_p.t1307 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3480 out_p.t1308 vp_p.t2880 vdd.t119 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3481 out_p.t1306 vp_p.t2881 vdd.t118 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3482 vdd.t117 vp_p.t2882 out_p.t1302 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3483 vdd.t116 vp_p.t2883 out_p.t1299 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3484 out_p.t2476 vp_p.t2884 vdd.t115 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3485 vdd.t114 vp_p.t2885 out_p.t1226 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3486 out_p.t2514 vp_p.t2886 vdd.t113 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3487 vdd.t112 vp_p.t2887 out_p.t2513 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3488 out_p.t2484 vp_p.t2888 vdd.t111 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3489 vdd.t110 vp_p.t2889 out_p.t2477 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3490 out_p.t2441 vp_p.t2890 vdd.t109 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3491 out_p.t1230 vp_p.t2891 vdd.t108 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3492 vdd.t107 vp_p.t2892 out_p.t1239 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3493 vdd.t106 vp_p.t2893 out_p.t1232 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3494 out_p.t1258 vp_p.t2894 vdd.t105 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3495 out_p.t1260 vp_p.t2895 vdd.t104 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3496 vdd.t103 vp_p.t2896 out_p.t1248 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3497 vdd.t102 vp_p.t2897 out_p.t1337 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3498 vdd.t101 vp_p.t2898 out_p.t1272 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3499 out_p.t1276 vp_p.t2899 vdd.t100 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3500 vdd.t99 vp_p.t2900 out_p.t1277 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3501 vdd.t98 vp_p.t2901 out_p.t1280 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3502 vdd.t97 vp_p.t2902 out_p.t1314 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3503 out_p.t1283 vp_p.t2903 vdd.t96 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3504 out_p.t1287 vp_p.t2904 vdd.t95 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3505 vdd.t94 vp_p.t2905 out_p.t1291 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3506 vdd.t93 vp_p.t2906 out_p.t1295 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3507 vdd.t92 vp_p.t2907 out_p.t1227 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3508 vdd.t91 vp_p.t2908 out_p.t2475 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3509 vdd.t90 vp_p.t2909 out_p.t2512 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3510 out_p.t2381 vp_p.t2910 vdd.t89 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3511 out_p.t2455 vp_p.t2911 vdd.t88 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3512 vdd.t87 vp_p.t2912 out_p.t439 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3513 vdd.t86 vp_p.t2913 out_p.t1240 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3514 out_p.t1236 vp_p.t2914 vdd.t85 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3515 out_p.t1261 vp_p.t2915 vdd.t84 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3516 vdd.t83 vp_p.t2916 out_p.t1247 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3517 out_p.t1254 vp_p.t2917 vdd.t82 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3518 vdd.t81 vp_p.t2918 out_p.t1340 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3519 vdd.t80 vp_p.t2919 out_p.t1271 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3520 out_p.t1332 vp_p.t2920 vdd.t79 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3521 out_p.t1335 vp_p.t2921 vdd.t78 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3522 vdd.t77 vp_p.t2922 out_p.t1275 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3523 vdd.t76 vp_p.t2923 out_p.t1326 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3524 out_p.t1324 vp_p.t2924 vdd.t75 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3525 vdd.t74 vp_p.t2925 out_p.t1321 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3526 out_p.t1279 vp_p.t2926 vdd.t73 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3527 out_p.t1316 vp_p.t2927 vdd.t72 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3528 out_p.t1311 vp_p.t2928 vdd.t71 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3529 vdd.t70 vp_p.t2929 out_p.t1286 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3530 out_p.t1259 vp_p.t2930 vdd.t69 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3531 out_p.t1290 vp_p.t2931 vdd.t68 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3532 out_p.t1303 vp_p.t2932 vdd.t67 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3533 vdd.t66 vp_p.t2933 out_p.t1294 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3534 vdd.t65 vp_p.t2934 out_p.t1296 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3535 out_p.t1297 vp_p.t2935 vdd.t64 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3536 out_p.t1298 vp_p.t2936 vdd.t63 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3537 vdd.t62 vp_p.t2937 out_p.t2492 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3538 out_p.t2488 vp_p.t2938 vdd.t61 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3539 vdd.t60 vp_p.t2939 out_p.t2427 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3540 vdd.t59 vp_p.t2940 out_p.t2485 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3541 vdd.t58 vp_p.t2941 out_p.t2403 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3542 vdd.t57 vp_p.t2942 out_p.t2408 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3543 vdd.t56 vp_p.t2943 out_p.t2445 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3544 vdd.t55 vp_p.t2944 out_p.t2474 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3545 out_p.t2442 vp_p.t2945 vdd.t54 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3546 vdd.t53 vp_p.t2946 out_p.t2438 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3547 vdd.t52 vp_p.t2947 out_p.t2404 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3548 out_p.t2432 vp_p.t2948 vdd.t51 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3549 out_p.t2437 vp_p.t2949 vdd.t50 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3550 out_p.t2433 vp_p.t2950 vdd.t49 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3551 out_p.t2435 vp_p.t2951 vdd.t48 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3552 vdd.t47 vp_p.t2952 out_p.t2451 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3553 out_p.t2447 vp_p.t2953 vdd.t46 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3554 out_p.t2431 vp_p.t2954 vdd.t45 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3555 out_p.t2444 vp_p.t2955 vdd.t44 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3556 out_p.t2440 vp_p.t2956 vdd.t43 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3557 out_p.t2443 vp_p.t2957 vdd.t42 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3558 out_p.t2428 vp_p.t2958 vdd.t41 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3559 out_p.t2426 vp_p.t2959 vdd.t40 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3560 vdd.t39 vp_p.t2960 out_p.t2450 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3561 vdd.t38 vp_p.t2961 out_p.t2430 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3562 out_p.t2446 vp_p.t2962 vdd.t37 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3563 out_p.t2439 vp_p.t2963 vdd.t36 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3564 vdd.t35 vp_p.t2964 out_p.t2456 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3565 vdd.t34 vp_p.t2965 out_p.t2405 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3566 out_p.t2407 vp_p.t2966 vdd.t33 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3567 vdd.t32 vp_p.t2967 out_p.t2436 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3568 vdd.t31 vp_p.t2968 out_p.t2429 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3569 out_p.t2399 vp_p.t2969 vdd.t30 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3570 vdd.t29 vp_p.t2970 out_p.t2434 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3571 out_p.t2400 vp_p.t2971 vdd.t28 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3572 out_p.t2402 vp_p.t2972 vdd.t27 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3573 vdd.t26 vp_p.t2973 out_p.t2406 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3574 out_p.t2401 vp_p.t2974 vdd.t25 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3575 out_p.t2380 vp_p.t2975 vdd.t24 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3576 out_p.t1228 vp_p.t2976 vdd.t23 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3577 out_p.t1222 vp_p.t2977 vdd.t22 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3578 vdd.t21 vp_p.t2978 out_p.t1225 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3579 vdd.t20 vp_p.t2979 out_p.t1238 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3580 out_p.t1233 vp_p.t2980 vdd.t19 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3581 out_p.t1231 vp_p.t2981 vdd.t18 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3582 out_p.t1249 vp_p.t2982 vdd.t17 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3583 vdd.t16 vp_p.t2983 out_p.t1270 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3584 out_p.t1329 vp_p.t2984 vdd.t15 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3585 vdd.t14 vp_p.t2985 out_p.t1325 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3586 vdd.t13 vp_p.t2986 out_p.t1278 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3587 vdd.t12 vp_p.t2987 out_p.t1250 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3588 out_p.t1309 vp_p.t2988 vdd.t11 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3589 out_p.t1301 vp_p.t2989 vdd.t10 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3590 out_p.t1300 vp_p.t2990 vdd.t9 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3591 out_p.t1357 vp_p.t2991 vdd.t8 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3592 vdd.t7 vp_p.t2992 out_p.t1354 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3593 out_p.t1347 vp_p.t2993 vdd.t6 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3594 vdd.t5 vp_p.t2994 out_p.t456 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3595 vdd.t4 vp_p.t2995 out_p.t457 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3596 vdd.t3 vp_p.t2996 out_p.t452 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3597 out_p.t453 vp_p.t2997 vdd.t2 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3598 out_p.t449 vp_p.t2998 vdd.t1 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3599 out_p.t451 vp_p.t2999 vdd.t0 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
C0 vdd out_p 11129.80fF
C1 vp_p out_p 1913.30fF
C2 out_p vp_n 344.46fF
C3 vdd vp_p 3055.12fF
R0 vp_p.n8624 vp_p.t569 716.572
R1 vp_p.n7205 vp_p.t2489 716.572
R2 vp_p.n7203 vp_p.t2237 716.572
R3 vp_p.n7210 vp_p.t694 716.572
R4 vp_p.n7208 vp_p.t442 716.572
R5 vp_p.n5786 vp_p.t1719 716.572
R6 vp_p.n7215 vp_p.t860 716.572
R7 vp_p.n7213 vp_p.t623 716.572
R8 vp_p.n5791 vp_p.t1148 716.572
R9 vp_p.n4368 vp_p.t895 716.572
R10 vp_p.n7220 vp_p.t2057 716.572
R11 vp_p.n7218 vp_p.t1807 716.572
R12 vp_p.n5796 vp_p.t2808 716.572
R13 vp_p.n4373 vp_p.t2564 716.572
R14 vp_p.n2949 vp_p.t1444 716.572
R15 vp_p.n7225 vp_p.t585 716.572
R16 vp_p.n7223 vp_p.t318 716.572
R17 vp_p.n5801 vp_p.t501 716.572
R18 vp_p.n4378 vp_p.t239 716.572
R19 vp_p.n2954 vp_p.t2114 716.572
R20 vp_p.n1529 vp_p.t1711 716.572
R21 vp_p.n7230 vp_p.t1501 716.572
R22 vp_p.n7228 vp_p.t1251 716.572
R23 vp_p.n5806 vp_p.t2152 716.572
R24 vp_p.n4383 vp_p.t1902 716.572
R25 vp_p.n2959 vp_p.t759 716.572
R26 vp_p.n1534 vp_p.t351 716.572
R27 vp_p.n50 vp_p.t100 716.572
R28 vp_p.n7235 vp_p.t2673 716.572
R29 vp_p.n7233 vp_p.t2422 716.572
R30 vp_p.n5811 vp_p.t836 716.572
R31 vp_p.n4388 vp_p.t601 716.572
R32 vp_p.n2964 vp_p.t2440 716.572
R33 vp_p.n1539 vp_p.t2049 716.572
R34 vp_p.n55 vp_p.t1799 716.572
R35 vp_p.n8794 vp_p.t671 716.572
R36 vp_p.n7240 vp_p.t876 716.572
R37 vp_p.n7238 vp_p.t634 716.572
R38 vp_p.n5816 vp_p.t2515 716.572
R39 vp_p.n4393 vp_p.t2254 716.572
R40 vp_p.n2969 vp_p.t1146 716.572
R41 vp_p.n1544 vp_p.t719 716.572
R42 vp_p.n60 vp_p.t485 716.572
R43 vp_p.n8799 vp_p.t2334 716.572
R44 vp_p.n10301 vp_p.t2801 716.572
R45 vp_p.n7592 vp_p.t1054 716.572
R46 vp_p.n7590 vp_p.t794 716.572
R47 vp_p.n6168 vp_p.t2818 716.572
R48 vp_p.n4745 vp_p.t2569 716.572
R49 vp_p.n3321 vp_p.t1455 716.572
R50 vp_p.n1896 vp_p.t1046 716.572
R51 vp_p.n470 vp_p.t786 716.572
R52 vp_p.n9216 vp_p.t2646 716.572
R53 vp_p.n10653 vp_p.t127 716.572
R54 vp_p.n12091 vp_p.t2011 716.572
R55 vp_p.n26294 vp_p.t2807 716.572
R56 vp_p.n24869 vp_p.t2392 716.572
R57 vp_p.n23447 vp_p.t2162 716.572
R58 vp_p.n22024 vp_p.t1034 716.572
R59 vp_p.n20600 vp_p.t1514 716.572
R60 vp_p.n19175 vp_p.t363 716.572
R61 vp_p.n17749 vp_p.t2208 716.572
R62 vp_p.n16322 vp_p.t2671 716.572
R63 vp_p.n14894 vp_p.t2271 716.572
R64 vp_p.n13828 vp_p.t1589 716.572
R65 vp_p.n7565 vp_p.t2232 716.572
R66 vp_p.n7563 vp_p.t2026 716.572
R67 vp_p.n6141 vp_p.t1500 716.572
R68 vp_p.n4718 vp_p.t1250 716.572
R69 vp_p.n3294 vp_p.t103 716.572
R70 vp_p.n1869 vp_p.t2687 716.572
R71 vp_p.n385 vp_p.t2444 716.572
R72 vp_p.n9124 vp_p.t1326 716.572
R73 vp_p.n10626 vp_p.t1800 716.572
R74 vp_p.n12064 vp_p.t673 716.572
R75 vp_p.n26268 vp_p.t1040 716.572
R76 vp_p.n24842 vp_p.t621 716.572
R77 vp_p.n23420 vp_p.t368 716.572
R78 vp_p.n21997 vp_p.t2212 716.572
R79 vp_p.n20573 vp_p.t2698 716.572
R80 vp_p.n19148 vp_p.t1582 716.572
R81 vp_p.n17722 vp_p.t425 716.572
R82 vp_p.n16295 vp_p.t1354 716.572
R83 vp_p.n14867 vp_p.t791 716.572
R84 vp_p.n13823 vp_p.t233 716.572
R85 vp_p.n7606 vp_p.t118 716.572
R86 vp_p.n7604 vp_p.t2862 716.572
R87 vp_p.n6182 vp_p.t1182 716.572
R88 vp_p.n4759 vp_p.t920 716.572
R89 vp_p.n3335 vp_p.t2775 716.572
R90 vp_p.n1910 vp_p.t2370 716.572
R91 vp_p.n484 vp_p.t2138 716.572
R92 vp_p.n9230 vp_p.t997 716.572
R93 vp_p.n10667 vp_p.t1482 716.572
R94 vp_p.n12105 vp_p.t337 716.572
R95 vp_p.n26308 vp_p.t1898 716.572
R96 vp_p.n24883 vp_p.t1491 716.572
R97 vp_p.n23461 vp_p.t1236 716.572
R98 vp_p.n22038 vp_p.t93 716.572
R99 vp_p.n20614 vp_p.t590 716.572
R100 vp_p.n19189 vp_p.t2423 716.572
R101 vp_p.n17763 vp_p.t1310 716.572
R102 vp_p.n16336 vp_p.t1030 716.572
R103 vp_p.n14908 vp_p.t1557 716.572
R104 vp_p.n13818 vp_p.t2907 716.572
R105 vp_p.n7560 vp_p.t729 716.572
R106 vp_p.n7558 vp_p.t492 716.572
R107 vp_p.n6136 vp_p.t828 716.572
R108 vp_p.n4713 vp_p.t595 716.572
R109 vp_p.n3289 vp_p.t2431 716.572
R110 vp_p.n1864 vp_p.t2046 716.572
R111 vp_p.n380 vp_p.t1790 716.572
R112 vp_p.n9119 vp_p.t661 716.572
R113 vp_p.n10621 vp_p.t1134 716.572
R114 vp_p.n12059 vp_p.t2993 716.572
R115 vp_p.n26263 vp_p.t2499 716.572
R116 vp_p.n24837 vp_p.t2097 716.572
R117 vp_p.n23415 vp_p.t1856 716.572
R118 vp_p.n21992 vp_p.t710 716.572
R119 vp_p.n20568 vp_p.t1195 716.572
R120 vp_p.n19143 vp_p.t44 716.572
R121 vp_p.n17717 vp_p.t1907 716.572
R122 vp_p.n16290 vp_p.t683 716.572
R123 vp_p.n14862 vp_p.t1646 716.572
R124 vp_p.n13813 vp_p.t2558 716.572
R125 vp_p.n7620 vp_p.t1937 716.572
R126 vp_p.n7618 vp_p.t1703 716.572
R127 vp_p.n6196 vp_p.t2477 716.572
R128 vp_p.n4773 vp_p.t2228 716.572
R129 vp_p.n3349 vp_p.t1112 716.572
R130 vp_p.n1924 vp_p.t699 716.572
R131 vp_p.n498 vp_p.t450 716.572
R132 vp_p.n9244 vp_p.t2295 716.572
R133 vp_p.n10681 vp_p.t2774 716.572
R134 vp_p.n12119 vp_p.t1663 716.572
R135 vp_p.n26322 vp_p.t713 716.572
R136 vp_p.n24897 vp_p.t279 716.572
R137 vp_p.n23475 vp_p.t52 716.572
R138 vp_p.n22052 vp_p.t1913 716.572
R139 vp_p.n20628 vp_p.t2381 716.572
R140 vp_p.n19203 vp_p.t1255 716.572
R141 vp_p.n17777 vp_p.t109 716.572
R142 vp_p.n16350 vp_p.t2333 716.572
R143 vp_p.n14922 vp_p.t149 716.572
R144 vp_p.n13808 vp_p.t1237 716.572
R145 vp_p.n7555 vp_p.t568 716.572
R146 vp_p.n7553 vp_p.t301 716.572
R147 vp_p.n6131 vp_p.t1402 716.572
R148 vp_p.n4708 vp_p.t1161 716.572
R149 vp_p.n3284 vp_p.t17 716.572
R150 vp_p.n1859 vp_p.t2575 716.572
R151 vp_p.n375 vp_p.t2347 716.572
R152 vp_p.n9114 vp_p.t1220 716.572
R153 vp_p.n10616 vp_p.t1704 716.572
R154 vp_p.n12054 vp_p.t564 716.572
R155 vp_p.n26258 vp_p.t2321 716.572
R156 vp_p.n24832 vp_p.t1915 716.572
R157 vp_p.n23410 vp_p.t1682 716.572
R158 vp_p.n21987 vp_p.t543 716.572
R159 vp_p.n20563 vp_p.t1018 716.572
R160 vp_p.n19138 vp_p.t2857 716.572
R161 vp_p.n17712 vp_p.t1745 716.572
R162 vp_p.n16285 vp_p.t1240 716.572
R163 vp_p.n14857 vp_p.t1025 716.572
R164 vp_p.n13803 vp_p.t136 716.572
R165 vp_p.n7634 vp_p.t739 716.572
R166 vp_p.n7632 vp_p.t511 716.572
R167 vp_p.n6210 vp_p.t797 716.572
R168 vp_p.n4787 vp_p.t572 716.572
R169 vp_p.n3363 vp_p.t2407 716.572
R170 vp_p.n1938 vp_p.t2024 716.572
R171 vp_p.n512 vp_p.t1770 716.572
R172 vp_p.n9258 vp_p.t637 716.572
R173 vp_p.n10695 vp_p.t1109 716.572
R174 vp_p.n12133 vp_p.t2968 716.572
R175 vp_p.n26336 vp_p.t2521 716.572
R176 vp_p.n24911 vp_p.t2108 716.572
R177 vp_p.n23489 vp_p.t1873 716.572
R178 vp_p.n22066 vp_p.t727 716.572
R179 vp_p.n20642 vp_p.t1211 716.572
R180 vp_p.n19217 vp_p.t67 716.572
R181 vp_p.n17791 vp_p.t1930 716.572
R182 vp_p.n16364 vp_p.t666 716.572
R183 vp_p.n14936 vp_p.t1751 716.572
R184 vp_p.n13798 vp_p.t2540 716.572
R185 vp_p.n7550 vp_p.t1616 716.572
R186 vp_p.n7548 vp_p.t1378 716.572
R187 vp_p.n6126 vp_p.t493 716.572
R188 vp_p.n4703 vp_p.t232 716.572
R189 vp_p.n3279 vp_p.t2106 716.572
R190 vp_p.n1854 vp_p.t1701 716.572
R191 vp_p.n370 vp_p.t1447 716.572
R192 vp_p.n9109 vp_p.t291 716.572
R193 vp_p.n10611 vp_p.t778 716.572
R194 vp_p.n12049 vp_p.t2638 716.572
R195 vp_p.n26253 vp_p.t385 716.572
R196 vp_p.n24827 vp_p.t2975 716.572
R197 vp_p.n23405 vp_p.t2713 716.572
R198 vp_p.n21982 vp_p.t1600 716.572
R199 vp_p.n20558 vp_p.t2081 716.572
R200 vp_p.n19133 vp_p.t928 716.572
R201 vp_p.n17707 vp_p.t2785 716.572
R202 vp_p.n16280 vp_p.t328 716.572
R203 vp_p.n14852 vp_p.t2493 716.572
R204 vp_p.n13793 vp_p.t2213 716.572
R205 vp_p.n7648 vp_p.t589 716.572
R206 vp_p.n7646 vp_p.t329 716.572
R207 vp_p.n6224 vp_p.t1372 716.572
R208 vp_p.n4801 vp_p.t1129 716.572
R209 vp_p.n3377 vp_p.t2987 716.572
R210 vp_p.n1952 vp_p.t2554 716.572
R211 vp_p.n526 vp_p.t2319 716.572
R212 vp_p.n9272 vp_p.t1202 716.572
R213 vp_p.n10709 vp_p.t1679 716.572
R214 vp_p.n12147 vp_p.t541 716.572
R215 vp_p.n26350 vp_p.t2348 716.572
R216 vp_p.n24925 vp_p.t1938 716.572
R217 vp_p.n23503 vp_p.t1708 716.572
R218 vp_p.n22080 vp_p.t565 716.572
R219 vp_p.n20656 vp_p.t1045 716.572
R220 vp_p.n19231 vp_p.t2882 716.572
R221 vp_p.n17805 vp_p.t1763 716.572
R222 vp_p.n16378 vp_p.t1223 716.572
R223 vp_p.n14950 vp_p.t1128 716.572
R224 vp_p.n13788 vp_p.t105 716.572
R225 vp_p.n7545 vp_p.t417 716.572
R226 vp_p.n7543 vp_p.t191 716.572
R227 vp_p.n6121 vp_p.t1806 716.572
R228 vp_p.n4698 vp_p.t1569 716.572
R229 vp_p.n3274 vp_p.t411 716.572
R230 vp_p.n1849 vp_p.t6 716.572
R231 vp_p.n365 vp_p.t2739 716.572
R232 vp_p.n9104 vp_p.t1623 716.572
R233 vp_p.n10606 vp_p.t2104 716.572
R234 vp_p.n12044 vp_p.t956 716.572
R235 vp_p.n26248 vp_p.t2191 716.572
R236 vp_p.n24822 vp_p.t1791 716.572
R237 vp_p.n23400 vp_p.t1555 716.572
R238 vp_p.n21977 vp_p.t398 716.572
R239 vp_p.n20553 vp_p.t886 716.572
R240 vp_p.n19128 vp_p.t2727 716.572
R241 vp_p.n17702 vp_p.t1612 716.572
R242 vp_p.n16275 vp_p.t1656 716.572
R243 vp_p.n14847 vp_p.t1098 716.572
R244 vp_p.n13783 vp_p.t556 716.572
R245 vp_p.n7662 vp_p.t2063 716.572
R246 vp_p.n7660 vp_p.t1816 716.572
R247 vp_p.n6238 vp_p.t707 716.572
R248 vp_p.n4815 vp_p.t459 716.572
R249 vp_p.n3391 vp_p.t2309 716.572
R250 vp_p.n1966 vp_p.t1901 716.572
R251 vp_p.n540 vp_p.t1669 716.572
R252 vp_p.n9286 vp_p.t530 716.572
R253 vp_p.n10723 vp_p.t1003 716.572
R254 vp_p.n12161 vp_p.t2846 716.572
R255 vp_p.n26364 vp_p.t822 716.572
R256 vp_p.n24939 vp_p.t400 716.572
R257 vp_p.n23517 vp_p.t170 716.572
R258 vp_p.n22094 vp_p.t2044 716.572
R259 vp_p.n20670 vp_p.t2502 716.572
R260 vp_p.n19245 vp_p.t1374 716.572
R261 vp_p.n17819 vp_p.t227 716.572
R262 vp_p.n16392 vp_p.t559 716.572
R263 vp_p.n14964 vp_p.t1981 716.572
R264 vp_p.n13778 vp_p.t2433 716.572
R265 vp_p.n7540 vp_p.t249 716.572
R266 vp_p.n7538 vp_p.t20 716.572
R267 vp_p.n6116 vp_p.t2356 716.572
R268 vp_p.n4693 vp_p.t2121 716.572
R269 vp_p.n3269 vp_p.t979 716.572
R270 vp_p.n1844 vp_p.t575 716.572
R271 vp_p.n360 vp_p.t315 716.572
R272 vp_p.n9099 vp_p.t2181 716.572
R273 vp_p.n10601 vp_p.t2655 716.572
R274 vp_p.n12039 vp_p.t1541 716.572
R275 vp_p.n26243 vp_p.t2047 716.572
R276 vp_p.n24817 vp_p.t1618 716.572
R277 vp_p.n23395 vp_p.t1379 716.572
R278 vp_p.n21972 vp_p.t230 716.572
R279 vp_p.n20548 vp_p.t715 716.572
R280 vp_p.n19123 vp_p.t2561 716.572
R281 vp_p.n17697 vp_p.t1441 716.572
R282 vp_p.n16270 vp_p.t2199 716.572
R283 vp_p.n14842 vp_p.t484 716.572
R284 vp_p.n13773 vp_p.t1116 716.572
R285 vp_p.n7676 vp_p.t99 716.572
R286 vp_p.n7674 vp_p.t2847 716.572
R287 vp_p.n6252 vp_p.t2779 716.572
R288 vp_p.n4829 vp_p.t2538 716.572
R289 vp_p.n3405 vp_p.t1417 716.572
R290 vp_p.n1980 vp_p.t998 716.572
R291 vp_p.n554 vp_p.t746 716.572
R292 vp_p.n9300 vp_p.t2599 716.572
R293 vp_p.n10737 vp_p.t88 716.572
R294 vp_p.n12175 vp_p.t1965 716.572
R295 vp_p.n26378 vp_p.t1890 716.572
R296 vp_p.n24953 vp_p.t1477 716.572
R297 vp_p.n23531 vp_p.t1227 716.572
R298 vp_p.n22108 vp_p.t82 716.572
R299 vp_p.n20684 vp_p.t574 716.572
R300 vp_p.n19259 vp_p.t2411 716.572
R301 vp_p.n17833 vp_p.t1295 716.572
R302 vp_p.n16406 vp_p.t2630 716.572
R303 vp_p.n14978 vp_p.t451 716.572
R304 vp_p.n13768 vp_p.t1553 716.572
R305 vp_p.n7535 vp_p.t2079 716.572
R306 vp_p.n7533 vp_p.t1838 716.572
R307 vp_p.n6111 vp_p.t686 716.572
R308 vp_p.n4688 vp_p.t424 716.572
R309 vp_p.n3264 vp_p.t2279 716.572
R310 vp_p.n1839 vp_p.t1885 716.572
R311 vp_p.n355 vp_p.t1640 716.572
R312 vp_p.n9094 vp_p.t510 716.572
R313 vp_p.n10596 vp_p.t974 716.572
R314 vp_p.n12034 vp_p.t2827 716.572
R315 vp_p.n26238 vp_p.t848 716.572
R316 vp_p.n24812 vp_p.t420 716.572
R317 vp_p.n23390 vp_p.t193 716.572
R318 vp_p.n21967 vp_p.t2064 716.572
R319 vp_p.n20543 vp_p.t2523 716.572
R320 vp_p.n19118 vp_p.t1400 716.572
R321 vp_p.n17692 vp_p.t246 716.572
R322 vp_p.n16265 vp_p.t535 716.572
R323 vp_p.n14837 vp_p.t2082 716.572
R324 vp_p.n13763 vp_p.t2408 716.572
R325 vp_p.n7690 vp_p.t2929 716.572
R326 vp_p.n7688 vp_p.t2684 716.572
R327 vp_p.n6266 vp_p.t356 716.572
R328 vp_p.n4843 vp_p.t104 716.572
R329 vp_p.n3419 vp_p.t1989 716.572
R330 vp_p.n1994 vp_p.t1572 716.572
R331 vp_p.n568 vp_p.t1327 716.572
R332 vp_p.n9314 vp_p.t187 716.572
R333 vp_p.n10751 vp_p.t675 716.572
R334 vp_p.n12189 vp_p.t2522 716.572
R335 vp_p.n26392 vp_p.t1727 716.572
R336 vp_p.n24967 vp_p.t1300 716.572
R337 vp_p.n23545 vp_p.t1061 716.572
R338 vp_p.n22122 vp_p.t2901 716.572
R339 vp_p.n20698 vp_p.t389 716.572
R340 vp_p.n19273 vp_p.t2239 716.572
R341 vp_p.n17847 vp_p.t1126 716.572
R342 vp_p.n16420 vp_p.t212 716.572
R343 vp_p.n14992 vp_p.t2812 716.572
R344 vp_p.n13758 vp_p.t2109 716.572
R345 vp_p.n7530 vp_p.t2581 716.572
R346 vp_p.n7528 vp_p.t2352 716.572
R347 vp_p.n6106 vp_p.t2326 716.572
R348 vp_p.n4683 vp_p.t2098 716.572
R349 vp_p.n3259 vp_p.t943 716.572
R350 vp_p.n1834 vp_p.t547 716.572
R351 vp_p.n350 vp_p.t280 716.572
R352 vp_p.n9089 vp_p.t2160 716.572
R353 vp_p.n10591 vp_p.t2617 716.572
R354 vp_p.n12029 vp_p.t1505 716.572
R355 vp_p.n26233 vp_p.t1384 716.572
R356 vp_p.n24807 vp_p.t951 716.572
R357 vp_p.n23385 vp_p.t717 716.572
R358 vp_p.n21962 vp_p.t2563 716.572
R359 vp_p.n20538 vp_p.t55 716.572
R360 vp_p.n19113 vp_p.t1918 716.572
R361 vp_p.n17687 vp_p.t773 716.572
R362 vp_p.n16260 vp_p.t2176 716.572
R363 vp_p.n14832 vp_p.t2648 716.572
R364 vp_p.n13753 vp_p.t1081 716.572
R365 vp_p.n7704 vp_p.t474 716.572
R366 vp_p.n7702 vp_p.t220 716.572
R367 vp_p.n6280 vp_p.t2029 716.572
R368 vp_p.n4857 vp_p.t1775 716.572
R369 vp_p.n3433 vp_p.t640 716.572
R370 vp_p.n2008 vp_p.t218 716.572
R371 vp_p.n582 vp_p.t2970 716.572
R372 vp_p.n9328 vp_p.t1849 716.572
R373 vp_p.n10765 vp_p.t2296 716.572
R374 vp_p.n12203 vp_p.t1186 716.572
R375 vp_p.n26406 vp_p.t2227 716.572
R376 vp_p.n24981 vp_p.t1840 716.572
R377 vp_p.n23559 vp_p.t1593 716.572
R378 vp_p.n22136 vp_p.t447 716.572
R379 vp_p.n20712 vp_p.t918 716.572
R380 vp_p.n19287 vp_p.t2771 716.572
R381 vp_p.n17861 vp_p.t1659 716.572
R382 vp_p.n16434 vp_p.t1871 716.572
R383 vp_p.n15006 vp_p.t401 716.572
R384 vp_p.n13748 vp_p.t751 716.572
R385 vp_p.n7525 vp_p.t1346 716.572
R386 vp_p.n7523 vp_p.t1090 716.572
R387 vp_p.n6101 vp_p.t1709 716.572
R388 vp_p.n4678 vp_p.t1449 716.572
R389 vp_p.n3254 vp_p.t297 716.572
R390 vp_p.n1829 vp_p.t2880 716.572
R391 vp_p.n345 vp_p.t2641 716.572
R392 vp_p.n9084 vp_p.t1522 716.572
R393 vp_p.n10586 vp_p.t2004 716.572
R394 vp_p.n12024 vp_p.t858 716.572
R395 vp_p.n26228 vp_p.t102 716.572
R396 vp_p.n24802 vp_p.t2685 716.572
R397 vp_p.n23380 vp_p.t2438 716.572
R398 vp_p.n21957 vp_p.t1323 716.572
R399 vp_p.n20533 vp_p.t1798 716.572
R400 vp_p.n19108 vp_p.t669 716.572
R401 vp_p.n17682 vp_p.t2517 716.572
R402 vp_p.n16255 vp_p.t1548 716.572
R403 vp_p.n14827 vp_p.t1175 716.572
R404 vp_p.n13743 vp_p.t431 716.572
R405 vp_p.n7718 vp_p.t2262 716.572
R406 vp_p.n7716 vp_p.t2048 716.572
R407 vp_p.n6294 vp_p.t322 716.572
R408 vp_p.n4871 vp_p.t80 716.572
R409 vp_p.n3447 vp_p.t1950 716.572
R410 vp_p.n2022 vp_p.t1544 716.572
R411 vp_p.n596 vp_p.t1292 716.572
R412 vp_p.n9342 vp_p.t154 716.572
R413 vp_p.n10779 vp_p.t638 716.572
R414 vp_p.n12217 vp_p.t2483 716.572
R415 vp_p.n26420 vp_p.t1062 716.572
R416 vp_p.n24995 vp_p.t652 716.572
R417 vp_p.n23573 vp_p.t390 716.572
R418 vp_p.n22150 vp_p.t2240 716.572
R419 vp_p.n20726 vp_p.t2717 716.572
R420 vp_p.n19301 vp_p.t1602 716.572
R421 vp_p.n17875 vp_p.t465 716.572
R422 vp_p.n16448 vp_p.t181 716.572
R423 vp_p.n15020 vp_p.t2025 716.572
R424 vp_p.n13738 vp_p.t2088 716.572
R425 vp_p.n7520 vp_p.t150 716.572
R426 vp_p.n7518 vp_p.t2890 716.572
R427 vp_p.n6096 vp_p.t10 716.572
R428 vp_p.n4673 vp_p.t2744 716.572
R429 vp_p.n3249 vp_p.t1627 716.572
R430 vp_p.n1824 vp_p.t1216 716.572
R431 vp_p.n340 vp_p.t959 716.572
R432 vp_p.n9079 vp_p.t2814 716.572
R433 vp_p.n10581 vp_p.t292 716.572
R434 vp_p.n12019 vp_p.t2167 716.572
R435 vp_p.n26223 vp_p.t1921 716.572
R436 vp_p.n24797 vp_p.t1519 716.572
R437 vp_p.n23375 vp_p.t1265 716.572
R438 vp_p.n21952 vp_p.t124 716.572
R439 vp_p.n20528 vp_p.t614 716.572
R440 vp_p.n19103 vp_p.t2459 716.572
R441 vp_p.n17677 vp_p.t1342 716.572
R442 vp_p.n16250 vp_p.t2838 716.572
R443 vp_p.n14822 vp_p.t2742 716.572
R444 vp_p.n13733 vp_p.t1756 716.572
R445 vp_p.n7732 vp_p.t1089 716.572
R446 vp_p.n7730 vp_p.t849 716.572
R447 vp_p.n6308 vp_p.t1650 716.572
R448 vp_p.n4885 vp_p.t1405 716.572
R449 vp_p.n3461 vp_p.t255 716.572
R450 vp_p.n2036 vp_p.t2831 716.572
R451 vp_p.n610 vp_p.t2586 716.572
R452 vp_p.n9356 vp_p.t1475 716.572
R453 vp_p.n10793 vp_p.t1946 716.572
R454 vp_p.n12231 vp_p.t800 716.572
R455 vp_p.n26434 vp_p.t2850 716.572
R456 vp_p.n25009 vp_p.t2435 716.572
R457 vp_p.n23587 vp_p.t2194 716.572
R458 vp_p.n22164 vp_p.t1074 716.572
R459 vp_p.n20740 vp_p.t1558 716.572
R460 vp_p.n19315 vp_p.t403 716.572
R461 vp_p.n17889 vp_p.t2255 716.572
R462 vp_p.n16462 vp_p.t1499 716.572
R463 vp_p.n15034 vp_p.t616 716.572
R464 vp_p.n13728 vp_p.t387 716.572
R465 vp_p.n7515 vp_p.t1967 716.572
R466 vp_p.n7513 vp_p.t1729 716.572
R467 vp_p.n6091 vp_p.t1330 716.572
R468 vp_p.n4668 vp_p.t1079 716.572
R469 vp_p.n3244 vp_p.t2936 716.572
R470 vp_p.n1819 vp_p.t2524 716.572
R471 vp_p.n335 vp_p.t2266 716.572
R472 vp_p.n9074 vp_p.t1162 716.572
R473 vp_p.n10576 vp_p.t1624 716.572
R474 vp_p.n12014 vp_p.t499 716.572
R475 vp_p.n26218 vp_p.t732 716.572
R476 vp_p.n24792 vp_p.t311 716.572
R477 vp_p.n23370 vp_p.t75 716.572
R478 vp_p.n21947 vp_p.t1940 716.572
R479 vp_p.n20523 vp_p.t2399 716.572
R480 vp_p.n19098 vp_p.t1282 716.572
R481 vp_p.n17672 vp_p.t142 716.572
R482 vp_p.n16245 vp_p.t1181 716.572
R483 vp_p.n14817 vp_p.t1366 716.572
R484 vp_p.n13723 vp_p.t72 716.572
R485 vp_p.n7746 vp_p.t174 716.572
R486 vp_p.n7744 vp_p.t2913 716.572
R487 vp_p.n6322 vp_p.t2985 716.572
R488 vp_p.n4899 vp_p.t2722 716.572
R489 vp_p.n3475 vp_p.t1607 716.572
R490 vp_p.n2050 vp_p.t1200 716.572
R491 vp_p.n624 vp_p.t936 716.572
R492 vp_p.n9370 vp_p.t2792 716.572
R493 vp_p.n10807 vp_p.t273 716.572
R494 vp_p.n12245 vp_p.t2153 716.572
R495 vp_p.n26448 vp_p.t1944 716.572
R496 vp_p.n25023 vp_p.t1542 716.572
R497 vp_p.n23601 vp_p.t1288 716.572
R498 vp_p.n22178 vp_p.t151 716.572
R499 vp_p.n20754 vp_p.t633 716.572
R500 vp_p.n19329 vp_p.t2476 716.572
R501 vp_p.n17903 vp_p.t1360 716.572
R502 vp_p.n16476 vp_p.t2821 716.572
R503 vp_p.n15048 vp_p.t2848 716.572
R504 vp_p.n13718 vp_p.t1738 716.572
R505 vp_p.n7510 vp_p.t764 716.572
R506 vp_p.n7508 vp_p.t537 716.572
R507 vp_p.n6086 vp_p.t2624 716.572
R508 vp_p.n4663 vp_p.t2383 716.572
R509 vp_p.n3239 vp_p.t1261 716.572
R510 vp_p.n1814 vp_p.t846 716.572
R511 vp_p.n330 vp_p.t609 716.572
R512 vp_p.n9069 vp_p.t2456 716.572
R513 vp_p.n10571 vp_p.t2930 716.572
R514 vp_p.n12009 vp_p.t1813 716.572
R515 vp_p.n26213 vp_p.t2536 716.572
R516 vp_p.n24787 vp_p.t2139 716.572
R517 vp_p.n23365 vp_p.t1892 716.572
R518 vp_p.n21942 vp_p.t744 716.572
R519 vp_p.n20518 vp_p.t1231 716.572
R520 vp_p.n19093 vp_p.t85 716.572
R521 vp_p.n17667 vp_p.t1961 716.572
R522 vp_p.n16240 vp_p.t2478 716.572
R523 vp_p.n14812 vp_p.t2954 716.572
R524 vp_p.n13713 vp_p.t1397 716.572
R525 vp_p.n7760 vp_p.t1994 716.572
R526 vp_p.n7758 vp_p.t1742 716.572
R527 vp_p.n6336 vp_p.t1304 716.572
R528 vp_p.n4913 vp_p.t1063 716.572
R529 vp_p.n3489 vp_p.t2908 716.572
R530 vp_p.n2064 vp_p.t2500 716.572
R531 vp_p.n638 vp_p.t2243 716.572
R532 vp_p.n9384 vp_p.t1130 716.572
R533 vp_p.n10821 vp_p.t1606 716.572
R534 vp_p.n12259 vp_p.t471 716.572
R535 vp_p.n26462 vp_p.t747 716.572
R536 vp_p.n25037 vp_p.t340 716.572
R537 vp_p.n23615 vp_p.t89 716.572
R538 vp_p.n22192 vp_p.t1968 716.572
R539 vp_p.n20768 vp_p.t2420 716.572
R540 vp_p.n19343 vp_p.t1302 716.572
R541 vp_p.n17917 vp_p.t166 716.572
R542 vp_p.n16490 vp_p.t1165 716.572
R543 vp_p.n15062 vp_p.t1472 716.572
R544 vp_p.n13708 vp_p.t50 716.572
R545 vp_p.n7505 vp_p.t613 716.572
R546 vp_p.n7503 vp_p.t359 716.572
R547 vp_p.n6081 vp_p.t208 716.572
R548 vp_p.n4658 vp_p.t2955 716.572
R549 vp_p.n3234 vp_p.t1833 716.572
R550 vp_p.n1809 vp_p.t1409 716.572
R551 vp_p.n325 vp_p.t1176 716.572
R552 vp_p.n9064 vp_p.t32 716.572
R553 vp_p.n10566 vp_p.t512 716.572
R554 vp_p.n12004 vp_p.t2364 716.572
R555 vp_p.n26208 vp_p.t2371 716.572
R556 vp_p.n24782 vp_p.t1971 716.572
R557 vp_p.n23360 vp_p.t1731 716.572
R558 vp_p.n21937 vp_p.t593 716.572
R559 vp_p.n20513 vp_p.t1067 716.572
R560 vp_p.n19088 vp_p.t2910 716.572
R561 vp_p.n17662 vp_p.t1788 716.572
R562 vp_p.n16235 vp_p.t53 716.572
R563 vp_p.n14807 vp_p.t2329 716.572
R564 vp_p.n13703 vp_p.t1958 716.572
R565 vp_p.n7774 vp_p.t455 716.572
R566 vp_p.n7772 vp_p.t214 716.572
R567 vp_p.n6350 vp_p.t643 716.572
R568 vp_p.n4927 vp_p.t386 716.572
R569 vp_p.n3503 vp_p.t2236 716.572
R570 vp_p.n2078 vp_p.t1853 716.572
R571 vp_p.n652 vp_p.t1601 716.572
R572 vp_p.n9398 vp_p.t462 716.572
R573 vp_p.n10835 vp_p.t927 716.572
R574 vp_p.n12273 vp_p.t2783 716.572
R575 vp_p.n26476 vp_p.t2209 716.572
R576 vp_p.n25051 vp_p.t1821 716.572
R577 vp_p.n23629 vp_p.t1578 716.572
R578 vp_p.n22206 vp_p.t422 716.572
R579 vp_p.n20782 vp_p.t905 716.572
R580 vp_p.n19357 vp_p.t2756 716.572
R581 vp_p.n17931 vp_p.t1639 716.572
R582 vp_p.n16504 vp_p.t494 716.572
R583 vp_p.n15076 vp_p.t2292 716.572
R584 vp_p.n13698 vp_p.t2375 716.572
R585 vp_p.n7500 vp_p.t1670 716.572
R586 vp_p.n7498 vp_p.t1420 716.572
R587 vp_p.n6076 vp_p.t2276 716.572
R588 vp_p.n4653 vp_p.t2065 716.572
R589 vp_p.n3229 vp_p.t910 716.572
R590 vp_p.n1804 vp_p.t507 716.572
R591 vp_p.n320 vp_p.t248 716.572
R592 vp_p.n9059 vp_p.t2122 716.572
R593 vp_p.n10561 vp_p.t2579 716.572
R594 vp_p.n11999 vp_p.t1468 716.572
R595 vp_p.n26203 vp_p.t426 716.572
R596 vp_p.n24777 vp_p.t26 716.572
R597 vp_p.n23355 vp_p.t2758 716.572
R598 vp_p.n21932 vp_p.t1641 716.572
R599 vp_p.n20508 vp_p.t2120 716.572
R600 vp_p.n19083 vp_p.t976 716.572
R601 vp_p.n17657 vp_p.t2828 716.572
R602 vp_p.n16230 vp_p.t2148 716.572
R603 vp_p.n14802 vp_p.t814 716.572
R604 vp_p.n13693 vp_p.t1052 716.572
R605 vp_p.n7788 vp_p.t269 716.572
R606 vp_p.n7786 vp_p.t40 716.572
R607 vp_p.n6364 vp_p.t1206 716.572
R608 vp_p.n4941 vp_p.t944 716.572
R609 vp_p.n3517 vp_p.t2800 716.572
R610 vp_p.n2092 vp_p.t2388 716.572
R611 vp_p.n666 vp_p.t2161 716.572
R612 vp_p.n9412 vp_p.t1027 716.572
R613 vp_p.n10849 vp_p.t1506 716.572
R614 vp_p.n12287 vp_p.t361 716.572
R615 vp_p.n26490 vp_p.t2069 716.572
R616 vp_p.n25065 vp_p.t1643 716.572
R617 vp_p.n23643 vp_p.t1404 716.572
R618 vp_p.n22220 vp_p.t251 716.572
R619 vp_p.n20796 vp_p.t734 716.572
R620 vp_p.n19371 vp_p.t2585 716.572
R621 vp_p.n17945 vp_p.t1474 716.572
R622 vp_p.n16518 vp_p.t1055 716.572
R623 vp_p.n15090 vp_p.t1702 716.572
R624 vp_p.n13688 vp_p.t2940 716.572
R625 vp_p.n7495 vp_p.t480 716.572
R626 vp_p.n7493 vp_p.t226 716.572
R627 vp_p.n6071 vp_p.t622 716.572
R628 vp_p.n4648 vp_p.t369 716.572
R629 vp_p.n3224 vp_p.t2214 716.572
R630 vp_p.n1799 vp_p.t1824 716.572
R631 vp_p.n315 vp_p.t1583 716.572
R632 vp_p.n9054 vp_p.t427 716.572
R633 vp_p.n10556 vp_p.t906 716.572
R634 vp_p.n11994 vp_p.t2757 716.572
R635 vp_p.n26198 vp_p.t2230 716.572
R636 vp_p.n24772 vp_p.t1846 716.572
R637 vp_p.n23350 vp_p.t1597 716.572
R638 vp_p.n21927 vp_p.t453 716.572
R639 vp_p.n20503 vp_p.t921 716.572
R640 vp_p.n19078 vp_p.t2776 716.572
R641 vp_p.n17652 vp_p.t1664 716.572
R642 vp_p.n16225 vp_p.t464 716.572
R643 vp_p.n14797 vp_p.t2398 716.572
R644 vp_p.n13683 vp_p.t2355 716.572
R645 vp_p.n7802 vp_p.t2102 716.572
R646 vp_p.n7800 vp_p.t1864 716.572
R647 vp_p.n6378 vp_p.t2509 716.572
R648 vp_p.n4955 vp_p.t2250 716.572
R649 vp_p.n3531 vp_p.t1143 716.572
R650 vp_p.n2106 vp_p.t718 716.572
R651 vp_p.n680 vp_p.t481 716.572
R652 vp_p.n9426 vp_p.t2330 716.572
R653 vp_p.n10863 vp_p.t2796 716.572
R654 vp_p.n12301 vp_p.t1689 716.572
R655 vp_p.n26504 vp_p.t878 716.572
R656 vp_p.n25079 vp_p.t457 716.572
R657 vp_p.n23657 vp_p.t215 716.572
R658 vp_p.n22234 vp_p.t2083 716.572
R659 vp_p.n20810 vp_p.t2539 716.572
R660 vp_p.n19385 vp_p.t1418 716.572
R661 vp_p.n17959 vp_p.t264 716.572
R662 vp_p.n16532 vp_p.t2357 716.572
R663 vp_p.n15104 vp_p.t274 716.572
R664 vp_p.n13678 vp_p.t1263 716.572
R665 vp_p.n7490 vp_p.t288 716.572
R666 vp_p.n7488 vp_p.t62 716.572
R667 vp_p.n6066 vp_p.t1184 716.572
R668 vp_p.n4643 vp_p.t924 716.572
R669 vp_p.n3219 vp_p.t2780 716.572
R670 vp_p.n1794 vp_p.t2372 716.572
R671 vp_p.n310 vp_p.t2140 716.572
R672 vp_p.n9049 vp_p.t999 716.572
R673 vp_p.n10551 vp_p.t1487 716.572
R674 vp_p.n11989 vp_p.t341 716.572
R675 vp_p.n26193 vp_p.t2089 716.572
R676 vp_p.n24767 vp_p.t1672 716.572
R677 vp_p.n23345 vp_p.t1421 716.572
R678 vp_p.n21922 vp_p.t270 716.572
R679 vp_p.n20498 vp_p.t749 716.572
R680 vp_p.n19073 vp_p.t2603 716.572
R681 vp_p.n17647 vp_p.t1495 716.572
R682 vp_p.n16220 vp_p.t1031 716.572
R683 vp_p.n14792 vp_p.t1796 716.572
R684 vp_p.n13673 vp_p.t2914 716.572
R685 vp_p.n7816 vp_p.t158 716.572
R686 vp_p.n7814 vp_p.t2897 716.572
R687 vp_p.n6392 vp_p.t1609 716.572
R688 vp_p.n4969 vp_p.t1368 716.572
R689 vp_p.n3545 vp_p.t224 716.572
R690 vp_p.n2120 vp_p.t2793 716.572
R691 vp_p.n694 vp_p.t2551 716.572
R692 vp_p.n9440 vp_p.t1430 716.572
R693 vp_p.n10877 vp_p.t1906 716.572
R694 vp_p.n12315 vp_p.t763 716.572
R695 vp_p.n26518 vp_p.t1931 716.572
R696 vp_p.n25093 vp_p.t1523 716.572
R697 vp_p.n23671 vp_p.t1271 716.572
R698 vp_p.n22248 vp_p.t128 716.572
R699 vp_p.n20824 vp_p.t619 716.572
R700 vp_p.n19399 vp_p.t2467 716.572
R701 vp_p.n17973 vp_p.t1348 716.572
R702 vp_p.n16546 vp_p.t1461 716.572
R703 vp_p.n15118 vp_p.t1772 716.572
R704 vp_p.n13668 vp_p.t355 716.572
R705 vp_p.n7485 vp_p.t1784 716.572
R706 vp_p.n7483 vp_p.t1545 716.572
R707 vp_p.n6061 vp_p.t519 716.572
R708 vp_p.n4638 vp_p.t256 716.572
R709 vp_p.n3214 vp_p.t2133 716.572
R710 vp_p.n1789 vp_p.t1725 716.572
R711 vp_p.n305 vp_p.t1478 716.572
R712 vp_p.n9044 vp_p.t330 716.572
R713 vp_p.n10546 vp_p.t801 716.572
R714 vp_p.n11984 vp_p.t2663 716.572
R715 vp_p.n26188 vp_p.t562 716.572
R716 vp_p.n24762 vp_p.t132 716.572
R717 vp_p.n23340 vp_p.t2878 716.572
R718 vp_p.n21917 vp_p.t1758 716.572
R719 vp_p.n20493 vp_p.t2215 716.572
R720 vp_p.n19068 vp_p.t1094 716.572
R721 vp_p.n17642 vp_p.t2956 716.572
R722 vp_p.n16215 vp_p.t357 716.572
R723 vp_p.n14787 vp_p.t2621 716.572
R724 vp_p.n13663 vp_p.t2238 716.572
R725 vp_p.n7830 vp_p.t2983 716.572
R726 vp_p.n7828 vp_p.t2721 716.572
R727 vp_p.n6406 vp_p.t2168 716.572
R728 vp_p.n4983 vp_p.t1925 716.572
R729 vp_p.n3559 vp_p.t781 716.572
R730 vp_p.n2134 vp_p.t372 716.572
R731 vp_p.n708 vp_p.t126 716.572
R732 vp_p.n9454 vp_p.t2007 716.572
R733 vp_p.n10891 vp_p.t2462 716.572
R734 vp_p.n12329 vp_p.t1345 716.572
R735 vp_p.n26532 vp_p.t1764 716.572
R736 vp_p.n25107 vp_p.t1355 716.572
R737 vp_p.n23685 vp_p.t1101 716.572
R738 vp_p.n22262 vp_p.t2961 716.572
R739 vp_p.n20838 vp_p.t436 716.572
R740 vp_p.n19413 vp_p.t2286 716.572
R741 vp_p.n17987 vp_p.t1178 716.572
R742 vp_p.n16560 vp_p.t2038 716.572
R743 vp_p.n15132 vp_p.t1155 716.572
R744 vp_p.n13658 vp_p.t911 716.572
R745 vp_p.n7480 vp_p.t600 716.572
R746 vp_p.n7478 vp_p.t345 716.572
R747 vp_p.n6056 vp_p.t1834 716.572
R748 vp_p.n4633 vp_p.t1590 716.572
R749 vp_p.n3209 vp_p.t444 716.572
R750 vp_p.n1784 vp_p.t33 716.572
R751 vp_p.n300 vp_p.t2769 716.572
R752 vp_p.n9039 vp_p.t1655 716.572
R753 vp_p.n10541 vp_p.t2129 716.572
R754 vp_p.n11979 vp_p.t989 716.572
R755 vp_p.n26183 vp_p.t2359 716.572
R756 vp_p.n24757 vp_p.t1951 716.572
R757 vp_p.n23335 vp_p.t1720 716.572
R758 vp_p.n21912 vp_p.t577 716.572
R759 vp_p.n20488 vp_p.t1056 716.572
R760 vp_p.n19063 vp_p.t2895 716.572
R761 vp_p.n17637 vp_p.t1779 716.572
R762 vp_p.n16210 vp_p.t1683 716.572
R763 vp_p.n14782 vp_p.t1235 716.572
R764 vp_p.n13653 vp_p.t587 716.572
R765 vp_p.n7844 vp_p.t1802 716.572
R766 vp_p.n7842 vp_p.t1563 716.572
R767 vp_p.n6420 vp_p.t497 716.572
R768 vp_p.n4997 vp_p.t235 716.572
R769 vp_p.n3573 vp_p.t2110 716.572
R770 vp_p.n2148 vp_p.t1705 716.572
R771 vp_p.n722 vp_p.t1450 716.572
R772 vp_p.n9468 vp_p.t296 716.572
R773 vp_p.n10905 vp_p.t779 716.572
R774 vp_p.n12343 vp_p.t2640 716.572
R775 vp_p.n26546 vp_p.t586 716.572
R776 vp_p.n25121 vp_p.t159 716.572
R777 vp_p.n23699 vp_p.t2898 716.572
R778 vp_p.n22276 vp_p.t1782 716.572
R779 vp_p.n20852 vp_p.t2233 716.572
R780 vp_p.n19427 vp_p.t1121 716.572
R781 vp_p.n18001 vp_p.t2978 716.572
R782 vp_p.n16574 vp_p.t335 716.572
R783 vp_p.n15146 vp_p.t2723 716.572
R784 vp_p.n13648 vp_p.t2218 716.572
R785 vp_p.n7475 vp_p.t2656 716.572
R786 vp_p.n7473 vp_p.t2403 716.572
R787 vp_p.n6051 vp_p.t171 716.572
R788 vp_p.n4628 vp_p.t2911 716.572
R789 vp_p.n3204 vp_p.t1789 716.572
R790 vp_p.n1779 vp_p.t1375 716.572
R791 vp_p.n295 vp_p.t1131 716.572
R792 vp_p.n9034 vp_p.t2988 716.572
R793 vp_p.n10536 vp_p.t472 716.572
R794 vp_p.n11974 vp_p.t2320 716.572
R795 vp_p.n26178 vp_p.t1442 716.572
R796 vp_p.n24752 vp_p.t1032 716.572
R797 vp_p.n23330 vp_p.t771 716.572
R798 vp_p.n21907 vp_p.t2631 716.572
R799 vp_p.n20483 vp_p.t113 716.572
R800 vp_p.n19058 vp_p.t1996 716.572
R801 vp_p.n17632 vp_p.t850 716.572
R802 vp_p.n16205 vp_p.t21 716.572
R803 vp_p.n14777 vp_p.t504 716.572
R804 vp_p.n13643 vp_p.t1912 716.572
R805 vp_p.n7858 vp_p.t2313 716.572
R806 vp_p.n7856 vp_p.t2092 716.572
R807 vp_p.n6434 vp_p.t2141 716.572
R808 vp_p.n5011 vp_p.t1897 716.572
R809 vp_p.n3587 vp_p.t752 716.572
R810 vp_p.n2162 vp_p.t343 716.572
R811 vp_p.n736 vp_p.t94 716.572
R812 vp_p.n9482 vp_p.t1975 716.572
R813 vp_p.n10919 vp_p.t2424 716.572
R814 vp_p.n12357 vp_p.t1311 716.572
R815 vp_p.n26560 vp_p.t1102 716.572
R816 vp_p.n25135 vp_p.t692 716.572
R817 vp_p.n23713 vp_p.t437 716.572
R818 vp_p.n22290 vp_p.t2287 716.572
R819 vp_p.n20866 vp_p.t2764 716.572
R820 vp_p.n19441 vp_p.t1651 716.572
R821 vp_p.n18015 vp_p.t520 716.572
R822 vp_p.n16588 vp_p.t2002 716.572
R823 vp_p.n15160 vp_p.t316 716.572
R824 vp_p.n13638 vp_p.t890 716.572
R825 vp_p.n7470 vp_p.t200 716.572
R826 vp_p.n7468 vp_p.t2945 716.572
R827 vp_p.n6046 vp_p.t1827 716.572
R828 vp_p.n4623 vp_p.t1584 716.572
R829 vp_p.n3199 vp_p.t432 716.572
R830 vp_p.n1774 vp_p.t28 716.572
R831 vp_p.n290 vp_p.t2759 716.572
R832 vp_p.n9029 vp_p.t1647 716.572
R833 vp_p.n10531 vp_p.t2126 716.572
R834 vp_p.n11969 vp_p.t982 716.572
R835 vp_p.n26173 vp_p.t1982 716.572
R836 vp_p.n24747 vp_p.t1565 716.572
R837 vp_p.n23325 vp_p.t1317 716.572
R838 vp_p.n21902 vp_p.t177 716.572
R839 vp_p.n20478 vp_p.t662 716.572
R840 vp_p.n19053 vp_p.t2510 716.572
R841 vp_p.n17627 vp_p.t1386 716.572
R842 vp_p.n16200 vp_p.t1680 716.572
R843 vp_p.n14772 vp_p.t1077 716.572
R844 vp_p.n13633 vp_p.t578 716.572
R845 vp_p.n7872 vp_p.t1825 716.572
R846 vp_p.n7870 vp_p.t1581 716.572
R847 vp_p.n6448 vp_p.t720 716.572
R848 vp_p.n5025 vp_p.t486 716.572
R849 vp_p.n3601 vp_p.t2335 716.572
R850 vp_p.n2176 vp_p.t1922 716.572
R851 vp_p.n750 vp_p.t1692 716.572
R852 vp_p.n9496 vp_p.t551 716.572
R853 vp_p.n10933 vp_p.t1028 716.572
R854 vp_p.n12371 vp_p.t2871 716.572
R855 vp_p.n26574 vp_p.t603 716.572
R856 vp_p.n25149 vp_p.t179 716.572
R857 vp_p.n23727 vp_p.t2922 716.572
R858 vp_p.n22304 vp_p.t1803 716.572
R859 vp_p.n20880 vp_p.t2252 716.572
R860 vp_p.n19455 vp_p.t1145 716.572
R861 vp_p.n18029 vp_p.t1 716.572
R862 vp_p.n16602 vp_p.t584 716.572
R863 vp_p.n15174 vp_p.t1952 716.572
R864 vp_p.n13628 vp_p.t2460 716.572
R865 vp_p.n7465 vp_p.t2022 716.572
R866 vp_p.n7463 vp_p.t1766 716.572
R867 vp_p.n6041 vp_p.t133 716.572
R868 vp_p.n4618 vp_p.t2877 716.572
R869 vp_p.n3194 vp_p.t1757 716.572
R870 vp_p.n1769 vp_p.t1350 716.572
R871 vp_p.n285 vp_p.t1095 716.572
R872 vp_p.n9024 vp_p.t2957 716.572
R873 vp_p.n10526 vp_p.t428 716.572
R874 vp_p.n11964 vp_p.t2280 716.572
R875 vp_p.n26168 vp_p.t774 716.572
R876 vp_p.n24742 vp_p.t364 716.572
R877 vp_p.n23320 vp_p.t114 716.572
R878 vp_p.n21897 vp_p.t2000 716.572
R879 vp_p.n20473 vp_p.t2450 716.572
R880 vp_p.n19048 vp_p.t1334 716.572
R881 vp_p.n17622 vp_p.t195 716.572
R882 vp_p.n16195 vp_p.t2984 716.572
R883 vp_p.n14767 vp_p.t2667 716.572
R884 vp_p.n13623 vp_p.t1887 716.572
R885 vp_p.n7886 vp_p.t2858 716.572
R886 vp_p.n7884 vp_p.t2615 716.572
R887 vp_p.n6462 vp_p.t2797 716.572
R888 vp_p.n5039 vp_p.t2553 716.572
R889 vp_p.n3615 vp_p.t1434 716.572
R890 vp_p.n2190 vp_p.t1024 716.572
R891 vp_p.n764 vp_p.t766 716.572
R892 vp_p.n9510 vp_p.t2622 716.572
R893 vp_p.n10947 vp_p.t106 716.572
R894 vp_p.n12385 vp_p.t1992 716.572
R895 vp_p.n26588 vp_p.t1660 716.572
R896 vp_p.n25163 vp_p.t1234 716.572
R897 vp_p.n23741 vp_p.t990 716.572
R898 vp_p.n22318 vp_p.t2836 716.572
R899 vp_p.n20894 vp_p.t326 716.572
R900 vp_p.n19469 vp_p.t2188 716.572
R901 vp_p.n18043 vp_p.t1064 716.572
R902 vp_p.n16616 vp_p.t2653 716.572
R903 vp_p.n15188 vp_p.t418 716.572
R904 vp_p.n13618 vp_p.t1573 716.572
R905 vp_p.n7460 vp_p.t1848 716.572
R906 vp_p.n7458 vp_p.t1598 716.572
R907 vp_p.n6036 vp_p.t702 716.572
R908 vp_p.n4613 vp_p.t458 716.572
R909 vp_p.n3189 vp_p.t2303 716.572
R910 vp_p.n1764 vp_p.t1900 716.572
R911 vp_p.n280 vp_p.t1668 716.572
R912 vp_p.n9019 vp_p.t528 716.572
R913 vp_p.n10521 vp_p.t1000 716.572
R914 vp_p.n11959 vp_p.t2843 716.572
R915 vp_p.n26163 vp_p.t620 716.572
R916 vp_p.n24737 vp_p.t201 716.572
R917 vp_p.n23315 vp_p.t2948 716.572
R918 vp_p.n21892 vp_p.t1822 716.572
R919 vp_p.n20468 vp_p.t2275 716.572
R920 vp_p.n19043 vp_p.t1170 716.572
R921 vp_p.n17617 vp_p.t25 716.572
R922 vp_p.n16190 vp_p.t557 716.572
R923 vp_p.n14762 vp_p.t2066 716.572
R924 vp_p.n13613 vp_p.t2427 716.572
R925 vp_p.n7900 vp_p.t1700 716.572
R926 vp_p.n7898 vp_p.t1446 716.572
R927 vp_p.n6476 vp_p.t1137 716.572
R928 vp_p.n5053 vp_p.t888 716.572
R929 vp_p.n3629 vp_p.t2732 716.572
R930 vp_p.n2204 vp_p.t2327 716.572
R931 vp_p.n778 vp_p.t2099 716.572
R932 vp_p.n9524 vp_p.t945 716.572
R933 vp_p.n10961 vp_p.t1431 716.572
R934 vp_p.n12399 vp_p.t281 716.572
R935 vp_p.n26602 vp_p.t466 716.572
R936 vp_p.n25177 vp_p.t45 716.572
R937 vp_p.n23755 vp_p.t2790 716.572
R938 vp_p.n22332 vp_p.t1676 716.572
R939 vp_p.n20908 vp_p.t2149 716.572
R940 vp_p.n19483 vp_p.t1016 716.572
R941 vp_p.n18057 vp_p.t2855 716.572
R942 vp_p.n16630 vp_p.t973 716.572
R943 vp_p.n15202 vp_p.t2043 716.572
R944 vp_p.n13608 vp_p.t2863 716.572
R945 vp_p.n7455 vp_p.t657 716.572
R946 vp_p.n7453 vp_p.t397 716.572
R947 vp_p.n6031 vp_p.t2032 716.572
R948 vp_p.n4608 vp_p.t1776 716.572
R949 vp_p.n3184 vp_p.t642 716.572
R950 vp_p.n1759 vp_p.t219 716.572
R951 vp_p.n275 vp_p.t2974 716.572
R952 vp_p.n9014 vp_p.t1852 716.572
R953 vp_p.n10516 vp_p.t2299 716.572
R954 vp_p.n11954 vp_p.t1190 716.572
R955 vp_p.n26158 vp_p.t2405 716.572
R956 vp_p.n24732 vp_p.t2021 716.572
R957 vp_p.n23310 vp_p.t1769 716.572
R958 vp_p.n21887 vp_p.t636 716.572
R959 vp_p.n20463 vp_p.t1107 716.572
R960 vp_p.n19038 vp_p.t2966 716.572
R961 vp_p.n17612 vp_p.t1845 716.572
R962 vp_p.n16185 vp_p.t1872 716.572
R963 vp_p.n14757 vp_p.t665 716.572
R964 vp_p.n13603 vp_p.t757 716.572
R965 vp_p.n7914 vp_p.t1527 716.572
R966 vp_p.n7912 vp_p.t1273 716.572
R967 vp_p.n6490 vp_p.t1710 716.572
R968 vp_p.n5067 vp_p.t1454 716.572
R969 vp_p.n3643 vp_p.t300 716.572
R970 vp_p.n2218 vp_p.t2883 716.572
R971 vp_p.n792 vp_p.t2644 716.572
R972 vp_p.n9538 vp_p.t1529 716.572
R973 vp_p.n10975 vp_p.t2008 716.572
R974 vp_p.n12413 vp_p.t863 716.572
R975 vp_p.n26616 vp_p.t276 716.572
R976 vp_p.n25191 vp_p.t2856 716.572
R977 vp_p.n23769 vp_p.t2614 716.572
R978 vp_p.n22346 vp_p.t1503 716.572
R979 vp_p.n20922 vp_p.t1986 716.572
R980 vp_p.n19497 vp_p.t840 716.572
R981 vp_p.n18071 vp_p.t2690 716.572
R982 vp_p.n16644 vp_p.t1552 716.572
R983 vp_p.n15216 vp_p.t1408 716.572
R984 vp_p.n13598 vp_p.t434 716.572
R985 vp_p.n7450 vp_p.t1722 716.572
R986 vp_p.n7448 vp_p.t1470 716.572
R987 vp_p.n6026 vp_p.t1111 716.572
R988 vp_p.n4603 vp_p.t872 716.572
R989 vp_p.n3179 vp_p.t2709 716.572
R990 vp_p.n1754 vp_p.t2294 716.572
R991 vp_p.n270 vp_p.t2077 716.572
R992 vp_p.n9009 vp_p.t923 716.572
R993 vp_p.n10511 vp_p.t1412 716.572
R994 vp_p.n11949 vp_p.t262 716.572
R995 vp_p.n26153 vp_p.t491 716.572
R996 vp_p.n24727 vp_p.t66 716.572
R997 vp_p.n23305 vp_p.t2809 716.572
R998 vp_p.n21882 vp_p.t1697 716.572
R999 vp_p.n20458 vp_p.t2163 716.572
R1000 vp_p.n19033 vp_p.t1038 716.572
R1001 vp_p.n17607 vp_p.t2875 716.572
R1002 vp_p.n16180 vp_p.t949 716.572
R1003 vp_p.n14752 vp_p.t2136 716.572
R1004 vp_p.n13593 vp_p.t2837 716.572
R1005 vp_p.n7928 vp_p.t321 716.572
R1006 vp_p.n7926 vp_p.t79 716.572
R1007 vp_p.n6504 vp_p.t16 716.572
R1008 vp_p.n5081 vp_p.t2745 716.572
R1009 vp_p.n3657 vp_p.t1630 716.572
R1010 vp_p.n2232 vp_p.t1218 716.572
R1011 vp_p.n806 vp_p.t962 716.572
R1012 vp_p.n9552 vp_p.t2817 716.572
R1013 vp_p.n10989 vp_p.t295 716.572
R1014 vp_p.n12427 vp_p.t2169 716.572
R1015 vp_p.n26630 vp_p.t2107 716.572
R1016 vp_p.n25205 vp_p.t1699 716.572
R1017 vp_p.n23783 vp_p.t1445 716.572
R1018 vp_p.n22360 vp_p.t290 716.572
R1019 vp_p.n20936 vp_p.t777 716.572
R1020 vp_p.n19511 vp_p.t2637 716.572
R1021 vp_p.n18085 vp_p.t1521 716.572
R1022 vp_p.n16658 vp_p.t2841 716.572
R1023 vp_p.n15230 vp_p.t5 716.572
R1024 vp_p.n13588 vp_p.t1761 716.572
R1025 vp_p.n7445 vp_p.t1209 716.572
R1026 vp_p.n7443 vp_p.t942 716.572
R1027 vp_p.n6021 vp_p.t2677 716.572
R1028 vp_p.n4598 vp_p.t2426 716.572
R1029 vp_p.n3174 vp_p.t1315 716.572
R1030 vp_p.n1749 vp_p.t892 716.572
R1031 vp_p.n265 vp_p.t659 716.572
R1032 vp_p.n9004 vp_p.t2507 716.572
R1033 vp_p.n10506 vp_p.t2990 716.572
R1034 vp_p.n11944 vp_p.t1865 716.572
R1035 vp_p.n26148 vp_p.t2972 716.572
R1036 vp_p.n24722 vp_p.t2544 716.572
R1037 vp_p.n23300 vp_p.t2293 716.572
R1038 vp_p.n21877 vp_p.t1187 716.572
R1039 vp_p.n20453 vp_p.t1662 716.572
R1040 vp_p.n19028 vp_p.t526 716.572
R1041 vp_p.n17602 vp_p.t2374 716.572
R1042 vp_p.n16175 vp_p.t2531 716.572
R1043 vp_p.n14747 vp_p.t745 716.572
R1044 vp_p.n13583 vp_p.t1436 716.572
R1045 vp_p.n7942 vp_p.t2143 716.572
R1046 vp_p.n7940 vp_p.t1896 716.572
R1047 vp_p.n6518 vp_p.t1333 716.572
R1048 vp_p.n5095 vp_p.t1083 716.572
R1049 vp_p.n3671 vp_p.t2939 716.572
R1050 vp_p.n2246 vp_p.t2525 716.572
R1051 vp_p.n820 vp_p.t2268 716.572
R1052 vp_p.n9566 vp_p.t1164 716.572
R1053 vp_p.n11003 vp_p.t1625 716.572
R1054 vp_p.n12441 vp_p.t500 716.572
R1055 vp_p.n26644 vp_p.t909 716.572
R1056 vp_p.n25219 vp_p.t508 716.572
R1057 vp_p.n23797 vp_p.t247 716.572
R1058 vp_p.n22374 vp_p.t2125 716.572
R1059 vp_p.n20950 vp_p.t2578 716.572
R1060 vp_p.n19525 vp_p.t1467 716.572
R1061 vp_p.n18099 vp_p.t314 716.572
R1062 vp_p.n16672 vp_p.t1183 716.572
R1063 vp_p.n15244 vp_p.t1605 716.572
R1064 vp_p.n13578 vp_p.t74 716.572
R1065 vp_p.n7440 vp_p.t15 716.572
R1066 vp_p.n7438 vp_p.t2747 716.572
R1067 vp_p.n6016 vp_p.t1008 716.572
R1068 vp_p.n4593 vp_p.t755 716.572
R1069 vp_p.n3169 vp_p.t2607 716.572
R1070 vp_p.n1744 vp_p.t2195 716.572
R1071 vp_p.n260 vp_p.t1974 716.572
R1072 vp_p.n8999 vp_p.t827 716.572
R1073 vp_p.n10501 vp_p.t1309 716.572
R1074 vp_p.n11939 vp_p.t173 716.572
R1075 vp_p.n26143 vp_p.t1787 716.572
R1076 vp_p.n24717 vp_p.t1373 716.572
R1077 vp_p.n23295 vp_p.t1133 716.572
R1078 vp_p.n21872 vp_p.t2989 716.572
R1079 vp_p.n20448 vp_p.t470 716.572
R1080 vp_p.n19023 vp_p.t2318 716.572
R1081 vp_p.n17597 vp_p.t1201 716.572
R1082 vp_p.n16170 vp_p.t856 716.572
R1083 vp_p.n14742 vp_p.t2350 716.572
R1084 vp_p.n13573 vp_p.t2734 716.572
R1085 vp_p.n7956 vp_p.t1222 716.572
R1086 vp_p.n7954 vp_p.t967 716.572
R1087 vp_p.n6532 vp_p.t2658 716.572
R1088 vp_p.n5109 vp_p.t2404 716.572
R1089 vp_p.n3685 vp_p.t1289 716.572
R1090 vp_p.n2260 vp_p.t875 716.572
R1091 vp_p.n834 vp_p.t635 716.572
R1092 vp_p.n9580 vp_p.t2481 716.572
R1093 vp_p.n11017 vp_p.t2965 716.572
R1094 vp_p.n12455 vp_p.t1844 716.572
R1095 vp_p.n26658 vp_p.t2996 716.572
R1096 vp_p.n25233 vp_p.t2560 716.572
R1097 vp_p.n23811 vp_p.t2325 716.572
R1098 vp_p.n22388 vp_p.t1205 716.572
R1099 vp_p.n20964 vp_p.t1685 716.572
R1100 vp_p.n19539 vp_p.t546 716.572
R1101 vp_p.n18113 vp_p.t2387 716.572
R1102 vp_p.n16686 vp_p.t2514 716.572
R1103 vp_p.n15258 vp_p.t866 716.572
R1104 vp_p.n13568 vp_p.t1416 716.572
R1105 vp_p.n7435 vp_p.t1832 716.572
R1106 vp_p.n7433 vp_p.t1587 716.572
R1107 vp_p.n6011 vp_p.t2304 716.572
R1108 vp_p.n4588 vp_p.t2087 716.572
R1109 vp_p.n3164 vp_p.t934 716.572
R1110 vp_p.n1739 vp_p.t529 716.572
R1111 vp_p.n255 vp_p.t266 716.572
R1112 vp_p.n8994 vp_p.t2147 716.572
R1113 vp_p.n10496 vp_p.t2601 716.572
R1114 vp_p.n11934 vp_p.t1494 716.572
R1115 vp_p.n26138 vp_p.t608 716.572
R1116 vp_p.n24712 vp_p.t186 716.572
R1117 vp_p.n23290 vp_p.t2928 716.572
R1118 vp_p.n21867 vp_p.t1810 716.572
R1119 vp_p.n20443 vp_p.t2260 716.572
R1120 vp_p.n19018 vp_p.t1154 716.572
R1121 vp_p.n17592 vp_p.t9 716.572
R1122 vp_p.n16165 vp_p.t2166 716.572
R1123 vp_p.n14737 vp_p.t941 716.572
R1124 vp_p.n13563 vp_p.t1072 716.572
R1125 vp_p.n7970 vp_p.t34 716.572
R1126 vp_p.n7968 vp_p.t2770 716.572
R1127 vp_p.n6546 vp_p.t978 716.572
R1128 vp_p.n5123 vp_p.t733 716.572
R1129 vp_p.n3699 vp_p.t2584 716.572
R1130 vp_p.n2274 vp_p.t2180 716.572
R1131 vp_p.n848 vp_p.t1942 716.572
R1132 vp_p.n9594 vp_p.t796 716.572
R1133 vp_p.n11031 vp_p.t1286 716.572
R1134 vp_p.n12469 vp_p.t147 716.572
R1135 vp_p.n26672 vp_p.t1815 716.572
R1136 vp_p.n25247 vp_p.t1399 716.572
R1137 vp_p.n23825 vp_p.t1159 716.572
R1138 vp_p.n22402 vp_p.t12 716.572
R1139 vp_p.n20978 vp_p.t496 716.572
R1140 vp_p.n19553 vp_p.t2345 716.572
R1141 vp_p.n18127 vp_p.t1217 716.572
R1142 vp_p.n16700 vp_p.t833 716.572
R1143 vp_p.n15272 vp_p.t2447 716.572
R1144 vp_p.n13558 vp_p.t2710 716.572
R1145 vp_p.n7430 vp_p.t1658 716.572
R1146 vp_p.n7428 vp_p.t1411 716.572
R1147 vp_p.n6006 vp_p.t2870 716.572
R1148 vp_p.n4583 vp_p.t2623 716.572
R1149 vp_p.n3159 vp_p.t1513 716.572
R1150 vp_p.n1734 vp_p.t1085 716.572
R1151 vp_p.n250 vp_p.t845 716.572
R1152 vp_p.n8989 vp_p.t2695 716.572
R1153 vp_p.n10491 vp_p.t190 716.572
R1154 vp_p.n11929 vp_p.t2060 716.572
R1155 vp_p.n26133 vp_p.t416 716.572
R1156 vp_p.n24707 vp_p.t14 716.572
R1157 vp_p.n23285 vp_p.t2746 716.572
R1158 vp_p.n21862 vp_p.t1631 716.572
R1159 vp_p.n20438 vp_p.t2112 716.572
R1160 vp_p.n19013 vp_p.t964 716.572
R1161 vp_p.n17587 vp_p.t2820 716.572
R1162 vp_p.n16160 vp_p.t2712 716.572
R1163 vp_p.n14732 vp_p.t325 716.572
R1164 vp_p.n13553 vp_p.t1633 716.572
R1165 vp_p.n7984 vp_p.t1512 716.572
R1166 vp_p.n7982 vp_p.t1260 716.572
R1167 vp_p.n6560 vp_p.t303 716.572
R1168 vp_p.n5137 vp_p.t71 716.572
R1169 vp_p.n3713 vp_p.t1936 716.572
R1170 vp_p.n2288 vp_p.t1531 716.572
R1171 vp_p.n862 vp_p.t1278 716.572
R1172 vp_p.n9608 vp_p.t139 716.572
R1173 vp_p.n11045 vp_p.t629 716.572
R1174 vp_p.n12483 vp_p.t2474 716.572
R1175 vp_p.n26686 vp_p.t263 716.572
R1176 vp_p.n25261 vp_p.t2842 716.572
R1177 vp_p.n23839 vp_p.t2598 716.572
R1178 vp_p.n22416 vp_p.t1490 716.572
R1179 vp_p.n20992 vp_p.t1966 716.572
R1180 vp_p.n19567 vp_p.t818 716.572
R1181 vp_p.n18141 vp_p.t2675 716.572
R1182 vp_p.n16714 vp_p.t168 716.572
R1183 vp_p.n15286 vp_p.t289 716.572
R1184 vp_p.n13548 vp_p.t2074 716.572
R1185 vp_p.n7425 vp_p.t2697 716.572
R1186 vp_p.n7423 vp_p.t2458 716.572
R1187 vp_p.n6001 vp_p.t1988 716.572
R1188 vp_p.n4578 vp_p.t1741 716.572
R1189 vp_p.n3154 vp_p.t607 716.572
R1190 vp_p.n1729 vp_p.t185 716.572
R1191 vp_p.n245 vp_p.t2927 716.572
R1192 vp_p.n8984 vp_p.t1809 716.572
R1193 vp_p.n10486 vp_p.t2259 716.572
R1194 vp_p.n11924 vp_p.t1152 716.572
R1195 vp_p.n26128 vp_p.t1496 716.572
R1196 vp_p.n24702 vp_p.t1073 716.572
R1197 vp_p.n23280 vp_p.t825 716.572
R1198 vp_p.n21857 vp_p.t2678 716.572
R1199 vp_p.n20433 vp_p.t172 716.572
R1200 vp_p.n19008 vp_p.t2045 716.572
R1201 vp_p.n17582 vp_p.t893 716.572
R1202 vp_p.n16155 vp_p.t1839 716.572
R1203 vp_p.n14727 vp_p.t1819 716.572
R1204 vp_p.n13543 vp_p.t724 716.572
R1205 vp_p.n7998 vp_p.t1344 716.572
R1206 vp_p.n7996 vp_p.t1087 716.572
R1207 vp_p.n6574 vp_p.t883 716.572
R1208 vp_p.n5151 vp_p.t647 716.572
R1209 vp_p.n3727 vp_p.t2492 716.572
R1210 vp_p.n2302 vp_p.t2094 716.572
R1211 vp_p.n876 vp_p.t1851 716.572
R1212 vp_p.n9622 vp_p.t706 716.572
R1213 vp_p.n11059 vp_p.t1189 716.572
R1214 vp_p.n12497 vp_p.t42 716.572
R1215 vp_p.n26700 vp_p.t98 716.572
R1216 vp_p.n25275 vp_p.t2682 716.572
R1217 vp_p.n23853 vp_p.t2430 716.572
R1218 vp_p.n22430 vp_p.t1319 716.572
R1219 vp_p.n21006 vp_p.t1794 716.572
R1220 vp_p.n19581 vp_p.t664 716.572
R1221 vp_p.n18155 vp_p.t2513 716.572
R1222 vp_p.n16728 vp_p.t726 716.572
R1223 vp_p.n15300 vp_p.t2672 716.572
R1224 vp_p.n13538 vp_p.t2610 716.572
R1225 vp_p.n7420 vp_p.t1535 716.572
R1226 vp_p.n7418 vp_p.t1280 716.572
R1227 vp_p.n5996 vp_p.t277 716.572
R1228 vp_p.n4573 vp_p.t49 716.572
R1229 vp_p.n3149 vp_p.t1911 716.572
R1230 vp_p.n1724 vp_p.t1504 716.572
R1231 vp_p.n240 vp_p.t1254 716.572
R1232 vp_p.n8979 vp_p.t108 716.572
R1233 vp_p.n10481 vp_p.t606 716.572
R1234 vp_p.n11919 vp_p.t2446 716.572
R1235 vp_p.n26123 vp_p.t284 716.572
R1236 vp_p.n24697 vp_p.t2869 716.572
R1237 vp_p.n23275 vp_p.t2620 716.572
R1238 vp_p.n21852 vp_p.t1510 716.572
R1239 vp_p.n20428 vp_p.t1991 716.572
R1240 vp_p.n19003 vp_p.t844 716.572
R1241 vp_p.n17577 vp_p.t2693 716.572
R1242 vp_p.n16150 vp_p.t141 716.572
R1243 vp_p.n14722 vp_p.t402 716.572
R1244 vp_p.n13533 vp_p.t2054 716.572
R1245 vp_p.n8012 vp_p.t146 716.572
R1246 vp_p.n8010 vp_p.t2889 716.572
R1247 vp_p.n6588 vp_p.t2187 716.572
R1248 vp_p.n5165 vp_p.t1957 716.572
R1249 vp_p.n3741 vp_p.t812 716.572
R1250 vp_p.n2316 vp_p.t392 716.572
R1251 vp_p.n890 vp_p.t157 716.572
R1252 vp_p.n9636 vp_p.t2037 716.572
R1253 vp_p.n11073 vp_p.t2485 716.572
R1254 vp_p.n12511 vp_p.t1365 716.572
R1255 vp_p.n26714 vp_p.t1920 716.572
R1256 vp_p.n25289 vp_p.t1516 716.572
R1257 vp_p.n23867 vp_p.t1262 716.572
R1258 vp_p.n22444 vp_p.t122 716.572
R1259 vp_p.n21020 vp_p.t612 716.572
R1260 vp_p.n19595 vp_p.t2455 716.572
R1261 vp_p.n18169 vp_p.t1339 716.572
R1262 vp_p.n16742 vp_p.t2055 716.572
R1263 vp_p.n15314 vp_p.t1285 716.572
R1264 vp_p.n13528 vp_p.t935 716.572
R1265 vp_p.n7415 vp_p.t70 716.572
R1266 vp_p.n7413 vp_p.t2811 716.572
R1267 vp_p.n5991 vp_p.t1204 716.572
R1268 vp_p.n4568 vp_p.t940 716.572
R1269 vp_p.n3144 vp_p.t2798 716.572
R1270 vp_p.n1719 vp_p.t2384 716.572
R1271 vp_p.n235 vp_p.t2158 716.572
R1272 vp_p.n8974 vp_p.t1023 716.572
R1273 vp_p.n10476 vp_p.t1502 716.572
R1274 vp_p.n11914 vp_p.t358 716.572
R1275 vp_p.n26118 vp_p.t1859 716.572
R1276 vp_p.n24692 vp_p.t1428 716.572
R1277 vp_p.n23270 vp_p.t1198 716.572
R1278 vp_p.n21847 vp_p.t48 716.572
R1279 vp_p.n20423 vp_p.t533 716.572
R1280 vp_p.n18998 vp_p.t2380 716.572
R1281 vp_p.n17572 vp_p.t1253 716.572
R1282 vp_p.n16145 vp_p.t1051 716.572
R1283 vp_p.n14717 vp_p.t1774 716.572
R1284 vp_p.n13523 vp_p.t2935 716.572
R1285 vp_p.n8026 vp_p.t2906 716.572
R1286 vp_p.n8024 vp_p.t2670 716.572
R1287 vp_p.n6602 vp_p.t1626 716.572
R1288 vp_p.n5179 vp_p.t1393 716.572
R1289 vp_p.n3755 vp_p.t237 716.572
R1290 vp_p.n2330 vp_p.t2813 716.572
R1291 vp_p.n904 vp_p.t2568 716.572
R1292 vp_p.n9650 vp_p.t1453 716.572
R1293 vp_p.n11087 vp_p.t1926 716.572
R1294 vp_p.n12525 vp_p.t784 716.572
R1295 vp_p.n26728 vp_p.t1716 716.572
R1296 vp_p.n25303 vp_p.t1281 716.572
R1297 vp_p.n23881 vp_p.t1047 716.572
R1298 vp_p.n22458 vp_p.t2887 716.572
R1299 vp_p.n21034 vp_p.t378 716.572
R1300 vp_p.n19609 vp_p.t2225 716.572
R1301 vp_p.n18183 vp_p.t1106 716.572
R1302 vp_p.n16756 vp_p.t1485 716.572
R1303 vp_p.n15328 vp_p.t1750 716.572
R1304 vp_p.n13518 vp_p.t375 716.572
R1305 vp_p.n7410 vp_p.t1551 716.572
R1306 vp_p.n7408 vp_p.t1301 716.572
R1307 vp_p.n5986 vp_p.t534 716.572
R1308 vp_p.n4563 vp_p.t272 716.572
R1309 vp_p.n3139 vp_p.t2151 716.572
R1310 vp_p.n1714 vp_p.t1737 716.572
R1311 vp_p.n230 vp_p.t1497 716.572
R1312 vp_p.n8969 vp_p.t350 716.572
R1313 vp_p.n10471 vp_p.t829 716.572
R1314 vp_p.n11909 vp_p.t2681 716.572
R1315 vp_p.n26113 vp_p.t309 716.572
R1316 vp_p.n24687 vp_p.t2888 716.572
R1317 vp_p.n23265 vp_p.t2649 716.572
R1318 vp_p.n21842 vp_p.t1534 716.572
R1319 vp_p.n20418 vp_p.t2014 716.572
R1320 vp_p.n18993 vp_p.t869 716.572
R1321 vp_p.n17567 vp_p.t2706 716.572
R1322 vp_p.n16140 vp_p.t377 716.572
R1323 vp_p.n14712 vp_p.t2597 716.572
R1324 vp_p.n13513 vp_p.t2258 716.572
R1325 vp_p.n8040 vp_p.t2730 716.572
R1326 vp_p.n8038 vp_p.t2501 716.572
R1327 vp_p.n6616 vp_p.t2183 716.572
R1328 vp_p.n5193 vp_p.t1948 716.572
R1329 vp_p.n3769 vp_p.t802 716.572
R1330 vp_p.n2344 vp_p.t388 716.572
R1331 vp_p.n918 vp_p.t153 716.572
R1332 vp_p.n9664 vp_p.t2031 716.572
R1333 vp_p.n11101 vp_p.t2480 716.572
R1334 vp_p.n12539 vp_p.t1363 716.572
R1335 vp_p.n26742 vp_p.t1537 716.572
R1336 vp_p.n25317 vp_p.t1110 716.572
R1337 vp_p.n23895 vp_p.t871 716.572
R1338 vp_p.n22472 vp_p.t2708 716.572
R1339 vp_p.n21048 vp_p.t211 716.572
R1340 vp_p.n19623 vp_p.t2078 716.572
R1341 vp_p.n18197 vp_p.t926 716.572
R1342 vp_p.n16770 vp_p.t2051 716.572
R1343 vp_p.n15342 vp_p.t1125 716.572
R1344 vp_p.n13508 vp_p.t929 716.572
R1345 vp_p.n7405 vp_p.t354 716.572
R1346 vp_p.n7403 vp_p.t101 716.572
R1347 vp_p.n5981 vp_p.t1858 716.572
R1348 vp_p.n4558 vp_p.t1604 716.572
R1349 vp_p.n3134 vp_p.t469 716.572
R1350 vp_p.n1709 vp_p.t47 716.572
R1351 vp_p.n225 vp_p.t2789 716.572
R1352 vp_p.n8964 vp_p.t1675 716.572
R1353 vp_p.n10466 vp_p.t2146 716.572
R1354 vp_p.n11904 vp_p.t1015 716.572
R1355 vp_p.n26108 vp_p.t2134 716.572
R1356 vp_p.n24682 vp_p.t1726 716.572
R1357 vp_p.n23260 vp_p.t1479 716.572
R1358 vp_p.n21837 vp_p.t331 716.572
R1359 vp_p.n20413 vp_p.t805 716.572
R1360 vp_p.n18988 vp_p.t2665 716.572
R1361 vp_p.n17562 vp_p.t1547 716.572
R1362 vp_p.n16135 vp_p.t1707 716.572
R1363 vp_p.n14707 vp_p.t1219 716.572
R1364 vp_p.n13503 vp_p.t602 716.572
R1365 vp_p.n8054 vp_p.t1571 716.572
R1366 vp_p.n8052 vp_p.t1325 716.572
R1367 vp_p.n6630 vp_p.t515 716.572
R1368 vp_p.n5207 vp_p.t250 716.572
R1369 vp_p.n3783 vp_p.t2128 716.572
R1370 vp_p.n2358 vp_p.t1724 716.572
R1371 vp_p.n932 vp_p.t1473 716.572
R1372 vp_p.n9678 vp_p.t323 716.572
R1373 vp_p.n11115 vp_p.t798 716.572
R1374 vp_p.n12553 vp_p.t2661 716.572
R1375 vp_p.n26756 vp_p.t339 716.572
R1376 vp_p.n25331 vp_p.t2905 716.572
R1377 vp_p.n23909 vp_p.t2669 716.572
R1378 vp_p.n22486 vp_p.t1550 716.572
R1379 vp_p.n21062 vp_p.t2036 716.572
R1380 vp_p.n19637 vp_p.t885 716.572
R1381 vp_p.n18211 vp_p.t2725 716.572
R1382 vp_p.n16784 vp_p.t353 716.572
R1383 vp_p.n15356 vp_p.t2703 716.572
R1384 vp_p.n13498 vp_p.t2235 716.572
R1385 vp_p.n7400 vp_p.t2415 716.572
R1386 vp_p.n7398 vp_p.t2179 716.572
R1387 vp_p.n5976 vp_p.t189 716.572
R1388 vp_p.n4553 vp_p.t2932 716.572
R1389 vp_p.n3129 vp_p.t1814 716.572
R1390 vp_p.n1704 vp_p.t1398 716.572
R1391 vp_p.n220 vp_p.t1158 716.572
R1392 vp_p.n8959 vp_p.t11 716.572
R1393 vp_p.n10461 vp_p.t495 716.572
R1394 vp_p.n11899 vp_p.t2344 716.572
R1395 vp_p.n26103 vp_p.t1214 716.572
R1396 vp_p.n24677 vp_p.t783 716.572
R1397 vp_p.n23255 vp_p.t554 716.572
R1398 vp_p.n21832 vp_p.t2395 716.572
R1399 vp_p.n20408 vp_p.t2873 716.572
R1400 vp_p.n18983 vp_p.t1753 716.572
R1401 vp_p.n17557 vp_p.t626 716.572
R1402 vp_p.n16130 vp_p.t37 716.572
R1403 vp_p.n14702 vp_p.t478 716.572
R1404 vp_p.n13493 vp_p.t1932 716.572
R1405 vp_p.n8068 vp_p.t374 716.572
R1406 vp_p.n8066 vp_p.t125 716.572
R1407 vp_p.n6644 vp_p.t1831 716.572
R1408 vp_p.n5221 vp_p.t1586 716.572
R1409 vp_p.n3797 vp_p.t441 716.572
R1410 vp_p.n2372 vp_p.t30 716.572
R1411 vp_p.n946 vp_p.t2763 716.572
R1412 vp_p.n9692 vp_p.t1649 716.572
R1413 vp_p.n11129 vp_p.t2127 716.572
R1414 vp_p.n12567 vp_p.t985 716.572
R1415 vp_p.n26770 vp_p.t2154 716.572
R1416 vp_p.n25345 vp_p.t1740 716.572
R1417 vp_p.n23923 vp_p.t1498 716.572
R1418 vp_p.n22500 vp_p.t352 716.572
R1419 vp_p.n21076 vp_p.t832 716.572
R1420 vp_p.n19651 vp_p.t2683 716.572
R1421 vp_p.n18225 vp_p.t1567 716.572
R1422 vp_p.n16798 vp_p.t1681 716.572
R1423 vp_p.n15370 vp_p.t1328 716.572
R1424 vp_p.n13488 vp_p.t583 716.572
R1425 vp_p.n7395 vp_p.t1244 716.572
R1426 vp_p.n7393 vp_p.t1001 716.572
R1427 vp_p.n5971 vp_p.t1509 716.572
R1428 vp_p.n4548 vp_p.t1256 716.572
R1429 vp_p.n3124 vp_p.t112 716.572
R1430 vp_p.n1699 vp_p.t2691 716.572
R1431 vp_p.n215 vp_p.t2448 716.572
R1432 vp_p.n8954 vp_p.t1332 716.572
R1433 vp_p.n10456 vp_p.t1808 716.572
R1434 vp_p.n11894 vp_p.t678 716.572
R1435 vp_p.n26098 vp_p.t24 716.572
R1436 vp_p.n24672 vp_p.t2583 716.572
R1437 vp_p.n23250 vp_p.t2354 716.572
R1438 vp_p.n21827 vp_p.t1226 716.572
R1439 vp_p.n20403 vp_p.t1718 716.572
R1440 vp_p.n18978 vp_p.t571 716.572
R1441 vp_p.n17552 vp_p.t2406 716.572
R1442 vp_p.n16125 vp_p.t1359 716.572
R1443 vp_p.n14697 vp_p.t2080 716.572
R1444 vp_p.n13483 vp_p.t242 716.572
R1445 vp_p.n8082 vp_p.t2178 716.572
R1446 vp_p.n8080 vp_p.t1943 716.572
R1447 vp_p.n6658 vp_p.t135 716.572
R1448 vp_p.n5235 vp_p.t2879 716.572
R1449 vp_p.n3811 vp_p.t1760 716.572
R1450 vp_p.n2386 vp_p.t1353 716.572
R1451 vp_p.n960 vp_p.t1097 716.572
R1452 vp_p.n9706 vp_p.t2960 716.572
R1453 vp_p.n11143 vp_p.t429 716.572
R1454 vp_p.n12581 vp_p.t2284 716.572
R1455 vp_p.n26784 vp_p.t955 716.572
R1456 vp_p.n25359 vp_p.t553 716.572
R1457 vp_p.n23937 vp_p.t287 716.572
R1458 vp_p.n22514 vp_p.t2165 716.572
R1459 vp_p.n21090 vp_p.t2628 716.572
R1460 vp_p.n19665 vp_p.t1517 716.572
R1461 vp_p.n18239 vp_p.t367 716.572
R1462 vp_p.n16812 vp_p.t2986 716.572
R1463 vp_p.n15384 vp_p.t2900 716.572
R1464 vp_p.n13478 vp_p.t1889 716.572
R1465 vp_p.n7390 vp_p.t58 716.572
R1466 vp_p.n7388 vp_p.t2795 716.572
R1467 vp_p.n5966 vp_p.t2799 716.572
R1468 vp_p.n4543 vp_p.t2555 716.572
R1469 vp_p.n3119 vp_p.t1435 716.572
R1470 vp_p.n1694 vp_p.t1026 716.572
R1471 vp_p.n210 vp_p.t767 716.572
R1472 vp_p.n8949 vp_p.t2626 716.572
R1473 vp_p.n10451 vp_p.t107 716.572
R1474 vp_p.n11889 vp_p.t1993 716.572
R1475 vp_p.n26093 vp_p.t1843 716.572
R1476 vp_p.n24667 vp_p.t1415 716.572
R1477 vp_p.n23245 vp_p.t1180 716.572
R1478 vp_p.n21822 vp_p.t39 716.572
R1479 vp_p.n20398 vp_p.t523 716.572
R1480 vp_p.n18973 vp_p.t2369 716.572
R1481 vp_p.n17547 vp_p.t1239 716.572
R1482 vp_p.n16120 vp_p.t2657 716.572
R1483 vp_p.n14692 vp_p.t682 716.572
R1484 vp_p.n13473 vp_p.t1574 716.572
R1485 vp_p.n8096 vp_p.t917 716.572
R1486 vp_p.n8094 vp_p.t687 716.572
R1487 vp_p.n6672 vp_p.t2486 716.572
R1488 vp_p.n5249 vp_p.t2231 716.572
R1489 vp_p.n3825 vp_p.t1120 716.572
R1490 vp_p.n2400 vp_p.t703 716.572
R1491 vp_p.n974 vp_p.t456 716.572
R1492 vp_p.n9720 vp_p.t2302 716.572
R1493 vp_p.n11157 vp_p.t2781 716.572
R1494 vp_p.n12595 vp_p.t1667 716.572
R1495 vp_p.n26798 vp_p.t2689 716.572
R1496 vp_p.n25373 vp_p.t2265 716.572
R1497 vp_p.n23951 vp_p.t2053 716.572
R1498 vp_p.n22528 vp_p.t901 716.572
R1499 vp_p.n21104 vp_p.t1389 716.572
R1500 vp_p.n19679 vp_p.t236 716.572
R1501 vp_p.n18253 vp_p.t2111 716.572
R1502 vp_p.n16826 vp_p.t2339 716.572
R1503 vp_p.n15398 vp_p.t1425 716.572
R1504 vp_p.n13468 vp_p.t1243 716.572
R1505 vp_p.n7385 vp_p.t1875 716.572
R1506 vp_p.n7383 vp_p.t1621 716.572
R1507 vp_p.n5961 vp_p.t1139 716.572
R1508 vp_p.n4538 vp_p.t889 716.572
R1509 vp_p.n3114 vp_p.t2733 716.572
R1510 vp_p.n1689 vp_p.t2328 716.572
R1511 vp_p.n205 vp_p.t2100 716.572
R1512 vp_p.n8944 vp_p.t948 716.572
R1513 vp_p.n10446 vp_p.t1433 716.572
R1514 vp_p.n11884 vp_p.t283 716.572
R1515 vp_p.n26088 vp_p.t654 716.572
R1516 vp_p.n24662 vp_p.t223 716.572
R1517 vp_p.n23240 vp_p.t2982 716.572
R1518 vp_p.n21817 vp_p.t1861 716.572
R1519 vp_p.n20393 vp_p.t2312 716.572
R1520 vp_p.n18968 vp_p.t1199 716.572
R1521 vp_p.n17542 vp_p.t51 716.572
R1522 vp_p.n16115 vp_p.t975 716.572
R1523 vp_p.n14687 vp_p.t2249 716.572
R1524 vp_p.n13463 vp_p.t2868 716.572
R1525 vp_p.n8110 vp_p.t2716 716.572
R1526 vp_p.n8108 vp_p.t2482 716.572
R1527 vp_p.n6686 vp_p.t804 716.572
R1528 vp_p.n5263 vp_p.t576 716.572
R1529 vp_p.n3839 vp_p.t2414 716.572
R1530 vp_p.n2414 vp_p.t2033 716.572
R1531 vp_p.n988 vp_p.t1778 716.572
R1532 vp_p.n9734 vp_p.t646 716.572
R1533 vp_p.n11171 vp_p.t1115 716.572
R1534 vp_p.n12609 vp_p.t2973 716.572
R1535 vp_p.n26812 vp_p.t1520 716.572
R1536 vp_p.n25387 vp_p.t1093 716.572
R1537 vp_p.n23965 vp_p.t855 716.572
R1538 vp_p.n22542 vp_p.t2700 716.572
R1539 vp_p.n21118 vp_p.t199 716.572
R1540 vp_p.n19693 vp_p.t2068 716.572
R1541 vp_p.n18267 vp_p.t913 716.572
R1542 vp_p.n16840 vp_p.t676 716.572
R1543 vp_p.n15412 vp_p.t27 716.572
R1544 vp_p.n13458 vp_p.t2546 716.572
R1545 vp_p.n7380 vp_p.t1714 716.572
R1546 vp_p.n7378 vp_p.t1459 716.572
R1547 vp_p.n5956 vp_p.t1715 716.572
R1548 vp_p.n4533 vp_p.t1460 716.572
R1549 vp_p.n3109 vp_p.t308 716.572
R1550 vp_p.n1684 vp_p.t2886 716.572
R1551 vp_p.n200 vp_p.t2645 716.572
R1552 vp_p.n8939 vp_p.t1530 716.572
R1553 vp_p.n10441 vp_p.t2010 716.572
R1554 vp_p.n11879 vp_p.t865 716.572
R1555 vp_p.n26083 vp_p.t479 716.572
R1556 vp_p.n24657 vp_p.t57 716.572
R1557 vp_p.n23235 vp_p.t2794 716.572
R1558 vp_p.n21812 vp_p.t1686 716.572
R1559 vp_p.n20388 vp_p.t2157 716.572
R1560 vp_p.n18963 vp_p.t1022 716.572
R1561 vp_p.n17537 vp_p.t2866 716.572
R1562 vp_p.n16110 vp_p.t1554 716.572
R1563 vp_p.n14682 vp_p.t1654 716.572
R1564 vp_p.n13453 vp_p.t443 716.572
R1565 vp_p.n8124 vp_p.t1556 716.572
R1566 vp_p.n8122 vp_p.t1308 716.572
R1567 vp_p.n6700 vp_p.t2132 716.572
R1568 vp_p.n5277 vp_p.t1886 716.572
R1569 vp_p.n3853 vp_p.t738 716.572
R1570 vp_p.n2428 vp_p.t324 716.572
R1571 vp_p.n1002 vp_p.t81 716.572
R1572 vp_p.n9748 vp_p.t1956 716.572
R1573 vp_p.n11185 vp_p.t2410 716.572
R1574 vp_p.n12623 vp_p.t1294 716.572
R1575 vp_p.n26826 vp_p.t313 716.572
R1576 vp_p.n25401 vp_p.t2893 716.572
R1577 vp_p.n23979 vp_p.t2654 716.572
R1578 vp_p.n22556 vp_p.t1540 716.572
R1579 vp_p.n21132 vp_p.t2020 716.572
R1580 vp_p.n19707 vp_p.t874 716.572
R1581 vp_p.n18281 vp_p.t2711 716.572
R1582 vp_p.n16854 vp_p.t1987 716.572
R1583 vp_p.n15426 vp_p.t1620 716.572
R1584 vp_p.n13448 vp_p.t881 716.572
R1585 vp_p.n7375 vp_p.t2736 716.572
R1586 vp_p.n7373 vp_p.t2506 716.572
R1587 vp_p.n5951 vp_p.t780 716.572
R1588 vp_p.n4528 vp_p.t552 716.572
R1589 vp_p.n3104 vp_p.t2394 716.572
R1590 vp_p.n1679 vp_p.t2006 716.572
R1591 vp_p.n195 vp_p.t1752 716.572
R1592 vp_p.n8934 vp_p.t625 716.572
R1593 vp_p.n10436 vp_p.t1088 716.572
R1594 vp_p.n11874 vp_p.t2949 716.572
R1595 vp_p.n26078 vp_p.t1543 716.572
R1596 vp_p.n24652 vp_p.t1119 716.572
R1597 vp_p.n23230 vp_p.t877 716.572
R1598 vp_p.n21807 vp_p.t2714 716.572
R1599 vp_p.n20383 vp_p.t216 716.572
R1600 vp_p.n18958 vp_p.t2085 716.572
R1601 vp_p.n17532 vp_p.t931 716.572
R1602 vp_p.n16105 vp_p.t651 716.572
R1603 vp_p.n14677 vp_p.t123 716.572
R1604 vp_p.n13443 vp_p.t2530 716.572
R1605 vp_p.n8138 vp_p.t1388 716.572
R1606 vp_p.n8136 vp_p.t1144 716.572
R1607 vp_p.n6714 vp_p.t2679 716.572
R1608 vp_p.n5291 vp_p.t2429 716.572
R1609 vp_p.n3867 vp_p.t1318 716.572
R1610 vp_p.n2442 vp_p.t894 716.572
R1611 vp_p.n1016 vp_p.t660 716.572
R1612 vp_p.n9762 vp_p.t2512 716.572
R1613 vp_p.n11199 vp_p.t2992 716.572
R1614 vp_p.n12637 vp_p.t1866 716.572
R1615 vp_p.n26840 vp_p.t156 716.572
R1616 vp_p.n25415 vp_p.t2719 716.572
R1617 vp_p.n23993 vp_p.t2484 716.572
R1618 vp_p.n22570 vp_p.t1364 716.572
R1619 vp_p.n21146 vp_p.t1847 716.572
R1620 vp_p.n19721 vp_p.t701 716.572
R1621 vp_p.n18295 vp_p.t2547 716.572
R1622 vp_p.n16868 vp_p.t2534 716.572
R1623 vp_p.n15440 vp_p.t996 716.572
R1624 vp_p.n13438 vp_p.t1438 716.572
R1625 vp_p.n7370 vp_p.t1233 716.572
R1626 vp_p.n7368 vp_p.t984 716.572
R1627 vp_p.n5946 vp_p.t117 716.572
R1628 vp_p.n4523 vp_p.t2865 716.572
R1629 vp_p.n3099 vp_p.t1748 716.572
R1630 vp_p.n1674 vp_p.t1338 716.572
R1631 vp_p.n190 vp_p.t1082 716.572
R1632 vp_p.n8929 vp_p.t2938 716.572
R1633 vp_p.n10431 vp_p.t412 716.572
R1634 vp_p.n11869 vp_p.t2267 716.572
R1635 vp_p.n26073 vp_p.t8 716.572
R1636 vp_p.n24647 vp_p.t2571 716.572
R1637 vp_p.n23225 vp_p.t2342 716.572
R1638 vp_p.n21802 vp_p.t1215 716.572
R1639 vp_p.n20378 vp_p.t1696 716.572
R1640 vp_p.n18953 vp_p.t558 716.572
R1641 vp_p.n17527 vp_p.t2397 716.572
R1642 vp_p.n16100 vp_p.t2969 716.572
R1643 vp_p.n14672 vp_p.t966 716.572
R1644 vp_p.n13433 vp_p.t1879 716.572
R1645 vp_p.n8152 vp_p.t198 716.572
R1646 vp_p.n8150 vp_p.t2941 716.572
R1647 vp_p.n6728 vp_p.t1011 716.572
R1648 vp_p.n5305 vp_p.t756 716.572
R1649 vp_p.n3881 vp_p.t2609 716.572
R1650 vp_p.n2456 vp_p.t2198 716.572
R1651 vp_p.n1030 vp_p.t1978 716.572
R1652 vp_p.n9776 vp_p.t831 716.572
R1653 vp_p.n11213 vp_p.t1314 716.572
R1654 vp_p.n12651 vp_p.t176 716.572
R1655 vp_p.n26854 vp_p.t1977 716.572
R1656 vp_p.n25429 vp_p.t1560 716.572
R1657 vp_p.n24007 vp_p.t1312 716.572
R1658 vp_p.n22584 vp_p.t175 716.572
R1659 vp_p.n21160 vp_p.t656 716.572
R1660 vp_p.n19735 vp_p.t2504 716.572
R1661 vp_p.n18309 vp_p.t1383 716.572
R1662 vp_p.n16882 vp_p.t857 716.572
R1663 vp_p.n15454 vp_p.t2577 716.572
R1664 vp_p.n13428 vp_p.t2735 716.572
R1665 vp_p.n7365 vp_p.t1066 716.572
R1666 vp_p.n7363 vp_p.t813 716.572
R1667 vp_p.n5941 vp_p.t693 716.572
R1668 vp_p.n4518 vp_p.t440 716.572
R1669 vp_p.n3094 vp_p.t2290 716.572
R1670 vp_p.n1669 vp_p.t1894 716.572
R1671 vp_p.n185 vp_p.t1653 716.572
R1672 vp_p.n8924 vp_p.t522 716.572
R1673 vp_p.n10426 vp_p.t983 716.572
R1674 vp_p.n11864 vp_p.t2832 716.572
R1675 vp_p.n26068 vp_p.t2819 716.572
R1676 vp_p.n24642 vp_p.t2401 716.572
R1677 vp_p.n23220 vp_p.t2170 716.572
R1678 vp_p.n21797 vp_p.t1048 716.572
R1679 vp_p.n20373 vp_p.t1526 716.572
R1680 vp_p.n18948 vp_p.t382 716.572
R1681 vp_p.n17522 vp_p.t2226 716.572
R1682 vp_p.n16095 vp_p.t542 716.572
R1683 vp_p.n14667 vp_p.t348 716.572
R1684 vp_p.n13423 vp_p.t2418 716.572
R1685 vp_p.n8166 vp_p.t1249 716.572
R1686 vp_p.n8164 vp_p.t1010 716.572
R1687 vp_p.n6742 vp_p.t92 716.572
R1688 vp_p.n5319 vp_p.t2840 716.572
R1689 vp_p.n3895 vp_p.t1732 716.572
R1690 vp_p.n2470 vp_p.t1307 716.572
R1691 vp_p.n1044 vp_p.t1068 716.572
R1692 vp_p.n9790 vp_p.t2912 716.572
R1693 vp_p.n11227 vp_p.t395 716.572
R1694 vp_p.n12665 vp_p.t2245 716.572
R1695 vp_p.n26868 vp_p.t29 716.572
R1696 vp_p.n25443 vp_p.t2591 716.572
R1697 vp_p.n24021 vp_p.t2362 716.572
R1698 vp_p.n22598 vp_p.t1230 716.572
R1699 vp_p.n21174 vp_p.t1721 716.572
R1700 vp_p.n19749 vp_p.t582 716.572
R1701 vp_p.n18323 vp_p.t2417 716.572
R1702 vp_p.n16896 vp_p.t2944 716.572
R1703 vp_p.n15468 vp_p.t1076 716.572
R1704 vp_p.n13418 vp_p.t1862 716.572
R1705 vp_p.n7360 vp_p.t2854 716.572
R1706 vp_p.n7358 vp_p.t2611 716.572
R1707 vp_p.n5936 vp_p.t2019 716.572
R1708 vp_p.n4513 vp_p.t1759 716.572
R1709 vp_p.n3089 vp_p.t632 716.572
R1710 vp_p.n1664 vp_p.t210 716.572
R1711 vp_p.n180 vp_p.t2959 716.572
R1712 vp_p.n8919 vp_p.t1837 716.572
R1713 vp_p.n10421 vp_p.t2283 716.572
R1714 vp_p.n11859 vp_p.t1177 716.572
R1715 vp_p.n26063 vp_p.t1652 716.572
R1716 vp_p.n24637 vp_p.t1232 716.572
R1717 vp_p.n23215 vp_p.t987 716.572
R1718 vp_p.n21792 vp_p.t2833 716.572
R1719 vp_p.n20368 vp_p.t320 716.572
R1720 vp_p.n18943 vp_p.t2185 716.572
R1721 vp_p.n17517 vp_p.t1060 716.572
R1722 vp_p.n16090 vp_p.t1863 716.572
R1723 vp_p.n14662 vp_p.t1949 716.572
R1724 vp_p.n13413 vp_p.t741 716.572
R1725 vp_p.n8180 vp_p.t2778 716.572
R1726 vp_p.n8178 vp_p.t2537 716.572
R1727 vp_p.n6756 vp_p.t1002 716.572
R1728 vp_p.n5333 vp_p.t748 716.572
R1729 vp_p.n3909 vp_p.t2602 716.572
R1730 vp_p.n2484 vp_p.t2193 716.572
R1731 vp_p.n1058 vp_p.t1973 716.572
R1732 vp_p.n9804 vp_p.t824 716.572
R1733 vp_p.n11241 vp_p.t1306 716.572
R1734 vp_p.n12679 vp_p.t169 716.572
R1735 vp_p.n26882 vp_p.t1580 716.572
R1736 vp_p.n25457 vp_p.t1167 716.572
R1737 vp_p.n24035 vp_p.t904 716.572
R1738 vp_p.n22612 vp_p.t2755 716.572
R1739 vp_p.n21188 vp_p.t245 716.572
R1740 vp_p.n19763 vp_p.t2119 716.572
R1741 vp_p.n18337 vp_p.t972 716.572
R1742 vp_p.n16910 vp_p.t853 716.572
R1743 vp_p.n15482 vp_p.t2421 716.572
R1744 vp_p.n13408 vp_p.t2729 716.572
R1745 vp_p.n7355 vp_p.t394 716.572
R1746 vp_p.n7353 vp_p.t161 716.572
R1747 vp_p.n5931 vp_p.t668 716.572
R1748 vp_p.n4508 vp_p.t405 716.572
R1749 vp_p.n3084 vp_p.t2257 716.572
R1750 vp_p.n1659 vp_p.t1869 716.572
R1751 vp_p.n175 vp_p.t1617 716.572
R1752 vp_p.n8914 vp_p.t490 716.572
R1753 vp_p.n10416 vp_p.t947 716.572
R1754 vp_p.n11854 vp_p.t2805 716.572
R1755 vp_p.n26058 vp_p.t2172 716.572
R1756 vp_p.n24632 vp_p.t1762 716.572
R1757 vp_p.n23210 vp_p.t1525 716.572
R1758 vp_p.n21787 vp_p.t381 716.572
R1759 vp_p.n20363 vp_p.t861 716.572
R1760 vp_p.n18938 vp_p.t2702 716.572
R1761 vp_p.n17512 vp_p.t1592 716.572
R1762 vp_p.n16085 vp_p.t514 716.572
R1763 vp_p.n14657 vp_p.t2526 716.572
R1764 vp_p.n13403 vp_p.t2389 716.572
R1765 vp_p.n8194 vp_p.t1270 716.572
R1766 vp_p.n8192 vp_p.t1033 716.572
R1767 vp_p.n6770 vp_p.t334 716.572
R1768 vp_p.n5347 vp_p.t84 716.572
R1769 vp_p.n3923 vp_p.t1960 716.572
R1770 vp_p.n2498 vp_p.t1546 716.572
R1771 vp_p.n1072 vp_p.t1297 716.572
R1772 vp_p.n9818 vp_p.t162 716.572
R1773 vp_p.n11255 vp_p.t645 716.572
R1774 vp_p.n12693 vp_p.t2491 716.572
R1775 vp_p.n26896 vp_p.t43 716.572
R1776 vp_p.n25471 vp_p.t2612 716.572
R1777 vp_p.n24049 vp_p.t2377 716.572
R1778 vp_p.n22626 vp_p.t1248 716.572
R1779 vp_p.n21202 vp_p.t1733 716.572
R1780 vp_p.n19777 vp_p.t599 716.572
R1781 vp_p.n18351 vp_p.t2437 716.572
R1782 vp_p.n16924 vp_p.t188 716.572
R1783 vp_p.n15496 vp_p.t268 716.572
R1784 vp_p.n13398 vp_p.t2093 716.572
R1785 vp_p.n7350 vp_p.t2471 716.572
R1786 vp_p.n7348 vp_p.t2216 716.572
R1787 vp_p.n5926 vp_p.t2009 716.572
R1788 vp_p.n4503 vp_p.t1754 716.572
R1789 vp_p.n3079 vp_p.t628 716.572
R1790 vp_p.n1654 vp_p.t205 716.572
R1791 vp_p.n170 vp_p.t2953 716.572
R1792 vp_p.n8909 vp_p.t1829 716.572
R1793 vp_p.n10411 vp_p.t2278 716.572
R1794 vp_p.n11849 vp_p.t1174 716.572
R1795 vp_p.n26053 vp_p.t1252 716.572
R1796 vp_p.n24627 vp_p.t839 716.572
R1797 vp_p.n23205 vp_p.t604 716.572
R1798 vp_p.n21782 vp_p.t2445 716.572
R1799 vp_p.n20358 vp_p.t2924 716.572
R1800 vp_p.n18933 vp_p.t1801 716.572
R1801 vp_p.n17507 vp_p.t674 716.572
R1802 vp_p.n16080 vp_p.t1860 716.572
R1803 vp_p.n14652 vp_p.t1793 716.572
R1804 vp_p.n13393 vp_p.t737 716.572
R1805 vp_p.n8208 vp_p.t78 716.572
R1806 vp_p.n8206 vp_p.t2823 716.572
R1807 vp_p.n6784 vp_p.t1657 716.572
R1808 vp_p.n5361 vp_p.t1410 716.572
R1809 vp_p.n3937 vp_p.t260 716.572
R1810 vp_p.n2512 vp_p.t2835 716.572
R1811 vp_p.n1086 vp_p.t2594 716.572
R1812 vp_p.n9832 vp_p.t1484 716.572
R1813 vp_p.n11269 vp_p.t1955 716.572
R1814 vp_p.n12707 vp_p.t811 716.572
R1815 vp_p.n26910 vp_p.t1867 716.572
R1816 vp_p.n25485 vp_p.t1443 716.572
R1817 vp_p.n24063 vp_p.t1208 716.572
R1818 vp_p.n22640 vp_p.t63 716.572
R1819 vp_p.n21216 vp_p.t545 716.572
R1820 vp_p.n19791 vp_p.t2386 716.572
R1821 vp_p.n18365 vp_p.t1264 716.572
R1822 vp_p.n16938 vp_p.t1507 716.572
R1823 vp_p.n15510 vp_p.t1884 716.572
R1824 vp_p.n13388 vp_p.t391 716.572
R1825 vp_p.n7345 vp_p.t1291 716.572
R1826 vp_p.n7343 vp_p.t1053 716.572
R1827 vp_p.n5921 vp_p.t299 716.572
R1828 vp_p.n4498 vp_p.t69 716.572
R1829 vp_p.n3074 vp_p.t1934 716.572
R1830 vp_p.n1649 vp_p.t1524 716.572
R1831 vp_p.n165 vp_p.t1272 716.572
R1832 vp_p.n8904 vp_p.t130 716.572
R1833 vp_p.n10406 vp_p.t624 716.572
R1834 vp_p.n11844 vp_p.t2470 716.572
R1835 vp_p.n26048 vp_p.t64 716.572
R1836 vp_p.n24622 vp_p.t2636 716.572
R1837 vp_p.n23200 vp_p.t2391 716.572
R1838 vp_p.n21777 vp_p.t1268 716.572
R1839 vp_p.n20353 vp_p.t1749 716.572
R1840 vp_p.n18928 vp_p.t617 716.572
R1841 vp_p.n17502 vp_p.t2465 716.572
R1842 vp_p.n16075 vp_p.t165 716.572
R1843 vp_p.n14647 vp_p.t384 716.572
R1844 vp_p.n13383 vp_p.t2072 716.572
R1845 vp_p.n8222 vp_p.t2896 716.572
R1846 vp_p.n8220 vp_p.t2660 716.572
R1847 vp_p.n6798 vp_p.t2200 716.572
R1848 vp_p.n5375 vp_p.t1980 716.572
R1849 vp_p.n3951 vp_p.t837 716.572
R1850 vp_p.n2526 vp_p.t406 716.572
R1851 vp_p.n1100 vp_p.t178 716.572
R1852 vp_p.n9846 vp_p.t2050 716.572
R1853 vp_p.n11283 vp_p.t2511 716.572
R1854 vp_p.n12721 vp_p.t1387 716.572
R1855 vp_p.n26924 vp_p.t1695 716.572
R1856 vp_p.n25499 vp_p.t1269 716.572
R1857 vp_p.n24077 vp_p.t1037 716.572
R1858 vp_p.n22654 vp_p.t2874 716.572
R1859 vp_p.n21230 vp_p.t366 716.572
R1860 vp_p.n19805 vp_p.t2211 716.572
R1861 vp_p.n18379 vp_p.t1092 716.572
R1862 vp_p.n16952 vp_p.t2073 716.572
R1863 vp_p.n15524 vp_p.t1259 716.572
R1864 vp_p.n13378 vp_p.t954 716.572
R1865 vp_p.n7340 vp_p.t91 716.572
R1866 vp_p.n7338 vp_p.t2839 716.572
R1867 vp_p.n5916 vp_p.t1629 716.572
R1868 vp_p.n4493 vp_p.t1395 716.572
R1869 vp_p.n3069 vp_p.t241 716.572
R1870 vp_p.n1644 vp_p.t2816 716.572
R1871 vp_p.n160 vp_p.t2570 716.572
R1872 vp_p.n8899 vp_p.t1458 716.572
R1873 vp_p.n10401 vp_p.t1927 716.572
R1874 vp_p.n11839 vp_p.t785 716.572
R1875 vp_p.n26043 vp_p.t1882 716.572
R1876 vp_p.n24617 vp_p.t1466 716.572
R1877 vp_p.n23195 vp_p.t1221 716.572
R1878 vp_p.n21772 vp_p.t77 716.572
R1879 vp_p.n20348 vp_p.t570 716.572
R1880 vp_p.n18923 vp_p.t2402 716.572
R1881 vp_p.n17497 vp_p.t1287 716.572
R1882 vp_p.n16070 vp_p.t1488 716.572
R1883 vp_p.n14642 vp_p.t1999 716.572
R1884 vp_p.n13373 vp_p.t376 716.572
R1885 vp_p.n8236 vp_p.t961 716.572
R1886 vp_p.n8234 vp_p.t725 716.572
R1887 vp_p.n6812 vp_p.t1313 716.572
R1888 vp_p.n5389 vp_p.t1069 716.572
R1889 vp_p.n3965 vp_p.t2918 716.572
R1890 vp_p.n2540 vp_p.t2505 716.572
R1891 vp_p.n1114 vp_p.t2247 716.572
R1892 vp_p.n9860 vp_p.t1138 716.572
R1893 vp_p.n11297 vp_p.t1610 716.572
R1894 vp_p.n12735 vp_p.t477 716.572
R1895 vp_p.n26938 vp_p.t2724 716.572
R1896 vp_p.n25513 vp_p.t2317 716.572
R1897 vp_p.n24091 vp_p.t2096 716.572
R1898 vp_p.n22668 vp_p.t937 716.572
R1899 vp_p.n21244 vp_p.t1427 716.572
R1900 vp_p.n19819 vp_p.t275 716.572
R1901 vp_p.n18393 vp_p.t2156 716.572
R1902 vp_p.n16966 vp_p.t1171 716.572
R1903 vp_p.n15538 vp_p.t2720 716.572
R1904 vp_p.n13368 vp_p.t56 716.572
R1905 vp_p.n7335 vp_p.t2573 716.572
R1906 vp_p.n7333 vp_p.t2343 716.572
R1907 vp_p.n5911 vp_p.t213 716.572
R1908 vp_p.n4488 vp_p.t2962 716.572
R1909 vp_p.n3064 vp_p.t1842 716.572
R1910 vp_p.n1639 vp_p.t1413 716.572
R1911 vp_p.n155 vp_p.t1179 716.572
R1912 vp_p.n8894 vp_p.t36 716.572
R1913 vp_p.n10396 vp_p.t521 716.572
R1914 vp_p.n11834 vp_p.t2367 716.572
R1915 vp_p.n26038 vp_p.t1371 716.572
R1916 vp_p.n24612 vp_p.t939 716.572
R1917 vp_p.n23190 vp_p.t712 716.572
R1918 vp_p.n21767 vp_p.t2552 716.572
R1919 vp_p.n20343 vp_p.t46 716.572
R1920 vp_p.n18918 vp_p.t1910 716.572
R1921 vp_p.n17492 vp_p.t765 716.572
R1922 vp_p.n16065 vp_p.t60 716.572
R1923 vp_p.n14637 vp_p.t618 716.572
R1924 vp_p.n13363 vp_p.t1964 716.572
R1925 vp_p.n8250 vp_p.t2762 716.572
R1926 vp_p.n8248 vp_p.t2532 716.572
R1927 vp_p.n6826 vp_p.t2605 716.572
R1928 vp_p.n5403 vp_p.t2373 716.572
R1929 vp_p.n3979 vp_p.t1242 716.572
R1930 vp_p.n2554 vp_p.t826 716.572
R1931 vp_p.n1128 vp_p.t594 716.572
R1932 vp_p.n9874 vp_p.t2428 716.572
R1933 vp_p.n11311 vp_p.t2916 716.572
R1934 vp_p.n12749 vp_p.t1792 716.572
R1935 vp_p.n26952 vp_p.t1566 716.572
R1936 vp_p.n25527 vp_p.t1151 716.572
R1937 vp_p.n24105 vp_p.t897 716.572
R1938 vp_p.n22682 vp_p.t2740 716.572
R1939 vp_p.n21258 vp_p.t231 716.572
R1940 vp_p.n19833 vp_p.t2105 716.572
R1941 vp_p.n18407 vp_p.t958 716.572
R1942 vp_p.n16980 vp_p.t2464 716.572
R1943 vp_p.n15552 vp_p.t1347 716.572
R1944 vp_p.n13358 vp_p.t1377 716.572
R1945 vp_p.n7330 vp_p.t1407 716.572
R1946 vp_p.n7328 vp_p.t1173 716.572
R1947 vp_p.n5906 vp_p.t1536 716.572
R1948 vp_p.n4483 vp_p.t1284 716.572
R1949 vp_p.n3059 vp_p.t145 716.572
R1950 vp_p.n1634 vp_p.t2707 716.572
R1951 vp_p.n150 vp_p.t2475 716.572
R1952 vp_p.n8889 vp_p.t1358 716.572
R1953 vp_p.n10391 vp_p.t1836 716.572
R1954 vp_p.n11829 vp_p.t695 716.572
R1955 vp_p.n26033 vp_p.t184 716.572
R1956 vp_p.n24607 vp_p.t2743 716.572
R1957 vp_p.n23185 vp_p.t2516 716.572
R1958 vp_p.n21762 vp_p.t1392 716.572
R1959 vp_p.n20338 vp_p.t1868 716.572
R1960 vp_p.n18913 vp_p.t723 716.572
R1961 vp_p.n17487 vp_p.t2567 716.572
R1962 vp_p.n16060 vp_p.t1382 716.572
R1963 vp_p.n14632 vp_p.t2197 716.572
R1964 vp_p.n13353 vp_p.t261 716.572
R1965 vp_p.n8264 vp_p.t2593 716.572
R1966 vp_p.n8262 vp_p.t2366 716.572
R1967 vp_p.n6840 vp_p.t194 716.572
R1968 vp_p.n5417 vp_p.t2934 716.572
R1969 vp_p.n3993 vp_p.t1817 716.572
R1970 vp_p.n2568 vp_p.t1401 716.572
R1971 vp_p.n1142 vp_p.t1160 716.572
R1972 vp_p.n9888 vp_p.t13 716.572
R1973 vp_p.n11325 vp_p.t498 716.572
R1974 vp_p.n12763 vp_p.t2346 716.572
R1975 vp_p.n26966 vp_p.t1396 716.572
R1976 vp_p.n25541 vp_p.t963 716.572
R1977 vp_p.n24119 vp_p.t728 716.572
R1978 vp_p.n22696 vp_p.t2572 716.572
R1979 vp_p.n21272 vp_p.t68 716.572
R1980 vp_p.n19847 vp_p.t1929 716.572
R1981 vp_p.n18421 vp_p.t788 716.572
R1982 vp_p.n16994 vp_p.t38 716.572
R1983 vp_p.n15566 vp_p.t716 716.572
R1984 vp_p.n13348 vp_p.t1935 716.572
R1985 vp_p.n7325 vp_p.t2454 716.572
R1986 vp_p.n7323 vp_p.t2204 716.572
R1987 vp_p.n5901 vp_p.t630 716.572
R1988 vp_p.n4478 vp_p.t373 716.572
R1989 vp_p.n3054 vp_p.t2222 716.572
R1990 vp_p.n1629 vp_p.t1830 716.572
R1991 vp_p.n145 vp_p.t1585 716.572
R1992 vp_p.n8884 vp_p.t439 716.572
R1993 vp_p.n10386 vp_p.t912 716.572
R1994 vp_p.n11824 vp_p.t2767 716.572
R1995 vp_p.n26028 vp_p.t1238 716.572
R1996 vp_p.n24602 vp_p.t817 716.572
R1997 vp_p.n23180 vp_p.t591 716.572
R1998 vp_p.n21757 vp_p.t2425 716.572
R1999 vp_p.n20333 vp_p.t2903 716.572
R2000 vp_p.n18908 vp_p.t1786 716.572
R2001 vp_p.n17482 vp_p.t655 716.572
R2002 vp_p.n16055 vp_p.t473 716.572
R2003 vp_p.n14627 vp_p.t696 716.572
R2004 vp_p.n13343 vp_p.t2363 716.572
R2005 vp_p.n8278 vp_p.t1426 716.572
R2006 vp_p.n8276 vp_p.t1192 716.572
R2007 vp_p.n6854 vp_p.t1511 716.572
R2008 vp_p.n5431 vp_p.t1258 716.572
R2009 vp_p.n4007 vp_p.t116 716.572
R2010 vp_p.n2582 vp_p.t2694 716.572
R2011 vp_p.n1156 vp_p.t2453 716.572
R2012 vp_p.n9902 vp_p.t1337 716.572
R2013 vp_p.n11339 vp_p.t1812 716.572
R2014 vp_p.n12777 vp_p.t680 716.572
R2015 vp_p.n26980 vp_p.t204 716.572
R2016 vp_p.n25555 vp_p.t2766 716.572
R2017 vp_p.n24133 vp_p.t2533 716.572
R2018 vp_p.n22710 vp_p.t1406 716.572
R2019 vp_p.n21286 vp_p.t1883 716.572
R2020 vp_p.n19861 vp_p.t735 716.572
R2021 vp_p.n18435 vp_p.t2589 716.572
R2022 vp_p.n17008 vp_p.t1362 716.572
R2023 vp_p.n15580 vp_p.t2298 716.572
R2024 vp_p.n13338 vp_p.t244 716.572
R2025 vp_p.n7320 vp_p.t2274 716.572
R2026 vp_p.n7318 vp_p.t2062 716.572
R2027 vp_p.n5896 vp_p.t1193 716.572
R2028 vp_p.n4473 vp_p.t930 716.572
R2029 vp_p.n3049 vp_p.t2787 716.572
R2030 vp_p.n1624 vp_p.t2378 716.572
R2031 vp_p.n140 vp_p.t2142 716.572
R2032 vp_p.n8879 vp_p.t1007 716.572
R2033 vp_p.n10381 vp_p.t1489 716.572
R2034 vp_p.n11819 vp_p.t344 716.572
R2035 vp_p.n26023 vp_p.t1071 716.572
R2036 vp_p.n24597 vp_p.t663 716.572
R2037 vp_p.n23175 vp_p.t399 716.572
R2038 vp_p.n21752 vp_p.t2251 716.572
R2039 vp_p.n20328 vp_p.t2728 716.572
R2040 vp_p.n18903 vp_p.t1613 716.572
R2041 vp_p.n17477 vp_p.t483 716.572
R2042 vp_p.n16050 vp_p.t1042 716.572
R2043 vp_p.n14622 vp_p.t65 716.572
R2044 vp_p.n13333 vp_p.t2921 716.572
R2045 vp_p.n8292 vp_p.t229 716.572
R2046 vp_p.n8290 vp_p.t2995 716.572
R2047 vp_p.n6868 vp_p.t2803 716.572
R2048 vp_p.n5445 vp_p.t2557 716.572
R2049 vp_p.n4021 vp_p.t1437 716.572
R2050 vp_p.n2596 vp_p.t1029 716.572
R2051 vp_p.n1170 vp_p.t768 716.572
R2052 vp_p.n9916 vp_p.t2627 716.572
R2053 vp_p.n11353 vp_p.t111 716.572
R2054 vp_p.n12791 vp_p.t1995 716.572
R2055 vp_p.n26994 vp_p.t2027 716.572
R2056 vp_p.n25569 vp_p.t1599 716.572
R2057 vp_p.n24147 vp_p.t1361 716.572
R2058 vp_p.n22724 vp_p.t217 716.572
R2059 vp_p.n21300 vp_p.t697 716.572
R2060 vp_p.n19875 vp_p.t2541 716.572
R2061 vp_p.n18449 vp_p.t1423 716.572
R2062 vp_p.n17022 vp_p.t2659 716.572
R2063 vp_p.n15594 vp_p.t908 716.572
R2064 vp_p.n13328 vp_p.t1576 716.572
R2065 vp_p.n7315 vp_p.t1105 716.572
R2066 vp_p.n7313 vp_p.t867 716.572
R2067 vp_p.n5891 vp_p.t2488 716.572
R2068 vp_p.n4468 vp_p.t2234 716.572
R2069 vp_p.n3044 vp_p.t1124 716.572
R2070 vp_p.n1619 vp_p.t705 716.572
R2071 vp_p.n135 vp_p.t461 716.572
R2072 vp_p.n8874 vp_p.t2308 716.572
R2073 vp_p.n10376 vp_p.t2784 716.572
R2074 vp_p.n11814 vp_p.t1671 716.572
R2075 vp_p.n26018 vp_p.t2864 716.572
R2076 vp_p.n24592 vp_p.t2452 716.572
R2077 vp_p.n23170 vp_p.t2205 716.572
R2078 vp_p.n21747 vp_p.t1084 716.572
R2079 vp_p.n20323 vp_p.t1570 716.572
R2080 vp_p.n18898 vp_p.t414 716.572
R2081 vp_p.n17472 vp_p.t2270 716.572
R2082 vp_p.n16045 vp_p.t2341 716.572
R2083 vp_p.n14617 vp_p.t1674 716.572
R2084 vp_p.n13323 vp_p.t1246 716.572
R2085 vp_p.n8306 vp_p.t1985 716.572
R2086 vp_p.n8304 vp_p.t1735 716.572
R2087 vp_p.n6882 vp_p.t2171 716.572
R2088 vp_p.n5459 vp_p.t1933 716.572
R2089 vp_p.n4035 vp_p.t790 716.572
R2090 vp_p.n2610 vp_p.t383 716.572
R2091 vp_p.n1184 vp_p.t134 716.572
R2092 vp_p.n9930 vp_p.t2015 716.572
R2093 vp_p.n11367 vp_p.t2469 716.572
R2094 vp_p.n12805 vp_p.t1351 716.572
R2095 vp_p.n27008 vp_p.t740 716.572
R2096 vp_p.n25583 vp_p.t327 716.572
R2097 vp_p.n24161 vp_p.t83 716.572
R2098 vp_p.n22738 vp_p.t1959 716.572
R2099 vp_p.n21314 vp_p.t2412 716.572
R2100 vp_p.n19889 vp_p.t1296 716.572
R2101 vp_p.n18463 vp_p.t160 716.572
R2102 vp_p.n17036 vp_p.t2041 716.572
R2103 vp_p.n15608 vp_p.t2400 716.572
R2104 vp_p.n13318 vp_p.t916 716.572
R2105 vp_p.n7310 vp_p.t2899 716.572
R2106 vp_p.n7308 vp_p.t2664 716.572
R2107 vp_p.n5886 vp_p.t810 716.572
R2108 vp_p.n4463 vp_p.t581 716.572
R2109 vp_p.n3039 vp_p.t2419 716.572
R2110 vp_p.n1614 vp_p.t2034 716.572
R2111 vp_p.n130 vp_p.t1780 716.572
R2112 vp_p.n8869 vp_p.t648 716.572
R2113 vp_p.n10371 vp_p.t1118 716.572
R2114 vp_p.n11809 vp_p.t2977 716.572
R2115 vp_p.n26013 vp_p.t1706 716.572
R2116 vp_p.n24587 vp_p.t1277 716.572
R2117 vp_p.n23165 vp_p.t1044 716.572
R2118 vp_p.n21742 vp_p.t2881 716.572
R2119 vp_p.n20318 vp_p.t371 716.572
R2120 vp_p.n18893 vp_p.t2220 716.572
R2121 vp_p.n17467 vp_p.t1100 716.572
R2122 vp_p.n16040 vp_p.t677 716.572
R2123 vp_p.n14612 vp_p.t254 716.572
R2124 vp_p.n13313 vp_p.t2549 716.572
R2125 vp_p.n8320 vp_p.t776 716.572
R2126 vp_p.n8318 vp_p.t549 716.572
R2127 vp_p.n6896 vp_p.t503 716.572
R2128 vp_p.n5473 vp_p.t240 716.572
R2129 vp_p.n4049 vp_p.t2117 716.572
R2130 vp_p.n2624 vp_p.t1713 716.572
R2131 vp_p.n1198 vp_p.t1457 716.572
R2132 vp_p.n9944 vp_p.t307 716.572
R2133 vp_p.n11381 vp_p.t787 716.572
R2134 vp_p.n12819 vp_p.t2647 716.572
R2135 vp_p.n27022 vp_p.t2548 716.572
R2136 vp_p.n25597 vp_p.t2150 716.572
R2137 vp_p.n24175 vp_p.t1899 716.572
R2138 vp_p.n22752 vp_p.t758 716.572
R2139 vp_p.n21328 vp_p.t1241 716.572
R2140 vp_p.n19903 vp_p.t97 716.572
R2141 vp_p.n18477 vp_p.t1979 716.572
R2142 vp_p.n17050 vp_p.t342 716.572
R2143 vp_p.n15622 vp_p.t1021 716.572
R2144 vp_p.n13308 vp_p.t2224 716.572
R2145 vp_p.n7305 vp_p.t2726 716.572
R2146 vp_p.n7303 vp_p.t2497 716.572
R2147 vp_p.n5881 vp_p.t1385 716.572
R2148 vp_p.n4458 vp_p.t1142 716.572
R2149 vp_p.n3034 vp_p.t2999 716.572
R2150 vp_p.n1609 vp_p.t2566 716.572
R2151 vp_p.n125 vp_p.t2332 716.572
R2152 vp_p.n8864 vp_p.t1210 716.572
R2153 vp_p.n10366 vp_p.t1688 716.572
R2154 vp_p.n11804 vp_p.t548 716.572
R2155 vp_p.n26008 vp_p.t1533 716.572
R2156 vp_p.n24582 vp_p.t1108 716.572
R2157 vp_p.n23160 vp_p.t868 716.572
R2158 vp_p.n21737 vp_p.t2705 716.572
R2159 vp_p.n20313 vp_p.t207 716.572
R2160 vp_p.n18888 vp_p.t2076 716.572
R2161 vp_p.n17462 vp_p.t919 716.572
R2162 vp_p.n16035 vp_p.t1228 716.572
R2163 vp_p.n14607 vp_p.t2625 716.572
R2164 vp_p.n13303 vp_p.t121 716.572
R2165 vp_p.n8334 vp_p.t2580 716.572
R2166 vp_p.n8332 vp_p.t2349 716.572
R2167 vp_p.n6910 vp_p.t1818 716.572
R2168 vp_p.n5487 vp_p.t1575 716.572
R2169 vp_p.n4063 vp_p.t419 716.572
R2170 vp_p.n2638 vp_p.t19 716.572
R2171 vp_p.n1212 vp_p.t2748 716.572
R2172 vp_p.n9958 vp_p.t1632 716.572
R2173 vp_p.n11395 vp_p.t2113 716.572
R2174 vp_p.n12833 vp_p.t965 716.572
R2175 vp_p.n27036 vp_p.t1381 716.572
R2176 vp_p.n25611 vp_p.t950 716.572
R2177 vp_p.n24189 vp_p.t714 716.572
R2178 vp_p.n22766 vp_p.t2562 716.572
R2179 vp_p.n21342 vp_p.t54 716.572
R2180 vp_p.n19917 vp_p.t1917 716.572
R2181 vp_p.n18491 vp_p.t770 716.572
R2182 vp_p.n17064 vp_p.t1666 716.572
R2183 vp_p.n15636 vp_p.t2596 716.572
R2184 vp_p.n13298 vp_p.t567 716.572
R2185 vp_p.n7300 vp_p.t2520 716.572
R2186 vp_p.n7298 vp_p.t2261 716.572
R2187 vp_p.n5876 vp_p.t799 716.572
R2188 vp_p.n4453 vp_p.t573 716.572
R2189 vp_p.n3029 vp_p.t2409 716.572
R2190 vp_p.n1604 vp_p.t2028 716.572
R2191 vp_p.n120 vp_p.t1773 716.572
R2192 vp_p.n8859 vp_p.t639 716.572
R2193 vp_p.n10361 vp_p.t1114 716.572
R2194 vp_p.n11799 vp_p.t2971 716.572
R2195 vp_p.n26003 vp_p.t1299 716.572
R2196 vp_p.n24577 vp_p.t884 716.572
R2197 vp_p.n23155 vp_p.t650 716.572
R2198 vp_p.n21732 vp_p.t2496 716.572
R2199 vp_p.n20308 vp_p.t2976 716.572
R2200 vp_p.n18883 vp_p.t1855 716.572
R2201 vp_p.n17457 vp_p.t709 716.572
R2202 vp_p.n16030 vp_p.t672 716.572
R2203 vp_p.n14602 vp_p.t96 716.572
R2204 vp_p.n13293 vp_p.t2543 716.572
R2205 vp_p.n8348 vp_p.t1156 716.572
R2206 vp_p.n8346 vp_p.t900 716.572
R2207 vp_p.n6924 vp_p.t2696 716.572
R2208 vp_p.n5501 vp_p.t2457 716.572
R2209 vp_p.n4077 vp_p.t1340 716.572
R2210 vp_p.n2652 vp_p.t907 716.572
R2211 vp_p.n1226 vp_p.t681 716.572
R2212 vp_p.n9972 vp_p.t2527 716.572
R2213 vp_p.n11409 vp_p.t18 716.572
R2214 vp_p.n12847 vp_p.t1881 716.572
R2215 vp_p.n27050 vp_p.t2902 716.572
R2216 vp_p.n25625 vp_p.t2498 716.572
R2217 vp_p.n24203 vp_p.t2242 716.572
R2218 vp_p.n22780 vp_p.t1127 716.572
R2219 vp_p.n21356 vp_p.t1603 716.572
R2220 vp_p.n19931 vp_p.t468 716.572
R2221 vp_p.n18505 vp_p.t2316 716.572
R2222 vp_p.n17078 vp_p.t2545 716.572
R2223 vp_p.n15650 vp_p.t969 716.572
R2224 vp_p.n13288 vp_p.t1465 716.572
R2225 vp_p.n7295 vp_p.t994 716.572
R2226 vp_p.n7293 vp_p.t743 716.572
R2227 vp_p.n5871 vp_p.t140 716.572
R2228 vp_p.n4448 vp_p.t2884 716.572
R2229 vp_p.n3024 vp_p.t1765 716.572
R2230 vp_p.n1599 vp_p.t1356 716.572
R2231 vp_p.n115 vp_p.t1103 716.572
R2232 vp_p.n8854 vp_p.t2963 716.572
R2233 vp_p.n10356 vp_p.t438 716.572
R2234 vp_p.n11794 vp_p.t2289 716.572
R2235 vp_p.n25998 vp_p.t2749 716.572
R2236 vp_p.n24572 vp_p.t2351 716.572
R2237 vp_p.n23150 vp_p.t2116 716.572
R2238 vp_p.n21727 vp_p.t968 716.572
R2239 vp_p.n20303 vp_p.t1456 716.572
R2240 vp_p.n18878 vp_p.t306 716.572
R2241 vp_p.n17452 vp_p.t2174 716.572
R2242 vp_p.n16025 vp_p.t2991 716.572
R2243 vp_p.n14597 vp_p.t938 716.572
R2244 vp_p.n13283 vp_p.t1893 716.572
R2245 vp_p.n8362 vp_p.t2952 716.572
R2246 vp_p.n8360 vp_p.t2699 716.572
R2247 vp_p.n6938 vp_p.t1036 716.572
R2248 vp_p.n5515 vp_p.t772 716.572
R2249 vp_p.n4091 vp_p.t2634 716.572
R2250 vp_p.n2666 vp_p.t2207 716.572
R2251 vp_p.n1240 vp_p.t1998 716.572
R2252 vp_p.n9986 vp_p.t852 716.572
R2253 vp_p.n11423 vp_p.t1336 716.572
R2254 vp_p.n12861 vp_p.t197 716.572
R2255 vp_p.n27064 vp_p.t1736 716.572
R2256 vp_p.n25639 vp_p.t1322 716.572
R2257 vp_p.n24217 vp_p.t1075 716.572
R2258 vp_p.n22794 vp_p.t2925 716.572
R2259 vp_p.n21370 vp_p.t404 716.572
R2260 vp_p.n19945 vp_p.t2256 716.572
R2261 vp_p.n18519 vp_p.t1150 716.572
R2262 vp_p.n17092 vp_p.t880 716.572
R2263 vp_p.n15664 vp_p.t2556 716.572
R2264 vp_p.n13278 vp_p.t2754 716.572
R2265 vp_p.n7290 vp_p.t821 716.572
R2266 vp_p.n7288 vp_p.t592 716.572
R2267 vp_p.n5866 vp_p.t708 716.572
R2268 vp_p.n4443 vp_p.t463 716.572
R2269 vp_p.n3019 vp_p.t2311 716.572
R2270 vp_p.n1594 vp_p.t1905 716.572
R2271 vp_p.n110 vp_p.t1673 716.572
R2272 vp_p.n8849 vp_p.t536 716.572
R2273 vp_p.n10351 vp_p.t1009 716.572
R2274 vp_p.n11789 vp_p.t2851 716.572
R2275 vp_p.n25993 vp_p.t2582 716.572
R2276 vp_p.n24567 vp_p.t2177 716.572
R2277 vp_p.n23145 vp_p.t1941 716.572
R2278 vp_p.n21722 vp_p.t795 716.572
R2279 vp_p.n20298 vp_p.t1283 716.572
R2280 vp_p.n18873 vp_p.t144 716.572
R2281 vp_p.n17447 vp_p.t2023 716.572
R2282 vp_p.n16020 vp_p.t563 716.572
R2283 vp_p.n14592 vp_p.t319 716.572
R2284 vp_p.n13273 vp_p.t2442 716.572
R2285 vp_p.n8376 vp_p.t1020 716.572
R2286 vp_p.n8374 vp_p.t762 716.572
R2287 vp_p.n6952 vp_p.t110 716.572
R2288 vp_p.n5529 vp_p.t2860 716.572
R2289 vp_p.n4105 vp_p.t1744 716.572
R2290 vp_p.n2680 vp_p.t1331 716.572
R2291 vp_p.n1254 vp_p.t1080 716.572
R2292 vp_p.n10000 vp_p.t2937 716.572
R2293 vp_p.n11437 vp_p.t409 716.572
R2294 vp_p.n12875 vp_p.t2264 716.572
R2295 vp_p.n27078 vp_p.t2773 716.572
R2296 vp_p.n25653 vp_p.t2368 716.572
R2297 vp_p.n24231 vp_p.t2135 716.572
R2298 vp_p.n22808 vp_p.t993 716.572
R2299 vp_p.n21384 vp_p.t1481 716.572
R2300 vp_p.n19959 vp_p.t333 716.572
R2301 vp_p.n18533 vp_p.t2190 716.572
R2302 vp_p.n17106 vp_p.t2967 716.572
R2303 vp_p.n15678 vp_p.t1059 716.572
R2304 vp_p.n13268 vp_p.t1874 716.572
R2305 vp_p.n7285 vp_p.t2619 716.572
R2306 vp_p.n7283 vp_p.t2382 716.572
R2307 vp_p.n5861 vp_p.t2039 716.572
R2308 vp_p.n4438 vp_p.t1785 716.572
R2309 vp_p.n3014 vp_p.t653 716.572
R2310 vp_p.n1589 vp_p.t222 716.572
R2311 vp_p.n105 vp_p.t2981 716.572
R2312 vp_p.n8844 vp_p.t1857 716.572
R2313 vp_p.n10346 vp_p.t2307 716.572
R2314 vp_p.n11784 vp_p.t1197 716.572
R2315 vp_p.n25988 vp_p.t1414 716.572
R2316 vp_p.n24562 vp_p.t995 716.572
R2317 vp_p.n23140 vp_p.t742 716.572
R2318 vp_p.n21717 vp_p.t2595 716.572
R2319 vp_p.n20293 vp_p.t87 716.572
R2320 vp_p.n18868 vp_p.t1963 716.572
R2321 vp_p.n17442 vp_p.t816 716.572
R2322 vp_p.n16015 vp_p.t1878 716.572
R2323 vp_p.n14587 vp_p.t1923 716.572
R2324 vp_p.n13263 vp_p.t761 716.572
R2325 vp_p.n8390 vp_p.t847 716.572
R2326 vp_p.n8388 vp_p.t611 716.572
R2327 vp_p.n6966 vp_p.t690 716.572
R2328 vp_p.n5543 vp_p.t430 716.572
R2329 vp_p.n4119 vp_p.t2282 716.572
R2330 vp_p.n2694 vp_p.t1891 716.572
R2331 vp_p.n1268 vp_p.t1645 716.572
R2332 vp_p.n10014 vp_p.t516 716.572
R2333 vp_p.n11451 vp_p.t981 716.572
R2334 vp_p.n12889 vp_p.t2830 716.572
R2335 vp_p.n27092 vp_p.t2600 716.572
R2336 vp_p.n25667 vp_p.t2192 716.572
R2337 vp_p.n24245 vp_p.t1970 716.572
R2338 vp_p.n22822 vp_p.t820 716.572
R2339 vp_p.n21398 vp_p.t1303 716.572
R2340 vp_p.n19973 vp_p.t167 716.572
R2341 vp_p.n18547 vp_p.t2042 716.572
R2342 vp_p.n17120 vp_p.t540 716.572
R2343 vp_p.n15692 vp_p.t421 716.572
R2344 vp_p.n13258 vp_p.t2413 716.572
R2345 vp_p.n7280 vp_p.t1452 716.572
R2346 vp_p.n7278 vp_p.t1213 716.572
R2347 vp_p.n5856 vp_p.t336 716.572
R2348 vp_p.n4433 vp_p.t86 716.572
R2349 vp_p.n3009 vp_p.t1962 716.572
R2350 vp_p.n1584 vp_p.t1549 716.572
R2351 vp_p.n100 vp_p.t1298 716.572
R2352 vp_p.n8839 vp_p.t164 716.572
R2353 vp_p.n10341 vp_p.t649 716.572
R2354 vp_p.n11779 vp_p.t2495 716.572
R2355 vp_p.n25983 vp_p.t221 716.572
R2356 vp_p.n24557 vp_p.t2791 716.572
R2357 vp_p.n23135 vp_p.t2550 716.572
R2358 vp_p.n21712 vp_p.t1429 716.572
R2359 vp_p.n20288 vp_p.t1904 716.572
R2360 vp_p.n18863 vp_p.t760 716.572
R2361 vp_p.n17437 vp_p.t2613 716.572
R2362 vp_p.n16010 vp_p.t192 716.572
R2363 vp_p.n14582 vp_p.t532 716.572
R2364 vp_p.n13253 vp_p.t2095 716.572
R2365 vp_p.n8404 vp_p.t2301 716.572
R2366 vp_p.n8402 vp_p.t2084 716.572
R2367 vp_p.n6980 vp_p.t22 716.572
R2368 vp_p.n5557 vp_p.t2751 716.572
R2369 vp_p.n4133 vp_p.t1636 716.572
R2370 vp_p.n2708 vp_p.t1224 716.572
R2371 vp_p.n1282 vp_p.t970 716.572
R2372 vp_p.n10028 vp_p.t2824 716.572
R2373 vp_p.n11465 vp_p.t305 716.572
R2374 vp_p.n12903 vp_p.t2173 716.572
R2375 vp_p.n27106 vp_p.t1091 716.572
R2376 vp_p.n25681 vp_p.t684 716.572
R2377 vp_p.n24259 vp_p.t423 716.572
R2378 vp_p.n22836 vp_p.t2277 716.572
R2379 vp_p.n21412 vp_p.t2753 716.572
R2380 vp_p.n19987 vp_p.t1638 716.572
R2381 vp_p.n18561 vp_p.t509 716.572
R2382 vp_p.n17134 vp_p.t2845 716.572
R2383 vp_p.n15706 vp_p.t1279 716.572
R2384 vp_p.n13248 vp_p.t1768 716.572
R2385 vp_p.n7275 vp_p.t531 716.572
R2386 vp_p.n7273 vp_p.t267 716.572
R2387 vp_p.n5851 vp_p.t1690 716.572
R2388 vp_p.n4428 vp_p.t1432 716.572
R2389 vp_p.n3004 vp_p.t282 716.572
R2390 vp_p.n1579 vp_p.t2867 716.572
R2391 vp_p.n95 vp_p.t2618 716.572
R2392 vp_p.n8834 vp_p.t1508 716.572
R2393 vp_p.n10336 vp_p.t1990 716.572
R2394 vp_p.n11774 vp_p.t843 716.572
R2395 vp_p.n25978 vp_p.t2281 716.572
R2396 vp_p.n24552 vp_p.t1888 716.572
R2397 vp_p.n23130 vp_p.t1642 716.572
R2398 vp_p.n21707 vp_p.t513 716.572
R2399 vp_p.n20283 vp_p.t977 716.572
R2400 vp_p.n18858 vp_p.t2829 716.572
R2401 vp_p.n17432 vp_p.t1723 716.572
R2402 vp_p.n16005 vp_p.t1539 716.572
R2403 vp_p.n14577 vp_p.t2765 716.572
R2404 vp_p.n13243 vp_p.t415 716.572
R2405 vp_p.n8418 vp_p.t1136 716.572
R2406 vp_p.n8416 vp_p.t887 716.572
R2407 vp_p.n6994 vp_p.t1341 716.572
R2408 vp_p.n5571 vp_p.t1086 716.572
R2409 vp_p.n4147 vp_p.t2947 716.572
R2410 vp_p.n2722 vp_p.t2529 716.572
R2411 vp_p.n1296 vp_p.t2273 716.572
R2412 vp_p.n10042 vp_p.t1169 716.572
R2413 vp_p.n11479 vp_p.t1635 716.572
R2414 vp_p.n12917 vp_p.t506 716.572
R2415 vp_p.n27120 vp_p.t2892 716.572
R2416 vp_p.n25695 vp_p.t2479 716.572
R2417 vp_p.n24273 vp_p.t2229 716.572
R2418 vp_p.n22850 vp_p.t1113 716.572
R2419 vp_p.n21426 vp_p.t1596 716.572
R2420 vp_p.n20001 vp_p.t452 716.572
R2421 vp_p.n18575 vp_p.t2297 716.572
R2422 vp_p.n17148 vp_p.t1191 716.572
R2423 vp_p.n15720 vp_p.t2859 716.572
R2424 vp_p.n13238 vp_p.t76 716.572
R2425 vp_p.n7270 vp_p.t2331 716.572
R2426 vp_p.n7268 vp_p.t2101 716.572
R2427 vp_p.n5846 vp_p.t2997 716.572
R2428 vp_p.n4423 vp_p.t2731 716.572
R2429 vp_p.n2999 vp_p.t1614 716.572
R2430 vp_p.n1574 vp_p.t1207 716.572
R2431 vp_p.n90 vp_p.t946 716.572
R2432 vp_p.n8829 vp_p.t2802 716.572
R2433 vp_p.n10331 vp_p.t278 716.572
R2434 vp_p.n11769 vp_p.t2159 716.572
R2435 vp_p.n25973 vp_p.t1117 716.572
R2436 vp_p.n24547 vp_p.t700 716.572
R2437 vp_p.n23125 vp_p.t454 716.572
R2438 vp_p.n21702 vp_p.t2300 716.572
R2439 vp_p.n20278 vp_p.t2777 716.572
R2440 vp_p.n18853 vp_p.t1665 716.572
R2441 vp_p.n17427 vp_p.t527 716.572
R2442 vp_p.n16000 vp_p.t2826 716.572
R2443 vp_p.n14572 vp_p.t1391 716.572
R2444 vp_p.n13233 vp_p.t1747 716.572
R2445 vp_p.n8432 vp_p.t2933 716.572
R2446 vp_p.n8430 vp_p.t2688 716.572
R2447 vp_p.n7008 vp_p.t2635 716.572
R2448 vp_p.n5585 vp_p.t2390 716.572
R2449 vp_p.n4161 vp_p.t1267 716.572
R2450 vp_p.n2736 vp_p.t854 716.572
R2451 vp_p.n1310 vp_p.t615 716.572
R2452 vp_p.n10056 vp_p.t2461 716.572
R2453 vp_p.n11493 vp_p.t2943 716.572
R2454 vp_p.n12931 vp_p.t1820 716.572
R2455 vp_p.n27134 vp_p.t1730 716.572
R2456 vp_p.n25709 vp_p.t1305 716.572
R2457 vp_p.n24287 vp_p.t1065 716.572
R2458 vp_p.n22864 vp_p.t2909 716.572
R2459 vp_p.n21440 vp_p.t393 716.572
R2460 vp_p.n20015 vp_p.t2244 716.572
R2461 vp_p.n18589 vp_p.t1132 716.572
R2462 vp_p.n17162 vp_p.t2487 716.572
R2463 vp_p.n15734 vp_p.t1486 716.572
R2464 vp_p.n13228 vp_p.t1403 716.572
R2465 vp_p.n7265 vp_p.t1163 716.572
R2466 vp_p.n7263 vp_p.t902 716.572
R2467 vp_p.n5841 vp_p.t1316 716.572
R2468 vp_p.n4418 vp_p.t1070 716.572
R2469 vp_p.n2994 vp_p.t2920 716.572
R2470 vp_p.n1569 vp_p.t2508 716.572
R2471 vp_p.n85 vp_p.t2248 716.572
R2472 vp_p.n8824 vp_p.t1141 716.572
R2473 vp_p.n10326 vp_p.t1611 716.572
R2474 vp_p.n11764 vp_p.t482 716.572
R2475 vp_p.n25968 vp_p.t2915 716.572
R2476 vp_p.n24542 vp_p.t2503 716.572
R2477 vp_p.n23120 vp_p.t2246 716.572
R2478 vp_p.n21697 vp_p.t1135 716.572
R2479 vp_p.n20273 vp_p.t1608 716.572
R2480 vp_p.n18848 vp_p.t476 716.572
R2481 vp_p.n17422 vp_p.t2324 716.572
R2482 vp_p.n15995 vp_p.t1172 716.572
R2483 vp_p.n14567 vp_p.t2980 716.572
R2484 vp_p.n13223 vp_p.t61 716.572
R2485 vp_p.n8446 vp_p.t2035 716.572
R2486 vp_p.n8444 vp_p.t1781 716.572
R2487 vp_p.n7022 vp_p.t988 716.572
R2488 vp_p.n5599 vp_p.t736 716.572
R2489 vp_p.n4175 vp_p.t2590 716.572
R2490 vp_p.n2750 vp_p.t2186 716.572
R2491 vp_p.n1324 vp_p.t1953 716.572
R2492 vp_p.n10070 vp_p.t808 716.572
R2493 vp_p.n11507 vp_p.t1293 716.572
R2494 vp_p.n12945 vp_p.t155 716.572
R2495 vp_p.n27148 vp_p.t789 716.572
R2496 vp_p.n25723 vp_p.t380 716.572
R2497 vp_p.n24301 vp_p.t129 716.572
R2498 vp_p.n22878 vp_p.t2013 716.572
R2499 vp_p.n21454 vp_p.t2468 716.572
R2500 vp_p.n20029 vp_p.t1349 716.572
R2501 vp_p.n18603 vp_p.t206 716.572
R2502 vp_p.n17176 vp_p.t841 716.572
R2503 vp_p.n15748 vp_p.t731 716.572
R2504 vp_p.n13218 vp_p.t2715 716.572
R2505 vp_p.n7260 vp_p.t2958 716.572
R2506 vp_p.n7258 vp_p.t2701 716.572
R2507 vp_p.n5836 vp_p.t2608 716.572
R2508 vp_p.n4413 vp_p.t2376 716.572
R2509 vp_p.n2989 vp_p.t1245 716.572
R2510 vp_p.n1564 vp_p.t830 716.572
R2511 vp_p.n80 vp_p.t596 716.572
R2512 vp_p.n8819 vp_p.t2432 716.572
R2513 vp_p.n10321 vp_p.t2917 716.572
R2514 vp_p.n11759 vp_p.t1795 716.572
R2515 vp_p.n25963 vp_p.t1743 716.572
R2516 vp_p.n24537 vp_p.t1329 716.572
R2517 vp_p.n23115 vp_p.t1078 716.572
R2518 vp_p.n21692 vp_p.t2931 716.572
R2519 vp_p.n20268 vp_p.t408 716.572
R2520 vp_p.n18843 vp_p.t2263 716.572
R2521 vp_p.n17417 vp_p.t1157 716.572
R2522 vp_p.n15990 vp_p.t2466 716.572
R2523 vp_p.n14562 vp_p.t1588 716.572
R2524 vp_p.n13213 vp_p.t1380 716.572
R2525 vp_p.n8460 vp_p.t835 716.572
R2526 vp_p.n8458 vp_p.t597 716.572
R2527 vp_p.n7036 vp_p.t2288 716.572
R2528 vp_p.n5613 vp_p.t2071 716.572
R2529 vp_p.n4189 vp_p.t915 716.572
R2530 vp_p.n2764 vp_p.t518 716.572
R2531 vp_p.n1338 vp_p.t253 716.572
R2532 vp_p.n10084 vp_p.t2131 716.572
R2533 vp_p.n11521 vp_p.t2587 716.572
R2534 vp_p.n12959 vp_p.t1476 716.572
R2535 vp_p.n27162 vp_p.t2588 716.572
R2536 vp_p.n25737 vp_p.t2184 716.572
R2537 vp_p.n24315 vp_p.t1947 716.572
R2538 vp_p.n22892 vp_p.t803 716.572
R2539 vp_p.n21468 vp_p.t1290 716.572
R2540 vp_p.n20043 vp_p.t152 716.572
R2541 vp_p.n18617 vp_p.t2030 716.572
R2542 vp_p.n17190 vp_p.t2155 716.572
R2543 vp_p.n15762 vp_p.t2323 716.572
R2544 vp_p.n13208 vp_p.t1057 716.572
R2545 vp_p.n7255 vp_p.t2441 716.572
R2546 vp_p.n7253 vp_p.t2196 716.572
R2547 vp_p.n5831 vp_p.t1212 716.572
R2548 vp_p.n4408 vp_p.t953 716.572
R2549 vp_p.n2984 vp_p.t2810 716.572
R2550 vp_p.n1559 vp_p.t2393 716.572
R2551 vp_p.n75 vp_p.t2164 716.572
R2552 vp_p.n8814 vp_p.t1041 716.572
R2553 vp_p.n10316 vp_p.t1518 716.572
R2554 vp_p.n11754 vp_p.t370 716.572
R2555 vp_p.n25958 vp_p.t1229 716.572
R2556 vp_p.n24532 vp_p.t807 716.572
R2557 vp_p.n23110 vp_p.t580 716.572
R2558 vp_p.n21687 vp_p.t2416 716.572
R2559 vp_p.n20263 vp_p.t2894 716.572
R2560 vp_p.n18838 vp_p.t1777 716.572
R2561 vp_p.n17412 vp_p.t644 716.572
R2562 vp_p.n15985 vp_p.t1058 716.572
R2563 vp_p.n14557 vp_p.t209 716.572
R2564 vp_p.n13203 vp_p.t2950 716.572
R2565 vp_p.n8474 vp_p.t2629 716.572
R2566 vp_p.n8472 vp_p.t2385 716.572
R2567 vp_p.n7050 vp_p.t631 716.572
R2568 vp_p.n5627 vp_p.t379 716.572
R2569 vp_p.n4203 vp_p.t2223 716.572
R2570 vp_p.n2778 vp_p.t1835 716.572
R2571 vp_p.n1352 vp_p.t1591 716.572
R2572 vp_p.n10098 vp_p.t446 716.572
R2573 vp_p.n11535 vp_p.t914 716.572
R2574 vp_p.n12973 vp_p.t2768 716.572
R2575 vp_p.n27176 vp_p.t1422 716.572
R2576 vp_p.n25751 vp_p.t1004 716.572
R2577 vp_p.n24329 vp_p.t750 716.572
R2578 vp_p.n22906 vp_p.t2604 716.572
R2579 vp_p.n21482 vp_p.t90 716.572
R2580 vp_p.n20057 vp_p.t1972 716.572
R2581 vp_p.n18631 vp_p.t823 716.572
R2582 vp_p.n17204 vp_p.t475 716.572
R2583 vp_p.n15776 vp_p.t922 716.572
R2584 vp_p.n13198 vp_p.t2365 716.572
R2585 vp_p.n7250 vp_p.t525 716.572
R2586 vp_p.n7248 vp_p.t258 716.572
R2587 vp_p.n5826 vp_p.t285 716.572
R2588 vp_p.n4403 vp_p.t59 716.572
R2589 vp_p.n2979 vp_p.t1919 716.572
R2590 vp_p.n1554 vp_p.t1515 716.572
R2591 vp_p.n70 vp_p.t1257 716.572
R2592 vp_p.n8809 vp_p.t115 716.572
R2593 vp_p.n10311 vp_p.t610 716.572
R2594 vp_p.n11749 vp_p.t2451 716.572
R2595 vp_p.n25953 vp_p.t2269 716.572
R2596 vp_p.n24527 vp_p.t1880 716.572
R2597 vp_p.n23105 vp_p.t1628 716.572
R2598 vp_p.n21682 vp_p.t502 716.572
R2599 vp_p.n20258 vp_p.t960 716.572
R2600 vp_p.n18833 vp_p.t2815 716.572
R2601 vp_p.n17407 vp_p.t1712 716.572
R2602 vp_p.n15980 vp_p.t148 716.572
R2603 vp_p.n14552 vp_p.t1694 716.572
R2604 vp_p.n13193 vp_p.t2059 716.572
R2605 vp_p.n8488 vp_p.t2463 716.572
R2606 vp_p.n8486 vp_p.t2206 716.572
R2607 vp_p.n7064 vp_p.t1194 716.572
R2608 vp_p.n5641 vp_p.t933 716.572
R2609 vp_p.n4217 vp_p.t2788 716.572
R2610 vp_p.n2792 vp_p.t2379 716.572
R2611 vp_p.n1366 vp_p.t2145 716.572
R2612 vp_p.n10112 vp_p.t1014 716.572
R2613 vp_p.n11549 vp_p.t1493 716.572
R2614 vp_p.n12987 vp_p.t347 716.572
R2615 vp_p.n27190 vp_p.t1247 716.572
R2616 vp_p.n25765 vp_p.t834 716.572
R2617 vp_p.n24343 vp_p.t598 716.572
R2618 vp_p.n22920 vp_p.t2436 716.572
R2619 vp_p.n21496 vp_p.t2919 716.572
R2620 vp_p.n20071 vp_p.t1797 716.572
R2621 vp_p.n18645 vp_p.t667 716.572
R2622 vp_p.n17218 vp_p.t1043 716.572
R2623 vp_p.n15790 vp_p.t294 716.572
R2624 vp_p.n13188 vp_p.t2923 716.572
R2625 vp_p.n7245 vp_p.t2310 716.572
R2626 vp_p.n7243 vp_p.t2091 716.572
R2627 vp_p.n5821 vp_p.t1615 716.572
R2628 vp_p.n4398 vp_p.t1376 716.572
R2629 vp_p.n2974 vp_p.t228 716.572
R2630 vp_p.n1549 vp_p.t2804 716.572
R2631 vp_p.n65 vp_p.t2559 716.572
R2632 vp_p.n8804 vp_p.t1440 716.572
R2633 vp_p.n10306 vp_p.t1914 716.572
R2634 vp_p.n11744 vp_p.t769 716.572
R2635 vp_p.n25948 vp_p.t1099 716.572
R2636 vp_p.n24522 vp_p.t691 716.572
R2637 vp_p.n23100 vp_p.t433 716.572
R2638 vp_p.n21677 vp_p.t2285 716.572
R2639 vp_p.n20253 vp_p.t2761 716.572
R2640 vp_p.n18828 vp_p.t1648 716.572
R2641 vp_p.n17402 vp_p.t517 716.572
R2642 vp_p.n15975 vp_p.t1471 716.572
R2643 vp_p.n14547 vp_p.t271 716.572
R2644 vp_p.n13183 vp_p.t362 716.572
R2645 vp_p.n8502 vp_p.t3 716.572
R2646 vp_p.n8500 vp_p.t2737 716.572
R2647 vp_p.n7078 vp_p.t2822 716.572
R2648 vp_p.n5655 vp_p.t2576 716.572
R2649 vp_p.n4231 vp_p.t1464 716.572
R2650 vp_p.n2806 vp_p.t1050 716.572
R2651 vp_p.n1380 vp_p.t793 716.572
R2652 vp_p.n10126 vp_p.t2650 716.572
R2653 vp_p.n11563 vp_p.t138 716.572
R2654 vp_p.n13001 vp_p.t2018 716.572
R2655 vp_p.n27204 vp_p.t1783 716.572
R2656 vp_p.n25779 vp_p.t1367 716.572
R2657 vp_p.n24357 vp_p.t1123 716.572
R2658 vp_p.n22934 vp_p.t2979 716.572
R2659 vp_p.n21510 vp_p.t460 716.572
R2660 vp_p.n20085 vp_p.t2306 716.572
R2661 vp_p.n18659 vp_p.t1196 716.572
R2662 vp_p.n17232 vp_p.t2674 716.572
R2663 vp_p.n15804 vp_p.t891 716.572
R2664 vp_p.n13178 vp_p.t1595 716.572
R2665 vp_p.n25943 vp_p.t2633 716.572
R2666 vp_p.n24517 vp_p.t2210 716.572
R2667 vp_p.n23095 vp_p.t1997 716.572
R2668 vp_p.n21672 vp_p.t851 716.572
R2669 vp_p.n20248 vp_p.t1335 716.572
R2670 vp_p.n18823 vp_p.t196 716.572
R2671 vp_p.n17397 vp_p.t2067 716.572
R2672 vp_p.n15970 vp_p.t2361 716.572
R2673 vp_p.n14542 vp_p.t1644 716.572
R2674 vp_p.n14381 vp_p.t1266 716.572
R2675 vp_p.n11739 vp_p.t1691 716.572
R2676 vp_p.n8516 vp_p.t721 716.572
R2677 vp_p.n8514 vp_p.t487 716.572
R2678 vp_p.n7092 vp_p.t2942 716.572
R2679 vp_p.n5669 vp_p.t2692 716.572
R2680 vp_p.n4245 vp_p.t1577 716.572
R2681 vp_p.n2820 vp_p.t1166 716.572
R2682 vp_p.n1394 vp_p.t903 716.572
R2683 vp_p.n10140 vp_p.t2750 716.572
R2684 vp_p.n11577 vp_p.t243 716.572
R2685 vp_p.n13017 vp_p.t2118 716.572
R2686 vp_p.n13173 vp_p.t1717 716.572
R2687 vp_p.n27218 vp_p.t2490 716.572
R2688 vp_p.n25793 vp_p.t2090 716.572
R2689 vp_p.n24371 vp_p.t1850 716.572
R2690 vp_p.n22948 vp_p.t704 716.572
R2691 vp_p.n21524 vp_p.t1188 716.572
R2692 vp_p.n20099 vp_p.t41 716.572
R2693 vp_p.n18673 vp_p.t1903 716.572
R2694 vp_p.n17246 vp_p.t2782 716.572
R2695 vp_p.n14537 vp_p.t1619 716.572
R2696 vp_p.n25938 vp_p.t1463 716.572
R2697 vp_p.n24512 vp_p.t1049 716.572
R2698 vp_p.n23090 vp_p.t792 716.572
R2699 vp_p.n21667 vp_p.t2652 716.572
R2700 vp_p.n20243 vp_p.t137 716.572
R2701 vp_p.n18818 vp_p.t2017 716.572
R2702 vp_p.n17392 vp_p.t870 716.572
R2703 vp_p.n15965 vp_p.t689 716.572
R2704 vp_p.n15824 vp_p.t234 716.572
R2705 vp_p.n13168 vp_p.t2565 716.572
R2706 vp_p.n11734 vp_p.t2998 716.572
R2707 vp_p.n10296 vp_p.t1140 716.572
R2708 vp_p.n8530 vp_p.t561 716.572
R2709 vp_p.n8528 vp_p.t293 716.572
R2710 vp_p.n7106 vp_p.t524 716.572
R2711 vp_p.n5683 vp_p.t257 716.572
R2712 vp_p.n4259 vp_p.t2137 716.572
R2713 vp_p.n2834 vp_p.t1728 716.572
R2714 vp_p.n1408 vp_p.t1480 716.572
R2715 vp_p.n10154 vp_p.t332 716.572
R2716 vp_p.n11593 vp_p.t806 716.572
R2717 vp_p.n11729 vp_p.t2666 716.572
R2718 vp_p.n13163 vp_p.t2241 716.572
R2719 vp_p.n14532 vp_p.t992 716.572
R2720 vp_p.n27232 vp_p.t2315 716.572
R2721 vp_p.n25807 vp_p.t1909 716.572
R2722 vp_p.n24385 vp_p.t1678 716.572
R2723 vp_p.n22962 vp_p.t539 716.572
R2724 vp_p.n21538 vp_p.t1013 716.572
R2725 vp_p.n20113 vp_p.t2853 716.572
R2726 vp_p.n18687 vp_p.t1739 716.572
R2727 vp_p.n15960 vp_p.t360 716.572
R2728 vp_p.n25933 vp_p.t259 716.572
R2729 vp_p.n24507 vp_p.t2834 716.572
R2730 vp_p.n23085 vp_p.t2592 716.572
R2731 vp_p.n21662 vp_p.t1483 716.572
R2732 vp_p.n20238 vp_p.t1954 716.572
R2733 vp_p.n18813 vp_p.t809 716.572
R2734 vp_p.n17387 vp_p.t2668 716.572
R2735 vp_p.n17266 vp_p.t2012 716.572
R2736 vp_p.n14527 vp_p.t1854 716.572
R2737 vp_p.n13158 vp_p.t896 716.572
R2738 vp_p.n11724 vp_p.t1321 716.572
R2739 vp_p.n10291 vp_p.t2434 716.572
R2740 vp_p.n8789 vp_p.t1984 716.572
R2741 vp_p.n8544 vp_p.t2358 716.572
R2742 vp_p.n8542 vp_p.t2124 716.572
R2743 vp_p.n7120 vp_p.t1841 716.572
R2744 vp_p.n5697 vp_p.t1594 716.572
R2745 vp_p.n4273 vp_p.t448 716.572
R2746 vp_p.n2848 vp_p.t35 716.572
R2747 vp_p.n1422 vp_p.t2772 716.572
R2748 vp_p.n10170 vp_p.t1661 716.572
R2749 vp_p.n10286 vp_p.t2130 716.572
R2750 vp_p.n11719 vp_p.t991 716.572
R2751 vp_p.n13153 vp_p.t588 716.572
R2752 vp_p.n14522 vp_p.t2574 716.572
R2753 vp_p.n15955 vp_p.t1687 716.572
R2754 vp_p.n27246 vp_p.t1149 716.572
R2755 vp_p.n25821 vp_p.t722 716.572
R2756 vp_p.n24399 vp_p.t489 716.572
R2757 vp_p.n22976 vp_p.t2338 716.572
R2758 vp_p.n21552 vp_p.t2806 716.572
R2759 vp_p.n20127 vp_p.t1693 716.572
R2760 vp_p.n17382 vp_p.t555 716.572
R2761 vp_p.n25928 vp_p.t2340 716.572
R2762 vp_p.n24502 vp_p.t1928 716.572
R2763 vp_p.n23080 vp_p.t1698 716.572
R2764 vp_p.n21657 vp_p.t560 716.572
R2765 vp_p.n20233 vp_p.t1039 716.572
R2766 vp_p.n18808 vp_p.t2876 716.572
R2767 vp_p.n18707 vp_p.t1755 716.572
R2768 vp_p.n15950 vp_p.t338 716.572
R2769 vp_p.n14517 vp_p.t1096 716.572
R2770 vp_p.n13148 vp_p.t2221 716.572
R2771 vp_p.n11714 vp_p.t2643 716.572
R2772 vp_p.n10281 vp_p.t782 716.572
R2773 vp_p.n8784 vp_p.t298 716.572
R2774 vp_p.n45 vp_p.t1451 716.572
R2775 vp_p.n8558 vp_p.t1185 716.572
R2776 vp_p.n8556 vp_p.t925 716.572
R2777 vp_p.n7134 vp_p.t143 716.572
R2778 vp_p.n5711 vp_p.t2885 716.572
R2779 vp_p.n4287 vp_p.t1767 716.572
R2780 vp_p.n2862 vp_p.t1357 716.572
R2781 vp_p.n1438 vp_p.t1104 716.572
R2782 vp_p.n8779 vp_p.t2964 716.572
R2783 vp_p.n10276 vp_p.t445 716.572
R2784 vp_p.n11709 vp_p.t2291 716.572
R2785 vp_p.n13143 vp_p.t1895 716.572
R2786 vp_p.n14512 vp_p.t1203 716.572
R2787 vp_p.n15945 vp_p.t2994 716.572
R2788 vp_p.n17377 vp_p.t2353 716.572
R2789 vp_p.n27260 vp_p.t2946 716.572
R2790 vp_p.n25835 vp_p.t2528 716.572
R2791 vp_p.n24413 vp_p.t2272 716.572
R2792 vp_p.n22990 vp_p.t1168 716.572
R2793 vp_p.n21566 vp_p.t1634 716.572
R2794 vp_p.n18803 vp_p.t505 716.572
R2795 vp_p.n25923 vp_p.t815 716.572
R2796 vp_p.n24497 vp_p.t396 716.572
R2797 vp_p.n23075 vp_p.t163 716.572
R2798 vp_p.n21652 vp_p.t2040 716.572
R2799 vp_p.n20228 vp_p.t2494 716.572
R2800 vp_p.n20147 vp_p.t1369 716.572
R2801 vp_p.n17372 vp_p.t225 716.572
R2802 vp_p.n15940 vp_p.t2662 716.572
R2803 vp_p.n14507 vp_p.t1945 716.572
R2804 vp_p.n13138 vp_p.t1579 716.572
R2805 vp_p.n11704 vp_p.t2001 716.572
R2806 vp_p.n10271 vp_p.t120 716.572
R2807 vp_p.n8774 vp_p.t2632 716.572
R2808 vp_p.n40 vp_p.t775 716.572
R2809 vp_p.n1524 vp_p.t1035 716.572
R2810 vp_p.n8572 vp_p.t1006 716.572
R2811 vp_p.n8570 vp_p.t754 716.572
R2812 vp_p.n7148 vp_p.t711 716.572
R2813 vp_p.n5725 vp_p.t467 716.572
R2814 vp_p.n4301 vp_p.t2314 716.572
R2815 vp_p.n2878 vp_p.t1908 716.572
R2816 vp_p.n35 vp_p.t1677 716.572
R2817 vp_p.n8769 vp_p.t538 716.572
R2818 vp_p.n10266 vp_p.t1012 716.572
R2819 vp_p.n11699 vp_p.t2852 716.572
R2820 vp_p.n13133 vp_p.t2443 716.572
R2821 vp_p.n14502 vp_p.t579 716.572
R2822 vp_p.n15935 vp_p.t566 716.572
R2823 vp_p.n17367 vp_p.t2182 716.572
R2824 vp_p.n18798 vp_p.t317 716.572
R2825 vp_p.n27274 vp_p.t2760 716.572
R2826 vp_p.n25849 vp_p.t2360 716.572
R2827 vp_p.n24427 vp_p.t2123 716.572
R2828 vp_p.n23004 vp_p.t980 716.572
R2829 vp_p.n20223 vp_p.t1469 716.572
R2830 vp_p.n25918 vp_p.t2616 716.572
R2831 vp_p.n24492 vp_p.t2202 716.572
R2832 vp_p.n23070 vp_p.t1983 716.572
R2833 vp_p.n21647 vp_p.t838 716.572
R2834 vp_p.n21586 vp_p.t1320 716.572
R2835 vp_p.n18793 vp_p.t180 716.572
R2836 vp_p.n17362 vp_p.t2052 716.572
R2837 vp_p.n15930 vp_p.t986 716.572
R2838 vp_p.n14497 vp_p.t550 716.572
R2839 vp_p.n13128 vp_p.t2872 716.572
R2840 vp_p.n11694 vp_p.t286 716.572
R2841 vp_p.n10261 vp_p.t1439 716.572
R2842 vp_p.n8764 vp_p.t952 716.572
R2843 vp_p.n30 vp_p.t2103 716.572
R2844 vp_p.n1519 vp_p.t2337 716.572
R2845 vp_p.n2944 vp_p.t2738 716.572
R2846 vp_p.n8586 vp_p.t2075 716.572
R2847 vp_p.n8584 vp_p.t1828 716.572
R2848 vp_p.n7162 vp_p.t2786 716.572
R2849 vp_p.n5739 vp_p.t2542 716.572
R2850 vp_p.n4317 vp_p.t1424 716.572
R2851 vp_p.n1514 vp_p.t1005 716.572
R2852 vp_p.n25 vp_p.t753 716.572
R2853 vp_p.n8759 vp_p.t2606 716.572
R2854 vp_p.n10256 vp_p.t95 716.572
R2855 vp_p.n11689 vp_p.t1976 716.572
R2856 vp_p.n13123 vp_p.t1559 716.572
R2857 vp_p.n14492 vp_p.t2061 716.572
R2858 vp_p.n15925 vp_p.t2639 716.572
R2859 vp_p.n17357 vp_p.t238 716.572
R2860 vp_p.n18788 vp_p.t1394 716.572
R2861 vp_p.n20218 vp_p.t2519 716.572
R2862 vp_p.n27288 vp_p.t842 716.572
R2863 vp_p.n25863 vp_p.t413 716.572
R2864 vp_p.n24441 vp_p.t183 716.572
R2865 vp_p.n21642 vp_p.t2056 716.572
R2866 vp_p.n25913 vp_p.t2449 716.572
R2867 vp_p.n24487 vp_p.t2058 716.572
R2868 vp_p.n23065 vp_p.t1811 716.572
R2869 vp_p.n23024 vp_p.t679 716.572
R2870 vp_p.n20213 vp_p.t1153 716.572
R2871 vp_p.n18783 vp_p.t7 716.572
R2872 vp_p.n17352 vp_p.t1877 716.572
R2873 vp_p.n15920 vp_p.t1562 716.572
R2874 vp_p.n14487 vp_p.t2904 716.572
R2875 vp_p.n13118 vp_p.t449 716.572
R2876 vp_p.n11684 vp_p.t873 716.572
R2877 vp_p.n10251 vp_p.t2016 716.572
R2878 vp_p.n8754 vp_p.t1538 716.572
R2879 vp_p.n20 vp_p.t2651 716.572
R2880 vp_p.n1509 vp_p.t2891 716.572
R2881 vp_p.n2939 vp_p.t312 716.572
R2882 vp_p.n4363 vp_p.t1462 716.572
R2883 vp_p.n8600 vp_p.t882 716.572
R2884 vp_p.n8598 vp_p.t641 716.572
R2885 vp_p.n7176 vp_p.t1122 716.572
R2886 vp_p.n5755 vp_p.t879 716.572
R2887 vp_p.n2934 vp_p.t2718 716.572
R2888 vp_p.n1504 vp_p.t2305 716.572
R2889 vp_p.n15 vp_p.t2086 716.572
R2890 vp_p.n8749 vp_p.t932 716.572
R2891 vp_p.n10246 vp_p.t1419 716.572
R2892 vp_p.n11679 vp_p.t265 716.572
R2893 vp_p.n13113 vp_p.t2844 716.572
R2894 vp_p.n14482 vp_p.t658 716.572
R2895 vp_p.n15915 vp_p.t957 716.572
R2896 vp_p.n17347 vp_p.t2070 716.572
R2897 vp_p.n18778 vp_p.t202 716.572
R2898 vp_p.n20208 vp_p.t1343 716.572
R2899 vp_p.n21637 vp_p.t859 716.572
R2900 vp_p.n27302 vp_p.t2642 716.572
R2901 vp_p.n25877 vp_p.t2219 716.572
R2902 vp_p.n23060 vp_p.t2005 716.572
R2903 vp_p.n25908 vp_p.t1275 716.572
R2904 vp_p.n24482 vp_p.t862 716.572
R2905 vp_p.n24461 vp_p.t627 716.572
R2906 vp_p.n21632 vp_p.t2473 716.572
R2907 vp_p.n20203 vp_p.t2951 716.572
R2908 vp_p.n18773 vp_p.t1826 716.572
R2909 vp_p.n17342 vp_p.t688 716.572
R2910 vp_p.n15910 vp_p.t2849 716.572
R2911 vp_p.n14477 vp_p.t1532 716.572
R2912 vp_p.n13108 vp_p.t1771 716.572
R2913 vp_p.n11674 vp_p.t2175 716.572
R2914 vp_p.n10241 vp_p.t310 716.572
R2915 vp_p.n8744 vp_p.t2825 716.572
R2916 vp_p.n10 vp_p.t971 716.572
R2917 vp_p.n1499 vp_p.t1225 716.572
R2918 vp_p.n2929 vp_p.t1637 716.572
R2919 vp_p.n4358 vp_p.t2752 716.572
R2920 vp_p.n5781 vp_p.t23 716.572
R2921 vp_p.n8614 vp_p.t365 716.572
R2922 vp_p.n8612 vp_p.t119 716.572
R2923 vp_p.n7192 vp_p.t2686 716.572
R2924 vp_p.n4353 vp_p.t2439 716.572
R2925 vp_p.n2924 vp_p.t1324 716.572
R2926 vp_p.n1494 vp_p.t899 716.572
R2927 vp_p.n5 vp_p.t670 716.572
R2928 vp_p.n8739 vp_p.t2518 716.572
R2929 vp_p.n10236 vp_p.t0 716.572
R2930 vp_p.n11669 vp_p.t1870 716.572
R2931 vp_p.n13103 vp_p.t1448 716.572
R2932 vp_p.n14472 vp_p.t2253 716.572
R2933 vp_p.n15905 vp_p.t2535 716.572
R2934 vp_p.n17337 vp_p.t1561 716.572
R2935 vp_p.n18768 vp_p.t2676 716.572
R2936 vp_p.n20198 vp_p.t819 716.572
R2937 vp_p.n21627 vp_p.t346 716.572
R2938 vp_p.n23055 vp_p.t1492 716.572
R2939 vp_p.n27316 vp_p.t2144 716.572
R2940 vp_p.n24477 vp_p.t1734 716.572
R2941 vp_p.n25903 vp_p.t2322 716.572
R2942 vp_p.n25897 vp_p.t1916 716.572
R2943 vp_p.n23050 vp_p.t1684 716.572
R2944 vp_p.n21622 vp_p.t544 716.572
R2945 vp_p.n20193 vp_p.t1019 716.572
R2946 vp_p.n18763 vp_p.t2861 716.572
R2947 vp_p.n17332 vp_p.t1746 716.572
R2948 vp_p.n15900 vp_p.t1969 716.572
R2949 vp_p.n14467 vp_p.t2 716.572
R2950 vp_p.n13098 vp_p.t864 716.572
R2951 vp_p.n11664 vp_p.t1276 716.572
R2952 vp_p.n10231 vp_p.t2396 716.572
R2953 vp_p.n8734 vp_p.t1939 716.572
R2954 vp_p.n0 vp_p.t73 716.572
R2955 vp_p.n1489 vp_p.t304 716.572
R2956 vp_p.n2919 vp_p.t730 716.572
R2957 vp_p.n4348 vp_p.t1876 716.572
R2958 vp_p.n5776 vp_p.t2115 716.572
R2959 vp_p.n8622 vp_p.t302 716.572
R2960 vp_p.n7580 vp_p.t435 716.572
R2961 vp_p.n7582 vp_p.t203 716.572
R2962 vp_p.n6146 vp_p.t182 716.572
R2963 vp_p.n4723 vp_p.t2926 716.572
R2964 vp_p.n3299 vp_p.t1804 716.572
R2965 vp_p.n1874 vp_p.t1390 716.572
R2966 vp_p.n390 vp_p.t1147 716.572
R2967 vp_p.n9129 vp_p.t4 716.572
R2968 vp_p.n10631 vp_p.t488 716.572
R2969 vp_p.n12069 vp_p.t2336 716.572
R2970 vp_p.n13833 vp_p.t1924 716.572
R2971 vp_p.n14872 vp_p.t2189 716.572
R2972 vp_p.n16300 vp_p.t31 716.572
R2973 vp_p.n17727 vp_p.t1622 716.572
R2974 vp_p.n19153 vp_p.t2741 716.572
R2975 vp_p.n20578 vp_p.t898 716.572
R2976 vp_p.n22002 vp_p.t410 716.572
R2977 vp_p.n23425 vp_p.t1568 716.572
R2978 vp_p.n24847 vp_p.t1805 716.572
R2979 vp_p.n26273 vp_p.t2203 716.572
R2980 vp_p.n26280 vp_p.t1017 716.572
R2981 vp_p.n24852 vp_p.t605 716.572
R2982 vp_p.n23430 vp_p.t349 716.572
R2983 vp_p.n22007 vp_p.t2201 716.572
R2984 vp_p.n20583 vp_p.t2680 716.572
R2985 vp_p.n19158 vp_p.t1564 716.572
R2986 vp_p.n17732 vp_p.t407 716.572
R2987 vp_p.n16305 vp_p.t1370 716.572
R2988 vp_p.n14877 vp_p.t698 716.572
R2989 vp_p.n13838 vp_p.t252 716.572
R2990 vp_p.n12074 vp_p.t685 716.572
R2991 vp_p.n10636 vp_p.t1823 716.572
R2992 vp_p.n9134 vp_p.t1352 716.572
R2993 vp_p.n395 vp_p.t2472 716.572
R2994 vp_p.n1879 vp_p.t2704 716.572
R2995 vp_p.n3304 vp_p.t131 716.572
R2996 vp_p.n4728 vp_p.t1274 716.572
R2997 vp_p.n6151 vp_p.t1528 716.572
R2998 vp_p.n7568 vp_p.t2003 716.572
R2999 vp_p.n7570 vp_p.t2217 716.572
R3000 vp_p.n14383 vp_p.n14380 18.301
R3001 vp_p.n13019 vp_p.n13016 18.301
R3002 vp_p.n15826 vp_p.n15823 18.301
R3003 vp_p.n11595 vp_p.n11592 18.301
R3004 vp_p.n17268 vp_p.n17265 18.301
R3005 vp_p.n10172 vp_p.n10169 18.301
R3006 vp_p.n18709 vp_p.n18706 18.301
R3007 vp_p.n1440 vp_p.n1437 18.301
R3008 vp_p.n20149 vp_p.n20146 18.301
R3009 vp_p.n2880 vp_p.n2877 18.301
R3010 vp_p.n21588 vp_p.n21585 18.301
R3011 vp_p.n4319 vp_p.n4316 18.301
R3012 vp_p.n23026 vp_p.n23023 18.301
R3013 vp_p.n5757 vp_p.n5754 18.301
R3014 vp_p.n24463 vp_p.n24460 18.301
R3015 vp_p.n7194 vp_p.n7191 18.301
R3016 vp_p.n25899 vp_p.n25896 18.301
R3017 vp_p.n7584 vp_p.n7581 18.301
R3018 vp_p.n7572 vp_p.n7571 18.301
R3019 vp_p.n24856 vp_p.n24855 18.301
R3020 vp_p.n24851 vp_p.n24850 18.301
R3021 vp_p.n6155 vp_p.n6154 18.301
R3022 vp_p.n6150 vp_p.n6149 18.301
R3023 vp_p.n23434 vp_p.n23433 18.301
R3024 vp_p.n23429 vp_p.n23428 18.301
R3025 vp_p.n4732 vp_p.n4731 18.301
R3026 vp_p.n4727 vp_p.n4726 18.301
R3027 vp_p.n22011 vp_p.n22010 18.301
R3028 vp_p.n22006 vp_p.n22005 18.301
R3029 vp_p.n3308 vp_p.n3307 18.301
R3030 vp_p.n3303 vp_p.n3302 18.301
R3031 vp_p.n20587 vp_p.n20586 18.301
R3032 vp_p.n20582 vp_p.n20581 18.301
R3033 vp_p.n1883 vp_p.n1882 18.301
R3034 vp_p.n1878 vp_p.n1877 18.301
R3035 vp_p.n19162 vp_p.n19161 18.301
R3036 vp_p.n19157 vp_p.n19156 18.301
R3037 vp_p.n399 vp_p.n398 18.301
R3038 vp_p.n394 vp_p.n393 18.301
R3039 vp_p.n17736 vp_p.n17735 18.301
R3040 vp_p.n17731 vp_p.n17730 18.301
R3041 vp_p.n9138 vp_p.n9137 18.301
R3042 vp_p.n9133 vp_p.n9132 18.301
R3043 vp_p.n16309 vp_p.n16308 18.301
R3044 vp_p.n16304 vp_p.n16303 18.301
R3045 vp_p.n10640 vp_p.n10639 18.301
R3046 vp_p.n10635 vp_p.n10634 18.301
R3047 vp_p.n14881 vp_p.n14880 18.301
R3048 vp_p.n14876 vp_p.n14875 18.301
R3049 vp_p.n12078 vp_p.n12077 18.301
R3050 vp_p.n12073 vp_p.n12072 18.301
R3051 vp_p.n13842 vp_p.n13841 18.301
R3052 vp_p.n13837 vp_p.n13836 18.301
R3053 vp_p.n13177 vp_p.n13176 18.301
R3054 vp_p.n13172 vp_p.n13171 18.301
R3055 vp_p.n13167 vp_p.n13166 18.301
R3056 vp_p.n13162 vp_p.n13161 18.301
R3057 vp_p.n13157 vp_p.n13156 18.301
R3058 vp_p.n13152 vp_p.n13151 18.301
R3059 vp_p.n13147 vp_p.n13146 18.301
R3060 vp_p.n13142 vp_p.n13141 18.301
R3061 vp_p.n13137 vp_p.n13136 18.301
R3062 vp_p.n13132 vp_p.n13131 18.301
R3063 vp_p.n13127 vp_p.n13126 18.301
R3064 vp_p.n13122 vp_p.n13121 18.301
R3065 vp_p.n13117 vp_p.n13116 18.301
R3066 vp_p.n13112 vp_p.n13111 18.301
R3067 vp_p.n13107 vp_p.n13106 18.301
R3068 vp_p.n13102 vp_p.n13101 18.301
R3069 vp_p.n11738 vp_p.n11737 18.301
R3070 vp_p.n11733 vp_p.n11732 18.301
R3071 vp_p.n11728 vp_p.n11727 18.301
R3072 vp_p.n11723 vp_p.n11722 18.301
R3073 vp_p.n11718 vp_p.n11717 18.301
R3074 vp_p.n11713 vp_p.n11712 18.301
R3075 vp_p.n11708 vp_p.n11707 18.301
R3076 vp_p.n11703 vp_p.n11702 18.301
R3077 vp_p.n11698 vp_p.n11697 18.301
R3078 vp_p.n11693 vp_p.n11692 18.301
R3079 vp_p.n11688 vp_p.n11687 18.301
R3080 vp_p.n11683 vp_p.n11682 18.301
R3081 vp_p.n11678 vp_p.n11677 18.301
R3082 vp_p.n11673 vp_p.n11672 18.301
R3083 vp_p.n11668 vp_p.n11667 18.301
R3084 vp_p.n14536 vp_p.n14535 18.301
R3085 vp_p.n14531 vp_p.n14530 18.301
R3086 vp_p.n14526 vp_p.n14525 18.301
R3087 vp_p.n14521 vp_p.n14520 18.301
R3088 vp_p.n14516 vp_p.n14515 18.301
R3089 vp_p.n14511 vp_p.n14510 18.301
R3090 vp_p.n14506 vp_p.n14505 18.301
R3091 vp_p.n14501 vp_p.n14500 18.301
R3092 vp_p.n14496 vp_p.n14495 18.301
R3093 vp_p.n14491 vp_p.n14490 18.301
R3094 vp_p.n14486 vp_p.n14485 18.301
R3095 vp_p.n14481 vp_p.n14480 18.301
R3096 vp_p.n14476 vp_p.n14475 18.301
R3097 vp_p.n14471 vp_p.n14470 18.301
R3098 vp_p.n10295 vp_p.n10294 18.301
R3099 vp_p.n10290 vp_p.n10289 18.301
R3100 vp_p.n10285 vp_p.n10284 18.301
R3101 vp_p.n10280 vp_p.n10279 18.301
R3102 vp_p.n10275 vp_p.n10274 18.301
R3103 vp_p.n10270 vp_p.n10269 18.301
R3104 vp_p.n10265 vp_p.n10264 18.301
R3105 vp_p.n10260 vp_p.n10259 18.301
R3106 vp_p.n10255 vp_p.n10254 18.301
R3107 vp_p.n10250 vp_p.n10249 18.301
R3108 vp_p.n10245 vp_p.n10244 18.301
R3109 vp_p.n10240 vp_p.n10239 18.301
R3110 vp_p.n10235 vp_p.n10234 18.301
R3111 vp_p.n15959 vp_p.n15958 18.301
R3112 vp_p.n15954 vp_p.n15953 18.301
R3113 vp_p.n15949 vp_p.n15948 18.301
R3114 vp_p.n15944 vp_p.n15943 18.301
R3115 vp_p.n15939 vp_p.n15938 18.301
R3116 vp_p.n15934 vp_p.n15933 18.301
R3117 vp_p.n15929 vp_p.n15928 18.301
R3118 vp_p.n15924 vp_p.n15923 18.301
R3119 vp_p.n15919 vp_p.n15918 18.301
R3120 vp_p.n15914 vp_p.n15913 18.301
R3121 vp_p.n15909 vp_p.n15908 18.301
R3122 vp_p.n15904 vp_p.n15903 18.301
R3123 vp_p.n8788 vp_p.n8787 18.301
R3124 vp_p.n8783 vp_p.n8782 18.301
R3125 vp_p.n8778 vp_p.n8777 18.301
R3126 vp_p.n8773 vp_p.n8772 18.301
R3127 vp_p.n8768 vp_p.n8767 18.301
R3128 vp_p.n8763 vp_p.n8762 18.301
R3129 vp_p.n8758 vp_p.n8757 18.301
R3130 vp_p.n8753 vp_p.n8752 18.301
R3131 vp_p.n8748 vp_p.n8747 18.301
R3132 vp_p.n8743 vp_p.n8742 18.301
R3133 vp_p.n8738 vp_p.n8737 18.301
R3134 vp_p.n17381 vp_p.n17380 18.301
R3135 vp_p.n17376 vp_p.n17375 18.301
R3136 vp_p.n17371 vp_p.n17370 18.301
R3137 vp_p.n17366 vp_p.n17365 18.301
R3138 vp_p.n17361 vp_p.n17360 18.301
R3139 vp_p.n17356 vp_p.n17355 18.301
R3140 vp_p.n17351 vp_p.n17350 18.301
R3141 vp_p.n17346 vp_p.n17345 18.301
R3142 vp_p.n17341 vp_p.n17340 18.301
R3143 vp_p.n17336 vp_p.n17335 18.301
R3144 vp_p.n44 vp_p.n43 18.301
R3145 vp_p.n39 vp_p.n38 18.301
R3146 vp_p.n34 vp_p.n33 18.301
R3147 vp_p.n29 vp_p.n28 18.301
R3148 vp_p.n24 vp_p.n23 18.301
R3149 vp_p.n19 vp_p.n18 18.301
R3150 vp_p.n14 vp_p.n13 18.301
R3151 vp_p.n9 vp_p.n8 18.301
R3152 vp_p.n4 vp_p.n3 18.301
R3153 vp_p.n18802 vp_p.n18801 18.301
R3154 vp_p.n18797 vp_p.n18796 18.301
R3155 vp_p.n18792 vp_p.n18791 18.301
R3156 vp_p.n18787 vp_p.n18786 18.301
R3157 vp_p.n18782 vp_p.n18781 18.301
R3158 vp_p.n18777 vp_p.n18776 18.301
R3159 vp_p.n18772 vp_p.n18771 18.301
R3160 vp_p.n18767 vp_p.n18766 18.301
R3161 vp_p.n1523 vp_p.n1522 18.301
R3162 vp_p.n1518 vp_p.n1517 18.301
R3163 vp_p.n1513 vp_p.n1512 18.301
R3164 vp_p.n1508 vp_p.n1507 18.301
R3165 vp_p.n1503 vp_p.n1502 18.301
R3166 vp_p.n1498 vp_p.n1497 18.301
R3167 vp_p.n1493 vp_p.n1492 18.301
R3168 vp_p.n20222 vp_p.n20221 18.301
R3169 vp_p.n20217 vp_p.n20216 18.301
R3170 vp_p.n20212 vp_p.n20211 18.301
R3171 vp_p.n20207 vp_p.n20206 18.301
R3172 vp_p.n20202 vp_p.n20201 18.301
R3173 vp_p.n20197 vp_p.n20196 18.301
R3174 vp_p.n2943 vp_p.n2942 18.301
R3175 vp_p.n2938 vp_p.n2937 18.301
R3176 vp_p.n2933 vp_p.n2932 18.301
R3177 vp_p.n2928 vp_p.n2927 18.301
R3178 vp_p.n2923 vp_p.n2922 18.301
R3179 vp_p.n21641 vp_p.n21640 18.301
R3180 vp_p.n21636 vp_p.n21635 18.301
R3181 vp_p.n21631 vp_p.n21630 18.301
R3182 vp_p.n21626 vp_p.n21625 18.301
R3183 vp_p.n4362 vp_p.n4361 18.301
R3184 vp_p.n4357 vp_p.n4356 18.301
R3185 vp_p.n4352 vp_p.n4351 18.301
R3186 vp_p.n23059 vp_p.n23058 18.301
R3187 vp_p.n23054 vp_p.n23053 18.301
R3188 vp_p.n5780 vp_p.n5779 18.301
R3189 vp_p.n8626 vp_p.n8625 18.301
R3190 vp_p.n12095 vp_p.n12094 18.301
R3191 vp_p.n10657 vp_p.n10656 18.301
R3192 vp_p.n9220 vp_p.n9219 18.301
R3193 vp_p.n474 vp_p.n473 18.301
R3194 vp_p.n1900 vp_p.n1899 18.301
R3195 vp_p.n3325 vp_p.n3324 18.301
R3196 vp_p.n4749 vp_p.n4748 18.301
R3197 vp_p.n6172 vp_p.n6171 18.301
R3198 vp_p.n7594 vp_p.n7593 18.301
R3199 vp_p.n14898 vp_p.n14897 18.301
R3200 vp_p.n16326 vp_p.n16325 18.301
R3201 vp_p.n17753 vp_p.n17752 18.301
R3202 vp_p.n19179 vp_p.n19178 18.301
R3203 vp_p.n20604 vp_p.n20603 18.301
R3204 vp_p.n22028 vp_p.n22027 18.301
R3205 vp_p.n23451 vp_p.n23450 18.301
R3206 vp_p.n24873 vp_p.n24872 18.301
R3207 vp_p.n26298 vp_p.n26297 18.301
R3208 vp_p.n12109 vp_p.n12108 18.301
R3209 vp_p.n10671 vp_p.n10670 18.301
R3210 vp_p.n9234 vp_p.n9233 18.301
R3211 vp_p.n488 vp_p.n487 18.301
R3212 vp_p.n1914 vp_p.n1913 18.301
R3213 vp_p.n3339 vp_p.n3338 18.301
R3214 vp_p.n4763 vp_p.n4762 18.301
R3215 vp_p.n6186 vp_p.n6185 18.301
R3216 vp_p.n7608 vp_p.n7607 18.301
R3217 vp_p.n14912 vp_p.n14911 18.301
R3218 vp_p.n16340 vp_p.n16339 18.301
R3219 vp_p.n17767 vp_p.n17766 18.301
R3220 vp_p.n19193 vp_p.n19192 18.301
R3221 vp_p.n20618 vp_p.n20617 18.301
R3222 vp_p.n22042 vp_p.n22041 18.301
R3223 vp_p.n23465 vp_p.n23464 18.301
R3224 vp_p.n24887 vp_p.n24886 18.301
R3225 vp_p.n26312 vp_p.n26311 18.301
R3226 vp_p.n12123 vp_p.n12122 18.301
R3227 vp_p.n10685 vp_p.n10684 18.301
R3228 vp_p.n9248 vp_p.n9247 18.301
R3229 vp_p.n502 vp_p.n501 18.301
R3230 vp_p.n1928 vp_p.n1927 18.301
R3231 vp_p.n3353 vp_p.n3352 18.301
R3232 vp_p.n4777 vp_p.n4776 18.301
R3233 vp_p.n6200 vp_p.n6199 18.301
R3234 vp_p.n7622 vp_p.n7621 18.301
R3235 vp_p.n14926 vp_p.n14925 18.301
R3236 vp_p.n16354 vp_p.n16353 18.301
R3237 vp_p.n17781 vp_p.n17780 18.301
R3238 vp_p.n19207 vp_p.n19206 18.301
R3239 vp_p.n20632 vp_p.n20631 18.301
R3240 vp_p.n22056 vp_p.n22055 18.301
R3241 vp_p.n23479 vp_p.n23478 18.301
R3242 vp_p.n24901 vp_p.n24900 18.301
R3243 vp_p.n26326 vp_p.n26325 18.301
R3244 vp_p.n12137 vp_p.n12136 18.301
R3245 vp_p.n10699 vp_p.n10698 18.301
R3246 vp_p.n9262 vp_p.n9261 18.301
R3247 vp_p.n516 vp_p.n515 18.301
R3248 vp_p.n1942 vp_p.n1941 18.301
R3249 vp_p.n3367 vp_p.n3366 18.301
R3250 vp_p.n4791 vp_p.n4790 18.301
R3251 vp_p.n6214 vp_p.n6213 18.301
R3252 vp_p.n7636 vp_p.n7635 18.301
R3253 vp_p.n14940 vp_p.n14939 18.301
R3254 vp_p.n16368 vp_p.n16367 18.301
R3255 vp_p.n17795 vp_p.n17794 18.301
R3256 vp_p.n19221 vp_p.n19220 18.301
R3257 vp_p.n20646 vp_p.n20645 18.301
R3258 vp_p.n22070 vp_p.n22069 18.301
R3259 vp_p.n23493 vp_p.n23492 18.301
R3260 vp_p.n24915 vp_p.n24914 18.301
R3261 vp_p.n26340 vp_p.n26339 18.301
R3262 vp_p.n12151 vp_p.n12150 18.301
R3263 vp_p.n10713 vp_p.n10712 18.301
R3264 vp_p.n9276 vp_p.n9275 18.301
R3265 vp_p.n530 vp_p.n529 18.301
R3266 vp_p.n1956 vp_p.n1955 18.301
R3267 vp_p.n3381 vp_p.n3380 18.301
R3268 vp_p.n4805 vp_p.n4804 18.301
R3269 vp_p.n6228 vp_p.n6227 18.301
R3270 vp_p.n7650 vp_p.n7649 18.301
R3271 vp_p.n14954 vp_p.n14953 18.301
R3272 vp_p.n16382 vp_p.n16381 18.301
R3273 vp_p.n17809 vp_p.n17808 18.301
R3274 vp_p.n19235 vp_p.n19234 18.301
R3275 vp_p.n20660 vp_p.n20659 18.301
R3276 vp_p.n22084 vp_p.n22083 18.301
R3277 vp_p.n23507 vp_p.n23506 18.301
R3278 vp_p.n24929 vp_p.n24928 18.301
R3279 vp_p.n26354 vp_p.n26353 18.301
R3280 vp_p.n12165 vp_p.n12164 18.301
R3281 vp_p.n10727 vp_p.n10726 18.301
R3282 vp_p.n9290 vp_p.n9289 18.301
R3283 vp_p.n544 vp_p.n543 18.301
R3284 vp_p.n1970 vp_p.n1969 18.301
R3285 vp_p.n3395 vp_p.n3394 18.301
R3286 vp_p.n4819 vp_p.n4818 18.301
R3287 vp_p.n6242 vp_p.n6241 18.301
R3288 vp_p.n7664 vp_p.n7663 18.301
R3289 vp_p.n14968 vp_p.n14967 18.301
R3290 vp_p.n16396 vp_p.n16395 18.301
R3291 vp_p.n17823 vp_p.n17822 18.301
R3292 vp_p.n19249 vp_p.n19248 18.301
R3293 vp_p.n20674 vp_p.n20673 18.301
R3294 vp_p.n22098 vp_p.n22097 18.301
R3295 vp_p.n23521 vp_p.n23520 18.301
R3296 vp_p.n24943 vp_p.n24942 18.301
R3297 vp_p.n26368 vp_p.n26367 18.301
R3298 vp_p.n12179 vp_p.n12178 18.301
R3299 vp_p.n10741 vp_p.n10740 18.301
R3300 vp_p.n9304 vp_p.n9303 18.301
R3301 vp_p.n558 vp_p.n557 18.301
R3302 vp_p.n1984 vp_p.n1983 18.301
R3303 vp_p.n3409 vp_p.n3408 18.301
R3304 vp_p.n4833 vp_p.n4832 18.301
R3305 vp_p.n6256 vp_p.n6255 18.301
R3306 vp_p.n7678 vp_p.n7677 18.301
R3307 vp_p.n14982 vp_p.n14981 18.301
R3308 vp_p.n16410 vp_p.n16409 18.301
R3309 vp_p.n17837 vp_p.n17836 18.301
R3310 vp_p.n19263 vp_p.n19262 18.301
R3311 vp_p.n20688 vp_p.n20687 18.301
R3312 vp_p.n22112 vp_p.n22111 18.301
R3313 vp_p.n23535 vp_p.n23534 18.301
R3314 vp_p.n24957 vp_p.n24956 18.301
R3315 vp_p.n26382 vp_p.n26381 18.301
R3316 vp_p.n12193 vp_p.n12192 18.301
R3317 vp_p.n10755 vp_p.n10754 18.301
R3318 vp_p.n9318 vp_p.n9317 18.301
R3319 vp_p.n572 vp_p.n571 18.301
R3320 vp_p.n1998 vp_p.n1997 18.301
R3321 vp_p.n3423 vp_p.n3422 18.301
R3322 vp_p.n4847 vp_p.n4846 18.301
R3323 vp_p.n6270 vp_p.n6269 18.301
R3324 vp_p.n7692 vp_p.n7691 18.301
R3325 vp_p.n14996 vp_p.n14995 18.301
R3326 vp_p.n16424 vp_p.n16423 18.301
R3327 vp_p.n17851 vp_p.n17850 18.301
R3328 vp_p.n19277 vp_p.n19276 18.301
R3329 vp_p.n20702 vp_p.n20701 18.301
R3330 vp_p.n22126 vp_p.n22125 18.301
R3331 vp_p.n23549 vp_p.n23548 18.301
R3332 vp_p.n24971 vp_p.n24970 18.301
R3333 vp_p.n26396 vp_p.n26395 18.301
R3334 vp_p.n12207 vp_p.n12206 18.301
R3335 vp_p.n10769 vp_p.n10768 18.301
R3336 vp_p.n9332 vp_p.n9331 18.301
R3337 vp_p.n586 vp_p.n585 18.301
R3338 vp_p.n2012 vp_p.n2011 18.301
R3339 vp_p.n3437 vp_p.n3436 18.301
R3340 vp_p.n4861 vp_p.n4860 18.301
R3341 vp_p.n6284 vp_p.n6283 18.301
R3342 vp_p.n7706 vp_p.n7705 18.301
R3343 vp_p.n15010 vp_p.n15009 18.301
R3344 vp_p.n16438 vp_p.n16437 18.301
R3345 vp_p.n17865 vp_p.n17864 18.301
R3346 vp_p.n19291 vp_p.n19290 18.301
R3347 vp_p.n20716 vp_p.n20715 18.301
R3348 vp_p.n22140 vp_p.n22139 18.301
R3349 vp_p.n23563 vp_p.n23562 18.301
R3350 vp_p.n24985 vp_p.n24984 18.301
R3351 vp_p.n26410 vp_p.n26409 18.301
R3352 vp_p.n12221 vp_p.n12220 18.301
R3353 vp_p.n10783 vp_p.n10782 18.301
R3354 vp_p.n9346 vp_p.n9345 18.301
R3355 vp_p.n600 vp_p.n599 18.301
R3356 vp_p.n2026 vp_p.n2025 18.301
R3357 vp_p.n3451 vp_p.n3450 18.301
R3358 vp_p.n4875 vp_p.n4874 18.301
R3359 vp_p.n6298 vp_p.n6297 18.301
R3360 vp_p.n7720 vp_p.n7719 18.301
R3361 vp_p.n15024 vp_p.n15023 18.301
R3362 vp_p.n16452 vp_p.n16451 18.301
R3363 vp_p.n17879 vp_p.n17878 18.301
R3364 vp_p.n19305 vp_p.n19304 18.301
R3365 vp_p.n20730 vp_p.n20729 18.301
R3366 vp_p.n22154 vp_p.n22153 18.301
R3367 vp_p.n23577 vp_p.n23576 18.301
R3368 vp_p.n24999 vp_p.n24998 18.301
R3369 vp_p.n26424 vp_p.n26423 18.301
R3370 vp_p.n12235 vp_p.n12234 18.301
R3371 vp_p.n10797 vp_p.n10796 18.301
R3372 vp_p.n9360 vp_p.n9359 18.301
R3373 vp_p.n614 vp_p.n613 18.301
R3374 vp_p.n2040 vp_p.n2039 18.301
R3375 vp_p.n3465 vp_p.n3464 18.301
R3376 vp_p.n4889 vp_p.n4888 18.301
R3377 vp_p.n6312 vp_p.n6311 18.301
R3378 vp_p.n7734 vp_p.n7733 18.301
R3379 vp_p.n15038 vp_p.n15037 18.301
R3380 vp_p.n16466 vp_p.n16465 18.301
R3381 vp_p.n17893 vp_p.n17892 18.301
R3382 vp_p.n19319 vp_p.n19318 18.301
R3383 vp_p.n20744 vp_p.n20743 18.301
R3384 vp_p.n22168 vp_p.n22167 18.301
R3385 vp_p.n23591 vp_p.n23590 18.301
R3386 vp_p.n25013 vp_p.n25012 18.301
R3387 vp_p.n26438 vp_p.n26437 18.301
R3388 vp_p.n12249 vp_p.n12248 18.301
R3389 vp_p.n10811 vp_p.n10810 18.301
R3390 vp_p.n9374 vp_p.n9373 18.301
R3391 vp_p.n628 vp_p.n627 18.301
R3392 vp_p.n2054 vp_p.n2053 18.301
R3393 vp_p.n3479 vp_p.n3478 18.301
R3394 vp_p.n4903 vp_p.n4902 18.301
R3395 vp_p.n6326 vp_p.n6325 18.301
R3396 vp_p.n7748 vp_p.n7747 18.301
R3397 vp_p.n15052 vp_p.n15051 18.301
R3398 vp_p.n16480 vp_p.n16479 18.301
R3399 vp_p.n17907 vp_p.n17906 18.301
R3400 vp_p.n19333 vp_p.n19332 18.301
R3401 vp_p.n20758 vp_p.n20757 18.301
R3402 vp_p.n22182 vp_p.n22181 18.301
R3403 vp_p.n23605 vp_p.n23604 18.301
R3404 vp_p.n25027 vp_p.n25026 18.301
R3405 vp_p.n26452 vp_p.n26451 18.301
R3406 vp_p.n12263 vp_p.n12262 18.301
R3407 vp_p.n10825 vp_p.n10824 18.301
R3408 vp_p.n9388 vp_p.n9387 18.301
R3409 vp_p.n642 vp_p.n641 18.301
R3410 vp_p.n2068 vp_p.n2067 18.301
R3411 vp_p.n3493 vp_p.n3492 18.301
R3412 vp_p.n4917 vp_p.n4916 18.301
R3413 vp_p.n6340 vp_p.n6339 18.301
R3414 vp_p.n7762 vp_p.n7761 18.301
R3415 vp_p.n15066 vp_p.n15065 18.301
R3416 vp_p.n16494 vp_p.n16493 18.301
R3417 vp_p.n17921 vp_p.n17920 18.301
R3418 vp_p.n19347 vp_p.n19346 18.301
R3419 vp_p.n20772 vp_p.n20771 18.301
R3420 vp_p.n22196 vp_p.n22195 18.301
R3421 vp_p.n23619 vp_p.n23618 18.301
R3422 vp_p.n25041 vp_p.n25040 18.301
R3423 vp_p.n26466 vp_p.n26465 18.301
R3424 vp_p.n12277 vp_p.n12276 18.301
R3425 vp_p.n10839 vp_p.n10838 18.301
R3426 vp_p.n9402 vp_p.n9401 18.301
R3427 vp_p.n656 vp_p.n655 18.301
R3428 vp_p.n2082 vp_p.n2081 18.301
R3429 vp_p.n3507 vp_p.n3506 18.301
R3430 vp_p.n4931 vp_p.n4930 18.301
R3431 vp_p.n6354 vp_p.n6353 18.301
R3432 vp_p.n7776 vp_p.n7775 18.301
R3433 vp_p.n15080 vp_p.n15079 18.301
R3434 vp_p.n16508 vp_p.n16507 18.301
R3435 vp_p.n17935 vp_p.n17934 18.301
R3436 vp_p.n19361 vp_p.n19360 18.301
R3437 vp_p.n20786 vp_p.n20785 18.301
R3438 vp_p.n22210 vp_p.n22209 18.301
R3439 vp_p.n23633 vp_p.n23632 18.301
R3440 vp_p.n25055 vp_p.n25054 18.301
R3441 vp_p.n26480 vp_p.n26479 18.301
R3442 vp_p.n12291 vp_p.n12290 18.301
R3443 vp_p.n10853 vp_p.n10852 18.301
R3444 vp_p.n9416 vp_p.n9415 18.301
R3445 vp_p.n670 vp_p.n669 18.301
R3446 vp_p.n2096 vp_p.n2095 18.301
R3447 vp_p.n3521 vp_p.n3520 18.301
R3448 vp_p.n4945 vp_p.n4944 18.301
R3449 vp_p.n6368 vp_p.n6367 18.301
R3450 vp_p.n7790 vp_p.n7789 18.301
R3451 vp_p.n15094 vp_p.n15093 18.301
R3452 vp_p.n16522 vp_p.n16521 18.301
R3453 vp_p.n17949 vp_p.n17948 18.301
R3454 vp_p.n19375 vp_p.n19374 18.301
R3455 vp_p.n20800 vp_p.n20799 18.301
R3456 vp_p.n22224 vp_p.n22223 18.301
R3457 vp_p.n23647 vp_p.n23646 18.301
R3458 vp_p.n25069 vp_p.n25068 18.301
R3459 vp_p.n26494 vp_p.n26493 18.301
R3460 vp_p.n12305 vp_p.n12304 18.301
R3461 vp_p.n10867 vp_p.n10866 18.301
R3462 vp_p.n9430 vp_p.n9429 18.301
R3463 vp_p.n684 vp_p.n683 18.301
R3464 vp_p.n2110 vp_p.n2109 18.301
R3465 vp_p.n3535 vp_p.n3534 18.301
R3466 vp_p.n4959 vp_p.n4958 18.301
R3467 vp_p.n6382 vp_p.n6381 18.301
R3468 vp_p.n7804 vp_p.n7803 18.301
R3469 vp_p.n15108 vp_p.n15107 18.301
R3470 vp_p.n16536 vp_p.n16535 18.301
R3471 vp_p.n17963 vp_p.n17962 18.301
R3472 vp_p.n19389 vp_p.n19388 18.301
R3473 vp_p.n20814 vp_p.n20813 18.301
R3474 vp_p.n22238 vp_p.n22237 18.301
R3475 vp_p.n23661 vp_p.n23660 18.301
R3476 vp_p.n25083 vp_p.n25082 18.301
R3477 vp_p.n26508 vp_p.n26507 18.301
R3478 vp_p.n12319 vp_p.n12318 18.301
R3479 vp_p.n10881 vp_p.n10880 18.301
R3480 vp_p.n9444 vp_p.n9443 18.301
R3481 vp_p.n698 vp_p.n697 18.301
R3482 vp_p.n2124 vp_p.n2123 18.301
R3483 vp_p.n3549 vp_p.n3548 18.301
R3484 vp_p.n4973 vp_p.n4972 18.301
R3485 vp_p.n6396 vp_p.n6395 18.301
R3486 vp_p.n7818 vp_p.n7817 18.301
R3487 vp_p.n15122 vp_p.n15121 18.301
R3488 vp_p.n16550 vp_p.n16549 18.301
R3489 vp_p.n17977 vp_p.n17976 18.301
R3490 vp_p.n19403 vp_p.n19402 18.301
R3491 vp_p.n20828 vp_p.n20827 18.301
R3492 vp_p.n22252 vp_p.n22251 18.301
R3493 vp_p.n23675 vp_p.n23674 18.301
R3494 vp_p.n25097 vp_p.n25096 18.301
R3495 vp_p.n26522 vp_p.n26521 18.301
R3496 vp_p.n12333 vp_p.n12332 18.301
R3497 vp_p.n10895 vp_p.n10894 18.301
R3498 vp_p.n9458 vp_p.n9457 18.301
R3499 vp_p.n712 vp_p.n711 18.301
R3500 vp_p.n2138 vp_p.n2137 18.301
R3501 vp_p.n3563 vp_p.n3562 18.301
R3502 vp_p.n4987 vp_p.n4986 18.301
R3503 vp_p.n6410 vp_p.n6409 18.301
R3504 vp_p.n7832 vp_p.n7831 18.301
R3505 vp_p.n15136 vp_p.n15135 18.301
R3506 vp_p.n16564 vp_p.n16563 18.301
R3507 vp_p.n17991 vp_p.n17990 18.301
R3508 vp_p.n19417 vp_p.n19416 18.301
R3509 vp_p.n20842 vp_p.n20841 18.301
R3510 vp_p.n22266 vp_p.n22265 18.301
R3511 vp_p.n23689 vp_p.n23688 18.301
R3512 vp_p.n25111 vp_p.n25110 18.301
R3513 vp_p.n26536 vp_p.n26535 18.301
R3514 vp_p.n12347 vp_p.n12346 18.301
R3515 vp_p.n10909 vp_p.n10908 18.301
R3516 vp_p.n9472 vp_p.n9471 18.301
R3517 vp_p.n726 vp_p.n725 18.301
R3518 vp_p.n2152 vp_p.n2151 18.301
R3519 vp_p.n3577 vp_p.n3576 18.301
R3520 vp_p.n5001 vp_p.n5000 18.301
R3521 vp_p.n6424 vp_p.n6423 18.301
R3522 vp_p.n7846 vp_p.n7845 18.301
R3523 vp_p.n15150 vp_p.n15149 18.301
R3524 vp_p.n16578 vp_p.n16577 18.301
R3525 vp_p.n18005 vp_p.n18004 18.301
R3526 vp_p.n19431 vp_p.n19430 18.301
R3527 vp_p.n20856 vp_p.n20855 18.301
R3528 vp_p.n22280 vp_p.n22279 18.301
R3529 vp_p.n23703 vp_p.n23702 18.301
R3530 vp_p.n25125 vp_p.n25124 18.301
R3531 vp_p.n26550 vp_p.n26549 18.301
R3532 vp_p.n12361 vp_p.n12360 18.301
R3533 vp_p.n10923 vp_p.n10922 18.301
R3534 vp_p.n9486 vp_p.n9485 18.301
R3535 vp_p.n740 vp_p.n739 18.301
R3536 vp_p.n2166 vp_p.n2165 18.301
R3537 vp_p.n3591 vp_p.n3590 18.301
R3538 vp_p.n5015 vp_p.n5014 18.301
R3539 vp_p.n6438 vp_p.n6437 18.301
R3540 vp_p.n7860 vp_p.n7859 18.301
R3541 vp_p.n15164 vp_p.n15163 18.301
R3542 vp_p.n16592 vp_p.n16591 18.301
R3543 vp_p.n18019 vp_p.n18018 18.301
R3544 vp_p.n19445 vp_p.n19444 18.301
R3545 vp_p.n20870 vp_p.n20869 18.301
R3546 vp_p.n22294 vp_p.n22293 18.301
R3547 vp_p.n23717 vp_p.n23716 18.301
R3548 vp_p.n25139 vp_p.n25138 18.301
R3549 vp_p.n26564 vp_p.n26563 18.301
R3550 vp_p.n12375 vp_p.n12374 18.301
R3551 vp_p.n10937 vp_p.n10936 18.301
R3552 vp_p.n9500 vp_p.n9499 18.301
R3553 vp_p.n754 vp_p.n753 18.301
R3554 vp_p.n2180 vp_p.n2179 18.301
R3555 vp_p.n3605 vp_p.n3604 18.301
R3556 vp_p.n5029 vp_p.n5028 18.301
R3557 vp_p.n6452 vp_p.n6451 18.301
R3558 vp_p.n7874 vp_p.n7873 18.301
R3559 vp_p.n15178 vp_p.n15177 18.301
R3560 vp_p.n16606 vp_p.n16605 18.301
R3561 vp_p.n18033 vp_p.n18032 18.301
R3562 vp_p.n19459 vp_p.n19458 18.301
R3563 vp_p.n20884 vp_p.n20883 18.301
R3564 vp_p.n22308 vp_p.n22307 18.301
R3565 vp_p.n23731 vp_p.n23730 18.301
R3566 vp_p.n25153 vp_p.n25152 18.301
R3567 vp_p.n26578 vp_p.n26577 18.301
R3568 vp_p.n12389 vp_p.n12388 18.301
R3569 vp_p.n10951 vp_p.n10950 18.301
R3570 vp_p.n9514 vp_p.n9513 18.301
R3571 vp_p.n768 vp_p.n767 18.301
R3572 vp_p.n2194 vp_p.n2193 18.301
R3573 vp_p.n3619 vp_p.n3618 18.301
R3574 vp_p.n5043 vp_p.n5042 18.301
R3575 vp_p.n6466 vp_p.n6465 18.301
R3576 vp_p.n7888 vp_p.n7887 18.301
R3577 vp_p.n15192 vp_p.n15191 18.301
R3578 vp_p.n16620 vp_p.n16619 18.301
R3579 vp_p.n18047 vp_p.n18046 18.301
R3580 vp_p.n19473 vp_p.n19472 18.301
R3581 vp_p.n20898 vp_p.n20897 18.301
R3582 vp_p.n22322 vp_p.n22321 18.301
R3583 vp_p.n23745 vp_p.n23744 18.301
R3584 vp_p.n25167 vp_p.n25166 18.301
R3585 vp_p.n26592 vp_p.n26591 18.301
R3586 vp_p.n12403 vp_p.n12402 18.301
R3587 vp_p.n10965 vp_p.n10964 18.301
R3588 vp_p.n9528 vp_p.n9527 18.301
R3589 vp_p.n782 vp_p.n781 18.301
R3590 vp_p.n2208 vp_p.n2207 18.301
R3591 vp_p.n3633 vp_p.n3632 18.301
R3592 vp_p.n5057 vp_p.n5056 18.301
R3593 vp_p.n6480 vp_p.n6479 18.301
R3594 vp_p.n7902 vp_p.n7901 18.301
R3595 vp_p.n15206 vp_p.n15205 18.301
R3596 vp_p.n16634 vp_p.n16633 18.301
R3597 vp_p.n18061 vp_p.n18060 18.301
R3598 vp_p.n19487 vp_p.n19486 18.301
R3599 vp_p.n20912 vp_p.n20911 18.301
R3600 vp_p.n22336 vp_p.n22335 18.301
R3601 vp_p.n23759 vp_p.n23758 18.301
R3602 vp_p.n25181 vp_p.n25180 18.301
R3603 vp_p.n26606 vp_p.n26605 18.301
R3604 vp_p.n12417 vp_p.n12416 18.301
R3605 vp_p.n10979 vp_p.n10978 18.301
R3606 vp_p.n9542 vp_p.n9541 18.301
R3607 vp_p.n796 vp_p.n795 18.301
R3608 vp_p.n2222 vp_p.n2221 18.301
R3609 vp_p.n3647 vp_p.n3646 18.301
R3610 vp_p.n5071 vp_p.n5070 18.301
R3611 vp_p.n6494 vp_p.n6493 18.301
R3612 vp_p.n7916 vp_p.n7915 18.301
R3613 vp_p.n15220 vp_p.n15219 18.301
R3614 vp_p.n16648 vp_p.n16647 18.301
R3615 vp_p.n18075 vp_p.n18074 18.301
R3616 vp_p.n19501 vp_p.n19500 18.301
R3617 vp_p.n20926 vp_p.n20925 18.301
R3618 vp_p.n22350 vp_p.n22349 18.301
R3619 vp_p.n23773 vp_p.n23772 18.301
R3620 vp_p.n25195 vp_p.n25194 18.301
R3621 vp_p.n26620 vp_p.n26619 18.301
R3622 vp_p.n12431 vp_p.n12430 18.301
R3623 vp_p.n10993 vp_p.n10992 18.301
R3624 vp_p.n9556 vp_p.n9555 18.301
R3625 vp_p.n810 vp_p.n809 18.301
R3626 vp_p.n2236 vp_p.n2235 18.301
R3627 vp_p.n3661 vp_p.n3660 18.301
R3628 vp_p.n5085 vp_p.n5084 18.301
R3629 vp_p.n6508 vp_p.n6507 18.301
R3630 vp_p.n7930 vp_p.n7929 18.301
R3631 vp_p.n15234 vp_p.n15233 18.301
R3632 vp_p.n16662 vp_p.n16661 18.301
R3633 vp_p.n18089 vp_p.n18088 18.301
R3634 vp_p.n19515 vp_p.n19514 18.301
R3635 vp_p.n20940 vp_p.n20939 18.301
R3636 vp_p.n22364 vp_p.n22363 18.301
R3637 vp_p.n23787 vp_p.n23786 18.301
R3638 vp_p.n25209 vp_p.n25208 18.301
R3639 vp_p.n26634 vp_p.n26633 18.301
R3640 vp_p.n12445 vp_p.n12444 18.301
R3641 vp_p.n11007 vp_p.n11006 18.301
R3642 vp_p.n9570 vp_p.n9569 18.301
R3643 vp_p.n824 vp_p.n823 18.301
R3644 vp_p.n2250 vp_p.n2249 18.301
R3645 vp_p.n3675 vp_p.n3674 18.301
R3646 vp_p.n5099 vp_p.n5098 18.301
R3647 vp_p.n6522 vp_p.n6521 18.301
R3648 vp_p.n7944 vp_p.n7943 18.301
R3649 vp_p.n15248 vp_p.n15247 18.301
R3650 vp_p.n16676 vp_p.n16675 18.301
R3651 vp_p.n18103 vp_p.n18102 18.301
R3652 vp_p.n19529 vp_p.n19528 18.301
R3653 vp_p.n20954 vp_p.n20953 18.301
R3654 vp_p.n22378 vp_p.n22377 18.301
R3655 vp_p.n23801 vp_p.n23800 18.301
R3656 vp_p.n25223 vp_p.n25222 18.301
R3657 vp_p.n26648 vp_p.n26647 18.301
R3658 vp_p.n12459 vp_p.n12458 18.301
R3659 vp_p.n11021 vp_p.n11020 18.301
R3660 vp_p.n9584 vp_p.n9583 18.301
R3661 vp_p.n838 vp_p.n837 18.301
R3662 vp_p.n2264 vp_p.n2263 18.301
R3663 vp_p.n3689 vp_p.n3688 18.301
R3664 vp_p.n5113 vp_p.n5112 18.301
R3665 vp_p.n6536 vp_p.n6535 18.301
R3666 vp_p.n7958 vp_p.n7957 18.301
R3667 vp_p.n15262 vp_p.n15261 18.301
R3668 vp_p.n16690 vp_p.n16689 18.301
R3669 vp_p.n18117 vp_p.n18116 18.301
R3670 vp_p.n19543 vp_p.n19542 18.301
R3671 vp_p.n20968 vp_p.n20967 18.301
R3672 vp_p.n22392 vp_p.n22391 18.301
R3673 vp_p.n23815 vp_p.n23814 18.301
R3674 vp_p.n25237 vp_p.n25236 18.301
R3675 vp_p.n26662 vp_p.n26661 18.301
R3676 vp_p.n12473 vp_p.n12472 18.301
R3677 vp_p.n11035 vp_p.n11034 18.301
R3678 vp_p.n9598 vp_p.n9597 18.301
R3679 vp_p.n852 vp_p.n851 18.301
R3680 vp_p.n2278 vp_p.n2277 18.301
R3681 vp_p.n3703 vp_p.n3702 18.301
R3682 vp_p.n5127 vp_p.n5126 18.301
R3683 vp_p.n6550 vp_p.n6549 18.301
R3684 vp_p.n7972 vp_p.n7971 18.301
R3685 vp_p.n15276 vp_p.n15275 18.301
R3686 vp_p.n16704 vp_p.n16703 18.301
R3687 vp_p.n18131 vp_p.n18130 18.301
R3688 vp_p.n19557 vp_p.n19556 18.301
R3689 vp_p.n20982 vp_p.n20981 18.301
R3690 vp_p.n22406 vp_p.n22405 18.301
R3691 vp_p.n23829 vp_p.n23828 18.301
R3692 vp_p.n25251 vp_p.n25250 18.301
R3693 vp_p.n26676 vp_p.n26675 18.301
R3694 vp_p.n12487 vp_p.n12486 18.301
R3695 vp_p.n11049 vp_p.n11048 18.301
R3696 vp_p.n9612 vp_p.n9611 18.301
R3697 vp_p.n866 vp_p.n865 18.301
R3698 vp_p.n2292 vp_p.n2291 18.301
R3699 vp_p.n3717 vp_p.n3716 18.301
R3700 vp_p.n5141 vp_p.n5140 18.301
R3701 vp_p.n6564 vp_p.n6563 18.301
R3702 vp_p.n7986 vp_p.n7985 18.301
R3703 vp_p.n15290 vp_p.n15289 18.301
R3704 vp_p.n16718 vp_p.n16717 18.301
R3705 vp_p.n18145 vp_p.n18144 18.301
R3706 vp_p.n19571 vp_p.n19570 18.301
R3707 vp_p.n20996 vp_p.n20995 18.301
R3708 vp_p.n22420 vp_p.n22419 18.301
R3709 vp_p.n23843 vp_p.n23842 18.301
R3710 vp_p.n25265 vp_p.n25264 18.301
R3711 vp_p.n26690 vp_p.n26689 18.301
R3712 vp_p.n12501 vp_p.n12500 18.301
R3713 vp_p.n11063 vp_p.n11062 18.301
R3714 vp_p.n9626 vp_p.n9625 18.301
R3715 vp_p.n880 vp_p.n879 18.301
R3716 vp_p.n2306 vp_p.n2305 18.301
R3717 vp_p.n3731 vp_p.n3730 18.301
R3718 vp_p.n5155 vp_p.n5154 18.301
R3719 vp_p.n6578 vp_p.n6577 18.301
R3720 vp_p.n8000 vp_p.n7999 18.301
R3721 vp_p.n15304 vp_p.n15303 18.301
R3722 vp_p.n16732 vp_p.n16731 18.301
R3723 vp_p.n18159 vp_p.n18158 18.301
R3724 vp_p.n19585 vp_p.n19584 18.301
R3725 vp_p.n21010 vp_p.n21009 18.301
R3726 vp_p.n22434 vp_p.n22433 18.301
R3727 vp_p.n23857 vp_p.n23856 18.301
R3728 vp_p.n25279 vp_p.n25278 18.301
R3729 vp_p.n26704 vp_p.n26703 18.301
R3730 vp_p.n12515 vp_p.n12514 18.301
R3731 vp_p.n11077 vp_p.n11076 18.301
R3732 vp_p.n9640 vp_p.n9639 18.301
R3733 vp_p.n894 vp_p.n893 18.301
R3734 vp_p.n2320 vp_p.n2319 18.301
R3735 vp_p.n3745 vp_p.n3744 18.301
R3736 vp_p.n5169 vp_p.n5168 18.301
R3737 vp_p.n6592 vp_p.n6591 18.301
R3738 vp_p.n8014 vp_p.n8013 18.301
R3739 vp_p.n15318 vp_p.n15317 18.301
R3740 vp_p.n16746 vp_p.n16745 18.301
R3741 vp_p.n18173 vp_p.n18172 18.301
R3742 vp_p.n19599 vp_p.n19598 18.301
R3743 vp_p.n21024 vp_p.n21023 18.301
R3744 vp_p.n22448 vp_p.n22447 18.301
R3745 vp_p.n23871 vp_p.n23870 18.301
R3746 vp_p.n25293 vp_p.n25292 18.301
R3747 vp_p.n26718 vp_p.n26717 18.301
R3748 vp_p.n12529 vp_p.n12528 18.301
R3749 vp_p.n11091 vp_p.n11090 18.301
R3750 vp_p.n9654 vp_p.n9653 18.301
R3751 vp_p.n908 vp_p.n907 18.301
R3752 vp_p.n2334 vp_p.n2333 18.301
R3753 vp_p.n3759 vp_p.n3758 18.301
R3754 vp_p.n5183 vp_p.n5182 18.301
R3755 vp_p.n6606 vp_p.n6605 18.301
R3756 vp_p.n8028 vp_p.n8027 18.301
R3757 vp_p.n15332 vp_p.n15331 18.301
R3758 vp_p.n16760 vp_p.n16759 18.301
R3759 vp_p.n18187 vp_p.n18186 18.301
R3760 vp_p.n19613 vp_p.n19612 18.301
R3761 vp_p.n21038 vp_p.n21037 18.301
R3762 vp_p.n22462 vp_p.n22461 18.301
R3763 vp_p.n23885 vp_p.n23884 18.301
R3764 vp_p.n25307 vp_p.n25306 18.301
R3765 vp_p.n26732 vp_p.n26731 18.301
R3766 vp_p.n12543 vp_p.n12542 18.301
R3767 vp_p.n11105 vp_p.n11104 18.301
R3768 vp_p.n9668 vp_p.n9667 18.301
R3769 vp_p.n922 vp_p.n921 18.301
R3770 vp_p.n2348 vp_p.n2347 18.301
R3771 vp_p.n3773 vp_p.n3772 18.301
R3772 vp_p.n5197 vp_p.n5196 18.301
R3773 vp_p.n6620 vp_p.n6619 18.301
R3774 vp_p.n8042 vp_p.n8041 18.301
R3775 vp_p.n15346 vp_p.n15345 18.301
R3776 vp_p.n16774 vp_p.n16773 18.301
R3777 vp_p.n18201 vp_p.n18200 18.301
R3778 vp_p.n19627 vp_p.n19626 18.301
R3779 vp_p.n21052 vp_p.n21051 18.301
R3780 vp_p.n22476 vp_p.n22475 18.301
R3781 vp_p.n23899 vp_p.n23898 18.301
R3782 vp_p.n25321 vp_p.n25320 18.301
R3783 vp_p.n26746 vp_p.n26745 18.301
R3784 vp_p.n12557 vp_p.n12556 18.301
R3785 vp_p.n11119 vp_p.n11118 18.301
R3786 vp_p.n9682 vp_p.n9681 18.301
R3787 vp_p.n936 vp_p.n935 18.301
R3788 vp_p.n2362 vp_p.n2361 18.301
R3789 vp_p.n3787 vp_p.n3786 18.301
R3790 vp_p.n5211 vp_p.n5210 18.301
R3791 vp_p.n6634 vp_p.n6633 18.301
R3792 vp_p.n8056 vp_p.n8055 18.301
R3793 vp_p.n15360 vp_p.n15359 18.301
R3794 vp_p.n16788 vp_p.n16787 18.301
R3795 vp_p.n18215 vp_p.n18214 18.301
R3796 vp_p.n19641 vp_p.n19640 18.301
R3797 vp_p.n21066 vp_p.n21065 18.301
R3798 vp_p.n22490 vp_p.n22489 18.301
R3799 vp_p.n23913 vp_p.n23912 18.301
R3800 vp_p.n25335 vp_p.n25334 18.301
R3801 vp_p.n26760 vp_p.n26759 18.301
R3802 vp_p.n12571 vp_p.n12570 18.301
R3803 vp_p.n11133 vp_p.n11132 18.301
R3804 vp_p.n9696 vp_p.n9695 18.301
R3805 vp_p.n950 vp_p.n949 18.301
R3806 vp_p.n2376 vp_p.n2375 18.301
R3807 vp_p.n3801 vp_p.n3800 18.301
R3808 vp_p.n5225 vp_p.n5224 18.301
R3809 vp_p.n6648 vp_p.n6647 18.301
R3810 vp_p.n8070 vp_p.n8069 18.301
R3811 vp_p.n15374 vp_p.n15373 18.301
R3812 vp_p.n16802 vp_p.n16801 18.301
R3813 vp_p.n18229 vp_p.n18228 18.301
R3814 vp_p.n19655 vp_p.n19654 18.301
R3815 vp_p.n21080 vp_p.n21079 18.301
R3816 vp_p.n22504 vp_p.n22503 18.301
R3817 vp_p.n23927 vp_p.n23926 18.301
R3818 vp_p.n25349 vp_p.n25348 18.301
R3819 vp_p.n26774 vp_p.n26773 18.301
R3820 vp_p.n12585 vp_p.n12584 18.301
R3821 vp_p.n11147 vp_p.n11146 18.301
R3822 vp_p.n9710 vp_p.n9709 18.301
R3823 vp_p.n964 vp_p.n963 18.301
R3824 vp_p.n2390 vp_p.n2389 18.301
R3825 vp_p.n3815 vp_p.n3814 18.301
R3826 vp_p.n5239 vp_p.n5238 18.301
R3827 vp_p.n6662 vp_p.n6661 18.301
R3828 vp_p.n8084 vp_p.n8083 18.301
R3829 vp_p.n15388 vp_p.n15387 18.301
R3830 vp_p.n16816 vp_p.n16815 18.301
R3831 vp_p.n18243 vp_p.n18242 18.301
R3832 vp_p.n19669 vp_p.n19668 18.301
R3833 vp_p.n21094 vp_p.n21093 18.301
R3834 vp_p.n22518 vp_p.n22517 18.301
R3835 vp_p.n23941 vp_p.n23940 18.301
R3836 vp_p.n25363 vp_p.n25362 18.301
R3837 vp_p.n26788 vp_p.n26787 18.301
R3838 vp_p.n12599 vp_p.n12598 18.301
R3839 vp_p.n11161 vp_p.n11160 18.301
R3840 vp_p.n9724 vp_p.n9723 18.301
R3841 vp_p.n978 vp_p.n977 18.301
R3842 vp_p.n2404 vp_p.n2403 18.301
R3843 vp_p.n3829 vp_p.n3828 18.301
R3844 vp_p.n5253 vp_p.n5252 18.301
R3845 vp_p.n6676 vp_p.n6675 18.301
R3846 vp_p.n8098 vp_p.n8097 18.301
R3847 vp_p.n15402 vp_p.n15401 18.301
R3848 vp_p.n16830 vp_p.n16829 18.301
R3849 vp_p.n18257 vp_p.n18256 18.301
R3850 vp_p.n19683 vp_p.n19682 18.301
R3851 vp_p.n21108 vp_p.n21107 18.301
R3852 vp_p.n22532 vp_p.n22531 18.301
R3853 vp_p.n23955 vp_p.n23954 18.301
R3854 vp_p.n25377 vp_p.n25376 18.301
R3855 vp_p.n26802 vp_p.n26801 18.301
R3856 vp_p.n12613 vp_p.n12612 18.301
R3857 vp_p.n11175 vp_p.n11174 18.301
R3858 vp_p.n9738 vp_p.n9737 18.301
R3859 vp_p.n992 vp_p.n991 18.301
R3860 vp_p.n2418 vp_p.n2417 18.301
R3861 vp_p.n3843 vp_p.n3842 18.301
R3862 vp_p.n5267 vp_p.n5266 18.301
R3863 vp_p.n6690 vp_p.n6689 18.301
R3864 vp_p.n8112 vp_p.n8111 18.301
R3865 vp_p.n15416 vp_p.n15415 18.301
R3866 vp_p.n16844 vp_p.n16843 18.301
R3867 vp_p.n18271 vp_p.n18270 18.301
R3868 vp_p.n19697 vp_p.n19696 18.301
R3869 vp_p.n21122 vp_p.n21121 18.301
R3870 vp_p.n22546 vp_p.n22545 18.301
R3871 vp_p.n23969 vp_p.n23968 18.301
R3872 vp_p.n25391 vp_p.n25390 18.301
R3873 vp_p.n26816 vp_p.n26815 18.301
R3874 vp_p.n12627 vp_p.n12626 18.301
R3875 vp_p.n11189 vp_p.n11188 18.301
R3876 vp_p.n9752 vp_p.n9751 18.301
R3877 vp_p.n1006 vp_p.n1005 18.301
R3878 vp_p.n2432 vp_p.n2431 18.301
R3879 vp_p.n3857 vp_p.n3856 18.301
R3880 vp_p.n5281 vp_p.n5280 18.301
R3881 vp_p.n6704 vp_p.n6703 18.301
R3882 vp_p.n8126 vp_p.n8125 18.301
R3883 vp_p.n15430 vp_p.n15429 18.301
R3884 vp_p.n16858 vp_p.n16857 18.301
R3885 vp_p.n18285 vp_p.n18284 18.301
R3886 vp_p.n19711 vp_p.n19710 18.301
R3887 vp_p.n21136 vp_p.n21135 18.301
R3888 vp_p.n22560 vp_p.n22559 18.301
R3889 vp_p.n23983 vp_p.n23982 18.301
R3890 vp_p.n25405 vp_p.n25404 18.301
R3891 vp_p.n26830 vp_p.n26829 18.301
R3892 vp_p.n12641 vp_p.n12640 18.301
R3893 vp_p.n11203 vp_p.n11202 18.301
R3894 vp_p.n9766 vp_p.n9765 18.301
R3895 vp_p.n1020 vp_p.n1019 18.301
R3896 vp_p.n2446 vp_p.n2445 18.301
R3897 vp_p.n3871 vp_p.n3870 18.301
R3898 vp_p.n5295 vp_p.n5294 18.301
R3899 vp_p.n6718 vp_p.n6717 18.301
R3900 vp_p.n8140 vp_p.n8139 18.301
R3901 vp_p.n15444 vp_p.n15443 18.301
R3902 vp_p.n16872 vp_p.n16871 18.301
R3903 vp_p.n18299 vp_p.n18298 18.301
R3904 vp_p.n19725 vp_p.n19724 18.301
R3905 vp_p.n21150 vp_p.n21149 18.301
R3906 vp_p.n22574 vp_p.n22573 18.301
R3907 vp_p.n23997 vp_p.n23996 18.301
R3908 vp_p.n25419 vp_p.n25418 18.301
R3909 vp_p.n26844 vp_p.n26843 18.301
R3910 vp_p.n12655 vp_p.n12654 18.301
R3911 vp_p.n11217 vp_p.n11216 18.301
R3912 vp_p.n9780 vp_p.n9779 18.301
R3913 vp_p.n1034 vp_p.n1033 18.301
R3914 vp_p.n2460 vp_p.n2459 18.301
R3915 vp_p.n3885 vp_p.n3884 18.301
R3916 vp_p.n5309 vp_p.n5308 18.301
R3917 vp_p.n6732 vp_p.n6731 18.301
R3918 vp_p.n8154 vp_p.n8153 18.301
R3919 vp_p.n15458 vp_p.n15457 18.301
R3920 vp_p.n16886 vp_p.n16885 18.301
R3921 vp_p.n18313 vp_p.n18312 18.301
R3922 vp_p.n19739 vp_p.n19738 18.301
R3923 vp_p.n21164 vp_p.n21163 18.301
R3924 vp_p.n22588 vp_p.n22587 18.301
R3925 vp_p.n24011 vp_p.n24010 18.301
R3926 vp_p.n25433 vp_p.n25432 18.301
R3927 vp_p.n26858 vp_p.n26857 18.301
R3928 vp_p.n12669 vp_p.n12668 18.301
R3929 vp_p.n11231 vp_p.n11230 18.301
R3930 vp_p.n9794 vp_p.n9793 18.301
R3931 vp_p.n1048 vp_p.n1047 18.301
R3932 vp_p.n2474 vp_p.n2473 18.301
R3933 vp_p.n3899 vp_p.n3898 18.301
R3934 vp_p.n5323 vp_p.n5322 18.301
R3935 vp_p.n6746 vp_p.n6745 18.301
R3936 vp_p.n8168 vp_p.n8167 18.301
R3937 vp_p.n15472 vp_p.n15471 18.301
R3938 vp_p.n16900 vp_p.n16899 18.301
R3939 vp_p.n18327 vp_p.n18326 18.301
R3940 vp_p.n19753 vp_p.n19752 18.301
R3941 vp_p.n21178 vp_p.n21177 18.301
R3942 vp_p.n22602 vp_p.n22601 18.301
R3943 vp_p.n24025 vp_p.n24024 18.301
R3944 vp_p.n25447 vp_p.n25446 18.301
R3945 vp_p.n26872 vp_p.n26871 18.301
R3946 vp_p.n12683 vp_p.n12682 18.301
R3947 vp_p.n11245 vp_p.n11244 18.301
R3948 vp_p.n9808 vp_p.n9807 18.301
R3949 vp_p.n1062 vp_p.n1061 18.301
R3950 vp_p.n2488 vp_p.n2487 18.301
R3951 vp_p.n3913 vp_p.n3912 18.301
R3952 vp_p.n5337 vp_p.n5336 18.301
R3953 vp_p.n6760 vp_p.n6759 18.301
R3954 vp_p.n8182 vp_p.n8181 18.301
R3955 vp_p.n15486 vp_p.n15485 18.301
R3956 vp_p.n16914 vp_p.n16913 18.301
R3957 vp_p.n18341 vp_p.n18340 18.301
R3958 vp_p.n19767 vp_p.n19766 18.301
R3959 vp_p.n21192 vp_p.n21191 18.301
R3960 vp_p.n22616 vp_p.n22615 18.301
R3961 vp_p.n24039 vp_p.n24038 18.301
R3962 vp_p.n25461 vp_p.n25460 18.301
R3963 vp_p.n26886 vp_p.n26885 18.301
R3964 vp_p.n12697 vp_p.n12696 18.301
R3965 vp_p.n11259 vp_p.n11258 18.301
R3966 vp_p.n9822 vp_p.n9821 18.301
R3967 vp_p.n1076 vp_p.n1075 18.301
R3968 vp_p.n2502 vp_p.n2501 18.301
R3969 vp_p.n3927 vp_p.n3926 18.301
R3970 vp_p.n5351 vp_p.n5350 18.301
R3971 vp_p.n6774 vp_p.n6773 18.301
R3972 vp_p.n8196 vp_p.n8195 18.301
R3973 vp_p.n15500 vp_p.n15499 18.301
R3974 vp_p.n16928 vp_p.n16927 18.301
R3975 vp_p.n18355 vp_p.n18354 18.301
R3976 vp_p.n19781 vp_p.n19780 18.301
R3977 vp_p.n21206 vp_p.n21205 18.301
R3978 vp_p.n22630 vp_p.n22629 18.301
R3979 vp_p.n24053 vp_p.n24052 18.301
R3980 vp_p.n25475 vp_p.n25474 18.301
R3981 vp_p.n26900 vp_p.n26899 18.301
R3982 vp_p.n12711 vp_p.n12710 18.301
R3983 vp_p.n11273 vp_p.n11272 18.301
R3984 vp_p.n9836 vp_p.n9835 18.301
R3985 vp_p.n1090 vp_p.n1089 18.301
R3986 vp_p.n2516 vp_p.n2515 18.301
R3987 vp_p.n3941 vp_p.n3940 18.301
R3988 vp_p.n5365 vp_p.n5364 18.301
R3989 vp_p.n6788 vp_p.n6787 18.301
R3990 vp_p.n8210 vp_p.n8209 18.301
R3991 vp_p.n15514 vp_p.n15513 18.301
R3992 vp_p.n16942 vp_p.n16941 18.301
R3993 vp_p.n18369 vp_p.n18368 18.301
R3994 vp_p.n19795 vp_p.n19794 18.301
R3995 vp_p.n21220 vp_p.n21219 18.301
R3996 vp_p.n22644 vp_p.n22643 18.301
R3997 vp_p.n24067 vp_p.n24066 18.301
R3998 vp_p.n25489 vp_p.n25488 18.301
R3999 vp_p.n26914 vp_p.n26913 18.301
R4000 vp_p.n12725 vp_p.n12724 18.301
R4001 vp_p.n11287 vp_p.n11286 18.301
R4002 vp_p.n9850 vp_p.n9849 18.301
R4003 vp_p.n1104 vp_p.n1103 18.301
R4004 vp_p.n2530 vp_p.n2529 18.301
R4005 vp_p.n3955 vp_p.n3954 18.301
R4006 vp_p.n5379 vp_p.n5378 18.301
R4007 vp_p.n6802 vp_p.n6801 18.301
R4008 vp_p.n8224 vp_p.n8223 18.301
R4009 vp_p.n15528 vp_p.n15527 18.301
R4010 vp_p.n16956 vp_p.n16955 18.301
R4011 vp_p.n18383 vp_p.n18382 18.301
R4012 vp_p.n19809 vp_p.n19808 18.301
R4013 vp_p.n21234 vp_p.n21233 18.301
R4014 vp_p.n22658 vp_p.n22657 18.301
R4015 vp_p.n24081 vp_p.n24080 18.301
R4016 vp_p.n25503 vp_p.n25502 18.301
R4017 vp_p.n26928 vp_p.n26927 18.301
R4018 vp_p.n12739 vp_p.n12738 18.301
R4019 vp_p.n11301 vp_p.n11300 18.301
R4020 vp_p.n9864 vp_p.n9863 18.301
R4021 vp_p.n1118 vp_p.n1117 18.301
R4022 vp_p.n2544 vp_p.n2543 18.301
R4023 vp_p.n3969 vp_p.n3968 18.301
R4024 vp_p.n5393 vp_p.n5392 18.301
R4025 vp_p.n6816 vp_p.n6815 18.301
R4026 vp_p.n8238 vp_p.n8237 18.301
R4027 vp_p.n15542 vp_p.n15541 18.301
R4028 vp_p.n16970 vp_p.n16969 18.301
R4029 vp_p.n18397 vp_p.n18396 18.301
R4030 vp_p.n19823 vp_p.n19822 18.301
R4031 vp_p.n21248 vp_p.n21247 18.301
R4032 vp_p.n22672 vp_p.n22671 18.301
R4033 vp_p.n24095 vp_p.n24094 18.301
R4034 vp_p.n25517 vp_p.n25516 18.301
R4035 vp_p.n26942 vp_p.n26941 18.301
R4036 vp_p.n12753 vp_p.n12752 18.301
R4037 vp_p.n11315 vp_p.n11314 18.301
R4038 vp_p.n9878 vp_p.n9877 18.301
R4039 vp_p.n1132 vp_p.n1131 18.301
R4040 vp_p.n2558 vp_p.n2557 18.301
R4041 vp_p.n3983 vp_p.n3982 18.301
R4042 vp_p.n5407 vp_p.n5406 18.301
R4043 vp_p.n6830 vp_p.n6829 18.301
R4044 vp_p.n8252 vp_p.n8251 18.301
R4045 vp_p.n15556 vp_p.n15555 18.301
R4046 vp_p.n16984 vp_p.n16983 18.301
R4047 vp_p.n18411 vp_p.n18410 18.301
R4048 vp_p.n19837 vp_p.n19836 18.301
R4049 vp_p.n21262 vp_p.n21261 18.301
R4050 vp_p.n22686 vp_p.n22685 18.301
R4051 vp_p.n24109 vp_p.n24108 18.301
R4052 vp_p.n25531 vp_p.n25530 18.301
R4053 vp_p.n26956 vp_p.n26955 18.301
R4054 vp_p.n12767 vp_p.n12766 18.301
R4055 vp_p.n11329 vp_p.n11328 18.301
R4056 vp_p.n9892 vp_p.n9891 18.301
R4057 vp_p.n1146 vp_p.n1145 18.301
R4058 vp_p.n2572 vp_p.n2571 18.301
R4059 vp_p.n3997 vp_p.n3996 18.301
R4060 vp_p.n5421 vp_p.n5420 18.301
R4061 vp_p.n6844 vp_p.n6843 18.301
R4062 vp_p.n8266 vp_p.n8265 18.301
R4063 vp_p.n15570 vp_p.n15569 18.301
R4064 vp_p.n16998 vp_p.n16997 18.301
R4065 vp_p.n18425 vp_p.n18424 18.301
R4066 vp_p.n19851 vp_p.n19850 18.301
R4067 vp_p.n21276 vp_p.n21275 18.301
R4068 vp_p.n22700 vp_p.n22699 18.301
R4069 vp_p.n24123 vp_p.n24122 18.301
R4070 vp_p.n25545 vp_p.n25544 18.301
R4071 vp_p.n26970 vp_p.n26969 18.301
R4072 vp_p.n12781 vp_p.n12780 18.301
R4073 vp_p.n11343 vp_p.n11342 18.301
R4074 vp_p.n9906 vp_p.n9905 18.301
R4075 vp_p.n1160 vp_p.n1159 18.301
R4076 vp_p.n2586 vp_p.n2585 18.301
R4077 vp_p.n4011 vp_p.n4010 18.301
R4078 vp_p.n5435 vp_p.n5434 18.301
R4079 vp_p.n6858 vp_p.n6857 18.301
R4080 vp_p.n8280 vp_p.n8279 18.301
R4081 vp_p.n15584 vp_p.n15583 18.301
R4082 vp_p.n17012 vp_p.n17011 18.301
R4083 vp_p.n18439 vp_p.n18438 18.301
R4084 vp_p.n19865 vp_p.n19864 18.301
R4085 vp_p.n21290 vp_p.n21289 18.301
R4086 vp_p.n22714 vp_p.n22713 18.301
R4087 vp_p.n24137 vp_p.n24136 18.301
R4088 vp_p.n25559 vp_p.n25558 18.301
R4089 vp_p.n26984 vp_p.n26983 18.301
R4090 vp_p.n12795 vp_p.n12794 18.301
R4091 vp_p.n11357 vp_p.n11356 18.301
R4092 vp_p.n9920 vp_p.n9919 18.301
R4093 vp_p.n1174 vp_p.n1173 18.301
R4094 vp_p.n2600 vp_p.n2599 18.301
R4095 vp_p.n4025 vp_p.n4024 18.301
R4096 vp_p.n5449 vp_p.n5448 18.301
R4097 vp_p.n6872 vp_p.n6871 18.301
R4098 vp_p.n8294 vp_p.n8293 18.301
R4099 vp_p.n15598 vp_p.n15597 18.301
R4100 vp_p.n17026 vp_p.n17025 18.301
R4101 vp_p.n18453 vp_p.n18452 18.301
R4102 vp_p.n19879 vp_p.n19878 18.301
R4103 vp_p.n21304 vp_p.n21303 18.301
R4104 vp_p.n22728 vp_p.n22727 18.301
R4105 vp_p.n24151 vp_p.n24150 18.301
R4106 vp_p.n25573 vp_p.n25572 18.301
R4107 vp_p.n26998 vp_p.n26997 18.301
R4108 vp_p.n12809 vp_p.n12808 18.301
R4109 vp_p.n11371 vp_p.n11370 18.301
R4110 vp_p.n9934 vp_p.n9933 18.301
R4111 vp_p.n1188 vp_p.n1187 18.301
R4112 vp_p.n2614 vp_p.n2613 18.301
R4113 vp_p.n4039 vp_p.n4038 18.301
R4114 vp_p.n5463 vp_p.n5462 18.301
R4115 vp_p.n6886 vp_p.n6885 18.301
R4116 vp_p.n8308 vp_p.n8307 18.301
R4117 vp_p.n15612 vp_p.n15611 18.301
R4118 vp_p.n17040 vp_p.n17039 18.301
R4119 vp_p.n18467 vp_p.n18466 18.301
R4120 vp_p.n19893 vp_p.n19892 18.301
R4121 vp_p.n21318 vp_p.n21317 18.301
R4122 vp_p.n22742 vp_p.n22741 18.301
R4123 vp_p.n24165 vp_p.n24164 18.301
R4124 vp_p.n25587 vp_p.n25586 18.301
R4125 vp_p.n27012 vp_p.n27011 18.301
R4126 vp_p.n12823 vp_p.n12822 18.301
R4127 vp_p.n11385 vp_p.n11384 18.301
R4128 vp_p.n9948 vp_p.n9947 18.301
R4129 vp_p.n1202 vp_p.n1201 18.301
R4130 vp_p.n2628 vp_p.n2627 18.301
R4131 vp_p.n4053 vp_p.n4052 18.301
R4132 vp_p.n5477 vp_p.n5476 18.301
R4133 vp_p.n6900 vp_p.n6899 18.301
R4134 vp_p.n8322 vp_p.n8321 18.301
R4135 vp_p.n15626 vp_p.n15625 18.301
R4136 vp_p.n17054 vp_p.n17053 18.301
R4137 vp_p.n18481 vp_p.n18480 18.301
R4138 vp_p.n19907 vp_p.n19906 18.301
R4139 vp_p.n21332 vp_p.n21331 18.301
R4140 vp_p.n22756 vp_p.n22755 18.301
R4141 vp_p.n24179 vp_p.n24178 18.301
R4142 vp_p.n25601 vp_p.n25600 18.301
R4143 vp_p.n27026 vp_p.n27025 18.301
R4144 vp_p.n12837 vp_p.n12836 18.301
R4145 vp_p.n11399 vp_p.n11398 18.301
R4146 vp_p.n9962 vp_p.n9961 18.301
R4147 vp_p.n1216 vp_p.n1215 18.301
R4148 vp_p.n2642 vp_p.n2641 18.301
R4149 vp_p.n4067 vp_p.n4066 18.301
R4150 vp_p.n5491 vp_p.n5490 18.301
R4151 vp_p.n6914 vp_p.n6913 18.301
R4152 vp_p.n8336 vp_p.n8335 18.301
R4153 vp_p.n15640 vp_p.n15639 18.301
R4154 vp_p.n17068 vp_p.n17067 18.301
R4155 vp_p.n18495 vp_p.n18494 18.301
R4156 vp_p.n19921 vp_p.n19920 18.301
R4157 vp_p.n21346 vp_p.n21345 18.301
R4158 vp_p.n22770 vp_p.n22769 18.301
R4159 vp_p.n24193 vp_p.n24192 18.301
R4160 vp_p.n25615 vp_p.n25614 18.301
R4161 vp_p.n27040 vp_p.n27039 18.301
R4162 vp_p.n12851 vp_p.n12850 18.301
R4163 vp_p.n11413 vp_p.n11412 18.301
R4164 vp_p.n9976 vp_p.n9975 18.301
R4165 vp_p.n1230 vp_p.n1229 18.301
R4166 vp_p.n2656 vp_p.n2655 18.301
R4167 vp_p.n4081 vp_p.n4080 18.301
R4168 vp_p.n5505 vp_p.n5504 18.301
R4169 vp_p.n6928 vp_p.n6927 18.301
R4170 vp_p.n8350 vp_p.n8349 18.301
R4171 vp_p.n15654 vp_p.n15653 18.301
R4172 vp_p.n17082 vp_p.n17081 18.301
R4173 vp_p.n18509 vp_p.n18508 18.301
R4174 vp_p.n19935 vp_p.n19934 18.301
R4175 vp_p.n21360 vp_p.n21359 18.301
R4176 vp_p.n22784 vp_p.n22783 18.301
R4177 vp_p.n24207 vp_p.n24206 18.301
R4178 vp_p.n25629 vp_p.n25628 18.301
R4179 vp_p.n27054 vp_p.n27053 18.301
R4180 vp_p.n12865 vp_p.n12864 18.301
R4181 vp_p.n11427 vp_p.n11426 18.301
R4182 vp_p.n9990 vp_p.n9989 18.301
R4183 vp_p.n1244 vp_p.n1243 18.301
R4184 vp_p.n2670 vp_p.n2669 18.301
R4185 vp_p.n4095 vp_p.n4094 18.301
R4186 vp_p.n5519 vp_p.n5518 18.301
R4187 vp_p.n6942 vp_p.n6941 18.301
R4188 vp_p.n8364 vp_p.n8363 18.301
R4189 vp_p.n15668 vp_p.n15667 18.301
R4190 vp_p.n17096 vp_p.n17095 18.301
R4191 vp_p.n18523 vp_p.n18522 18.301
R4192 vp_p.n19949 vp_p.n19948 18.301
R4193 vp_p.n21374 vp_p.n21373 18.301
R4194 vp_p.n22798 vp_p.n22797 18.301
R4195 vp_p.n24221 vp_p.n24220 18.301
R4196 vp_p.n25643 vp_p.n25642 18.301
R4197 vp_p.n27068 vp_p.n27067 18.301
R4198 vp_p.n12879 vp_p.n12878 18.301
R4199 vp_p.n11441 vp_p.n11440 18.301
R4200 vp_p.n10004 vp_p.n10003 18.301
R4201 vp_p.n1258 vp_p.n1257 18.301
R4202 vp_p.n2684 vp_p.n2683 18.301
R4203 vp_p.n4109 vp_p.n4108 18.301
R4204 vp_p.n5533 vp_p.n5532 18.301
R4205 vp_p.n6956 vp_p.n6955 18.301
R4206 vp_p.n8378 vp_p.n8377 18.301
R4207 vp_p.n15682 vp_p.n15681 18.301
R4208 vp_p.n17110 vp_p.n17109 18.301
R4209 vp_p.n18537 vp_p.n18536 18.301
R4210 vp_p.n19963 vp_p.n19962 18.301
R4211 vp_p.n21388 vp_p.n21387 18.301
R4212 vp_p.n22812 vp_p.n22811 18.301
R4213 vp_p.n24235 vp_p.n24234 18.301
R4214 vp_p.n25657 vp_p.n25656 18.301
R4215 vp_p.n27082 vp_p.n27081 18.301
R4216 vp_p.n12893 vp_p.n12892 18.301
R4217 vp_p.n11455 vp_p.n11454 18.301
R4218 vp_p.n10018 vp_p.n10017 18.301
R4219 vp_p.n1272 vp_p.n1271 18.301
R4220 vp_p.n2698 vp_p.n2697 18.301
R4221 vp_p.n4123 vp_p.n4122 18.301
R4222 vp_p.n5547 vp_p.n5546 18.301
R4223 vp_p.n6970 vp_p.n6969 18.301
R4224 vp_p.n8392 vp_p.n8391 18.301
R4225 vp_p.n15696 vp_p.n15695 18.301
R4226 vp_p.n17124 vp_p.n17123 18.301
R4227 vp_p.n18551 vp_p.n18550 18.301
R4228 vp_p.n19977 vp_p.n19976 18.301
R4229 vp_p.n21402 vp_p.n21401 18.301
R4230 vp_p.n22826 vp_p.n22825 18.301
R4231 vp_p.n24249 vp_p.n24248 18.301
R4232 vp_p.n25671 vp_p.n25670 18.301
R4233 vp_p.n27096 vp_p.n27095 18.301
R4234 vp_p.n12907 vp_p.n12906 18.301
R4235 vp_p.n11469 vp_p.n11468 18.301
R4236 vp_p.n10032 vp_p.n10031 18.301
R4237 vp_p.n1286 vp_p.n1285 18.301
R4238 vp_p.n2712 vp_p.n2711 18.301
R4239 vp_p.n4137 vp_p.n4136 18.301
R4240 vp_p.n5561 vp_p.n5560 18.301
R4241 vp_p.n6984 vp_p.n6983 18.301
R4242 vp_p.n8406 vp_p.n8405 18.301
R4243 vp_p.n15710 vp_p.n15709 18.301
R4244 vp_p.n17138 vp_p.n17137 18.301
R4245 vp_p.n18565 vp_p.n18564 18.301
R4246 vp_p.n19991 vp_p.n19990 18.301
R4247 vp_p.n21416 vp_p.n21415 18.301
R4248 vp_p.n22840 vp_p.n22839 18.301
R4249 vp_p.n24263 vp_p.n24262 18.301
R4250 vp_p.n25685 vp_p.n25684 18.301
R4251 vp_p.n27110 vp_p.n27109 18.301
R4252 vp_p.n12921 vp_p.n12920 18.301
R4253 vp_p.n11483 vp_p.n11482 18.301
R4254 vp_p.n10046 vp_p.n10045 18.301
R4255 vp_p.n1300 vp_p.n1299 18.301
R4256 vp_p.n2726 vp_p.n2725 18.301
R4257 vp_p.n4151 vp_p.n4150 18.301
R4258 vp_p.n5575 vp_p.n5574 18.301
R4259 vp_p.n6998 vp_p.n6997 18.301
R4260 vp_p.n8420 vp_p.n8419 18.301
R4261 vp_p.n15724 vp_p.n15723 18.301
R4262 vp_p.n17152 vp_p.n17151 18.301
R4263 vp_p.n18579 vp_p.n18578 18.301
R4264 vp_p.n20005 vp_p.n20004 18.301
R4265 vp_p.n21430 vp_p.n21429 18.301
R4266 vp_p.n22854 vp_p.n22853 18.301
R4267 vp_p.n24277 vp_p.n24276 18.301
R4268 vp_p.n25699 vp_p.n25698 18.301
R4269 vp_p.n27124 vp_p.n27123 18.301
R4270 vp_p.n12935 vp_p.n12934 18.301
R4271 vp_p.n11497 vp_p.n11496 18.301
R4272 vp_p.n10060 vp_p.n10059 18.301
R4273 vp_p.n1314 vp_p.n1313 18.301
R4274 vp_p.n2740 vp_p.n2739 18.301
R4275 vp_p.n4165 vp_p.n4164 18.301
R4276 vp_p.n5589 vp_p.n5588 18.301
R4277 vp_p.n7012 vp_p.n7011 18.301
R4278 vp_p.n8434 vp_p.n8433 18.301
R4279 vp_p.n15738 vp_p.n15737 18.301
R4280 vp_p.n17166 vp_p.n17165 18.301
R4281 vp_p.n18593 vp_p.n18592 18.301
R4282 vp_p.n20019 vp_p.n20018 18.301
R4283 vp_p.n21444 vp_p.n21443 18.301
R4284 vp_p.n22868 vp_p.n22867 18.301
R4285 vp_p.n24291 vp_p.n24290 18.301
R4286 vp_p.n25713 vp_p.n25712 18.301
R4287 vp_p.n27138 vp_p.n27137 18.301
R4288 vp_p.n12949 vp_p.n12948 18.301
R4289 vp_p.n11511 vp_p.n11510 18.301
R4290 vp_p.n10074 vp_p.n10073 18.301
R4291 vp_p.n1328 vp_p.n1327 18.301
R4292 vp_p.n2754 vp_p.n2753 18.301
R4293 vp_p.n4179 vp_p.n4178 18.301
R4294 vp_p.n5603 vp_p.n5602 18.301
R4295 vp_p.n7026 vp_p.n7025 18.301
R4296 vp_p.n8448 vp_p.n8447 18.301
R4297 vp_p.n15752 vp_p.n15751 18.301
R4298 vp_p.n17180 vp_p.n17179 18.301
R4299 vp_p.n18607 vp_p.n18606 18.301
R4300 vp_p.n20033 vp_p.n20032 18.301
R4301 vp_p.n21458 vp_p.n21457 18.301
R4302 vp_p.n22882 vp_p.n22881 18.301
R4303 vp_p.n24305 vp_p.n24304 18.301
R4304 vp_p.n25727 vp_p.n25726 18.301
R4305 vp_p.n27152 vp_p.n27151 18.301
R4306 vp_p.n12963 vp_p.n12962 18.301
R4307 vp_p.n11525 vp_p.n11524 18.301
R4308 vp_p.n10088 vp_p.n10087 18.301
R4309 vp_p.n1342 vp_p.n1341 18.301
R4310 vp_p.n2768 vp_p.n2767 18.301
R4311 vp_p.n4193 vp_p.n4192 18.301
R4312 vp_p.n5617 vp_p.n5616 18.301
R4313 vp_p.n7040 vp_p.n7039 18.301
R4314 vp_p.n8462 vp_p.n8461 18.301
R4315 vp_p.n15766 vp_p.n15765 18.301
R4316 vp_p.n17194 vp_p.n17193 18.301
R4317 vp_p.n18621 vp_p.n18620 18.301
R4318 vp_p.n20047 vp_p.n20046 18.301
R4319 vp_p.n21472 vp_p.n21471 18.301
R4320 vp_p.n22896 vp_p.n22895 18.301
R4321 vp_p.n24319 vp_p.n24318 18.301
R4322 vp_p.n25741 vp_p.n25740 18.301
R4323 vp_p.n27166 vp_p.n27165 18.301
R4324 vp_p.n12977 vp_p.n12976 18.301
R4325 vp_p.n11539 vp_p.n11538 18.301
R4326 vp_p.n10102 vp_p.n10101 18.301
R4327 vp_p.n1356 vp_p.n1355 18.301
R4328 vp_p.n2782 vp_p.n2781 18.301
R4329 vp_p.n4207 vp_p.n4206 18.301
R4330 vp_p.n5631 vp_p.n5630 18.301
R4331 vp_p.n7054 vp_p.n7053 18.301
R4332 vp_p.n8476 vp_p.n8475 18.301
R4333 vp_p.n15780 vp_p.n15779 18.301
R4334 vp_p.n17208 vp_p.n17207 18.301
R4335 vp_p.n18635 vp_p.n18634 18.301
R4336 vp_p.n20061 vp_p.n20060 18.301
R4337 vp_p.n21486 vp_p.n21485 18.301
R4338 vp_p.n22910 vp_p.n22909 18.301
R4339 vp_p.n24333 vp_p.n24332 18.301
R4340 vp_p.n25755 vp_p.n25754 18.301
R4341 vp_p.n27180 vp_p.n27179 18.301
R4342 vp_p.n12991 vp_p.n12990 18.301
R4343 vp_p.n11553 vp_p.n11552 18.301
R4344 vp_p.n10116 vp_p.n10115 18.301
R4345 vp_p.n1370 vp_p.n1369 18.301
R4346 vp_p.n2796 vp_p.n2795 18.301
R4347 vp_p.n4221 vp_p.n4220 18.301
R4348 vp_p.n5645 vp_p.n5644 18.301
R4349 vp_p.n7068 vp_p.n7067 18.301
R4350 vp_p.n8490 vp_p.n8489 18.301
R4351 vp_p.n15794 vp_p.n15793 18.301
R4352 vp_p.n17222 vp_p.n17221 18.301
R4353 vp_p.n18649 vp_p.n18648 18.301
R4354 vp_p.n20075 vp_p.n20074 18.301
R4355 vp_p.n21500 vp_p.n21499 18.301
R4356 vp_p.n22924 vp_p.n22923 18.301
R4357 vp_p.n24347 vp_p.n24346 18.301
R4358 vp_p.n25769 vp_p.n25768 18.301
R4359 vp_p.n27194 vp_p.n27193 18.301
R4360 vp_p.n13005 vp_p.n13004 18.301
R4361 vp_p.n11567 vp_p.n11566 18.301
R4362 vp_p.n10130 vp_p.n10129 18.301
R4363 vp_p.n1384 vp_p.n1383 18.301
R4364 vp_p.n2810 vp_p.n2809 18.301
R4365 vp_p.n4235 vp_p.n4234 18.301
R4366 vp_p.n5659 vp_p.n5658 18.301
R4367 vp_p.n7082 vp_p.n7081 18.301
R4368 vp_p.n8504 vp_p.n8503 18.301
R4369 vp_p.n15808 vp_p.n15807 18.301
R4370 vp_p.n17236 vp_p.n17235 18.301
R4371 vp_p.n18663 vp_p.n18662 18.301
R4372 vp_p.n20089 vp_p.n20088 18.301
R4373 vp_p.n21514 vp_p.n21513 18.301
R4374 vp_p.n22938 vp_p.n22937 18.301
R4375 vp_p.n24361 vp_p.n24360 18.301
R4376 vp_p.n25783 vp_p.n25782 18.301
R4377 vp_p.n27208 vp_p.n27207 18.301
R4378 vp_p.n11581 vp_p.n11580 18.301
R4379 vp_p.n10144 vp_p.n10143 18.301
R4380 vp_p.n1398 vp_p.n1397 18.301
R4381 vp_p.n2824 vp_p.n2823 18.301
R4382 vp_p.n4249 vp_p.n4248 18.301
R4383 vp_p.n5673 vp_p.n5672 18.301
R4384 vp_p.n7096 vp_p.n7095 18.301
R4385 vp_p.n8518 vp_p.n8517 18.301
R4386 vp_p.n17250 vp_p.n17249 18.301
R4387 vp_p.n18677 vp_p.n18676 18.301
R4388 vp_p.n20103 vp_p.n20102 18.301
R4389 vp_p.n21528 vp_p.n21527 18.301
R4390 vp_p.n22952 vp_p.n22951 18.301
R4391 vp_p.n24375 vp_p.n24374 18.301
R4392 vp_p.n25797 vp_p.n25796 18.301
R4393 vp_p.n27222 vp_p.n27221 18.301
R4394 vp_p.n10158 vp_p.n10157 18.301
R4395 vp_p.n1412 vp_p.n1411 18.301
R4396 vp_p.n2838 vp_p.n2837 18.301
R4397 vp_p.n4263 vp_p.n4262 18.301
R4398 vp_p.n5687 vp_p.n5686 18.301
R4399 vp_p.n7110 vp_p.n7109 18.301
R4400 vp_p.n8532 vp_p.n8531 18.301
R4401 vp_p.n18691 vp_p.n18690 18.301
R4402 vp_p.n20117 vp_p.n20116 18.301
R4403 vp_p.n21542 vp_p.n21541 18.301
R4404 vp_p.n22966 vp_p.n22965 18.301
R4405 vp_p.n24389 vp_p.n24388 18.301
R4406 vp_p.n25811 vp_p.n25810 18.301
R4407 vp_p.n27236 vp_p.n27235 18.301
R4408 vp_p.n1426 vp_p.n1425 18.301
R4409 vp_p.n2852 vp_p.n2851 18.301
R4410 vp_p.n4277 vp_p.n4276 18.301
R4411 vp_p.n5701 vp_p.n5700 18.301
R4412 vp_p.n7124 vp_p.n7123 18.301
R4413 vp_p.n8546 vp_p.n8545 18.301
R4414 vp_p.n20131 vp_p.n20130 18.301
R4415 vp_p.n21556 vp_p.n21555 18.301
R4416 vp_p.n22980 vp_p.n22979 18.301
R4417 vp_p.n24403 vp_p.n24402 18.301
R4418 vp_p.n25825 vp_p.n25824 18.301
R4419 vp_p.n27250 vp_p.n27249 18.301
R4420 vp_p.n2866 vp_p.n2865 18.301
R4421 vp_p.n4291 vp_p.n4290 18.301
R4422 vp_p.n5715 vp_p.n5714 18.301
R4423 vp_p.n7138 vp_p.n7137 18.301
R4424 vp_p.n8560 vp_p.n8559 18.301
R4425 vp_p.n21570 vp_p.n21569 18.301
R4426 vp_p.n22994 vp_p.n22993 18.301
R4427 vp_p.n24417 vp_p.n24416 18.301
R4428 vp_p.n25839 vp_p.n25838 18.301
R4429 vp_p.n27264 vp_p.n27263 18.301
R4430 vp_p.n4305 vp_p.n4304 18.301
R4431 vp_p.n5729 vp_p.n5728 18.301
R4432 vp_p.n7152 vp_p.n7151 18.301
R4433 vp_p.n8574 vp_p.n8573 18.301
R4434 vp_p.n23008 vp_p.n23007 18.301
R4435 vp_p.n24431 vp_p.n24430 18.301
R4436 vp_p.n25853 vp_p.n25852 18.301
R4437 vp_p.n27278 vp_p.n27277 18.301
R4438 vp_p.n5743 vp_p.n5742 18.301
R4439 vp_p.n7166 vp_p.n7165 18.301
R4440 vp_p.n8588 vp_p.n8587 18.301
R4441 vp_p.n24445 vp_p.n24444 18.301
R4442 vp_p.n25867 vp_p.n25866 18.301
R4443 vp_p.n27292 vp_p.n27291 18.301
R4444 vp_p.n7180 vp_p.n7179 18.301
R4445 vp_p.n8602 vp_p.n8601 18.301
R4446 vp_p.n25881 vp_p.n25880 18.301
R4447 vp_p.n27306 vp_p.n27305 18.301
R4448 vp_p.n8616 vp_p.n8615 18.301
R4449 vp_p.n27320 vp_p.n27319 18.301
R4450 vp_p.n13005 vp_p.n13002 16.403
R4451 vp_p.n12991 vp_p.n12988 16.403
R4452 vp_p.n12977 vp_p.n12974 16.403
R4453 vp_p.n12963 vp_p.n12960 16.403
R4454 vp_p.n12949 vp_p.n12946 16.403
R4455 vp_p.n12935 vp_p.n12932 16.403
R4456 vp_p.n12921 vp_p.n12918 16.403
R4457 vp_p.n12907 vp_p.n12904 16.403
R4458 vp_p.n12893 vp_p.n12890 16.403
R4459 vp_p.n12879 vp_p.n12876 16.403
R4460 vp_p.n12865 vp_p.n12862 16.403
R4461 vp_p.n12851 vp_p.n12848 16.403
R4462 vp_p.n12837 vp_p.n12834 16.403
R4463 vp_p.n12823 vp_p.n12820 16.403
R4464 vp_p.n12809 vp_p.n12806 16.403
R4465 vp_p.n12795 vp_p.n12792 16.403
R4466 vp_p.n12781 vp_p.n12778 16.403
R4467 vp_p.n12767 vp_p.n12764 16.403
R4468 vp_p.n12753 vp_p.n12750 16.403
R4469 vp_p.n12739 vp_p.n12736 16.403
R4470 vp_p.n12725 vp_p.n12722 16.403
R4471 vp_p.n12711 vp_p.n12708 16.403
R4472 vp_p.n12697 vp_p.n12694 16.403
R4473 vp_p.n12683 vp_p.n12680 16.403
R4474 vp_p.n12669 vp_p.n12666 16.403
R4475 vp_p.n12655 vp_p.n12652 16.403
R4476 vp_p.n12641 vp_p.n12638 16.403
R4477 vp_p.n12627 vp_p.n12624 16.403
R4478 vp_p.n12613 vp_p.n12610 16.403
R4479 vp_p.n12599 vp_p.n12596 16.403
R4480 vp_p.n12585 vp_p.n12582 16.403
R4481 vp_p.n12571 vp_p.n12568 16.403
R4482 vp_p.n12557 vp_p.n12554 16.403
R4483 vp_p.n12543 vp_p.n12540 16.403
R4484 vp_p.n12529 vp_p.n12526 16.403
R4485 vp_p.n12515 vp_p.n12512 16.403
R4486 vp_p.n12501 vp_p.n12498 16.403
R4487 vp_p.n12487 vp_p.n12484 16.403
R4488 vp_p.n12473 vp_p.n12470 16.403
R4489 vp_p.n12459 vp_p.n12456 16.403
R4490 vp_p.n12445 vp_p.n12442 16.403
R4491 vp_p.n12431 vp_p.n12428 16.403
R4492 vp_p.n12417 vp_p.n12414 16.403
R4493 vp_p.n12403 vp_p.n12400 16.403
R4494 vp_p.n12389 vp_p.n12386 16.403
R4495 vp_p.n12375 vp_p.n12372 16.403
R4496 vp_p.n12361 vp_p.n12358 16.403
R4497 vp_p.n12347 vp_p.n12344 16.403
R4498 vp_p.n12333 vp_p.n12330 16.403
R4499 vp_p.n12319 vp_p.n12316 16.403
R4500 vp_p.n12305 vp_p.n12302 16.403
R4501 vp_p.n12291 vp_p.n12288 16.403
R4502 vp_p.n12277 vp_p.n12274 16.403
R4503 vp_p.n12263 vp_p.n12260 16.403
R4504 vp_p.n12249 vp_p.n12246 16.403
R4505 vp_p.n12235 vp_p.n12232 16.403
R4506 vp_p.n12221 vp_p.n12218 16.403
R4507 vp_p.n12207 vp_p.n12204 16.403
R4508 vp_p.n12193 vp_p.n12190 16.403
R4509 vp_p.n12179 vp_p.n12176 16.403
R4510 vp_p.n12165 vp_p.n12162 16.403
R4511 vp_p.n12151 vp_p.n12148 16.403
R4512 vp_p.n12137 vp_p.n12134 16.403
R4513 vp_p.n12123 vp_p.n12120 16.403
R4514 vp_p.n12109 vp_p.n12106 16.403
R4515 vp_p.n12095 vp_p.n12092 16.403
R4516 vp_p.n15808 vp_p.n15805 16.403
R4517 vp_p.n15794 vp_p.n15791 16.403
R4518 vp_p.n15780 vp_p.n15777 16.403
R4519 vp_p.n15766 vp_p.n15763 16.403
R4520 vp_p.n15752 vp_p.n15749 16.403
R4521 vp_p.n15738 vp_p.n15735 16.403
R4522 vp_p.n15724 vp_p.n15721 16.403
R4523 vp_p.n15710 vp_p.n15707 16.403
R4524 vp_p.n15696 vp_p.n15693 16.403
R4525 vp_p.n15682 vp_p.n15679 16.403
R4526 vp_p.n15668 vp_p.n15665 16.403
R4527 vp_p.n15654 vp_p.n15651 16.403
R4528 vp_p.n15640 vp_p.n15637 16.403
R4529 vp_p.n15626 vp_p.n15623 16.403
R4530 vp_p.n15612 vp_p.n15609 16.403
R4531 vp_p.n15598 vp_p.n15595 16.403
R4532 vp_p.n15584 vp_p.n15581 16.403
R4533 vp_p.n15570 vp_p.n15567 16.403
R4534 vp_p.n15556 vp_p.n15553 16.403
R4535 vp_p.n15542 vp_p.n15539 16.403
R4536 vp_p.n15528 vp_p.n15525 16.403
R4537 vp_p.n15514 vp_p.n15511 16.403
R4538 vp_p.n15500 vp_p.n15497 16.403
R4539 vp_p.n15486 vp_p.n15483 16.403
R4540 vp_p.n15472 vp_p.n15469 16.403
R4541 vp_p.n15458 vp_p.n15455 16.403
R4542 vp_p.n15444 vp_p.n15441 16.403
R4543 vp_p.n15430 vp_p.n15427 16.403
R4544 vp_p.n15416 vp_p.n15413 16.403
R4545 vp_p.n15402 vp_p.n15399 16.403
R4546 vp_p.n15388 vp_p.n15385 16.403
R4547 vp_p.n15374 vp_p.n15371 16.403
R4548 vp_p.n15360 vp_p.n15357 16.403
R4549 vp_p.n15346 vp_p.n15343 16.403
R4550 vp_p.n15332 vp_p.n15329 16.403
R4551 vp_p.n15318 vp_p.n15315 16.403
R4552 vp_p.n15304 vp_p.n15301 16.403
R4553 vp_p.n15290 vp_p.n15287 16.403
R4554 vp_p.n15276 vp_p.n15273 16.403
R4555 vp_p.n15262 vp_p.n15259 16.403
R4556 vp_p.n15248 vp_p.n15245 16.403
R4557 vp_p.n15234 vp_p.n15231 16.403
R4558 vp_p.n15220 vp_p.n15217 16.403
R4559 vp_p.n15206 vp_p.n15203 16.403
R4560 vp_p.n15192 vp_p.n15189 16.403
R4561 vp_p.n15178 vp_p.n15175 16.403
R4562 vp_p.n15164 vp_p.n15161 16.403
R4563 vp_p.n15150 vp_p.n15147 16.403
R4564 vp_p.n15136 vp_p.n15133 16.403
R4565 vp_p.n15122 vp_p.n15119 16.403
R4566 vp_p.n15108 vp_p.n15105 16.403
R4567 vp_p.n15094 vp_p.n15091 16.403
R4568 vp_p.n15080 vp_p.n15077 16.403
R4569 vp_p.n15066 vp_p.n15063 16.403
R4570 vp_p.n15052 vp_p.n15049 16.403
R4571 vp_p.n15038 vp_p.n15035 16.403
R4572 vp_p.n15024 vp_p.n15021 16.403
R4573 vp_p.n15010 vp_p.n15007 16.403
R4574 vp_p.n14996 vp_p.n14993 16.403
R4575 vp_p.n14982 vp_p.n14979 16.403
R4576 vp_p.n14968 vp_p.n14965 16.403
R4577 vp_p.n14954 vp_p.n14951 16.403
R4578 vp_p.n14940 vp_p.n14937 16.403
R4579 vp_p.n14926 vp_p.n14923 16.403
R4580 vp_p.n14912 vp_p.n14909 16.403
R4581 vp_p.n14898 vp_p.n14895 16.403
R4582 vp_p.n11581 vp_p.n11578 16.403
R4583 vp_p.n11567 vp_p.n11564 16.403
R4584 vp_p.n11553 vp_p.n11550 16.403
R4585 vp_p.n11539 vp_p.n11536 16.403
R4586 vp_p.n11525 vp_p.n11522 16.403
R4587 vp_p.n11511 vp_p.n11508 16.403
R4588 vp_p.n11497 vp_p.n11494 16.403
R4589 vp_p.n11483 vp_p.n11480 16.403
R4590 vp_p.n11469 vp_p.n11466 16.403
R4591 vp_p.n11455 vp_p.n11452 16.403
R4592 vp_p.n11441 vp_p.n11438 16.403
R4593 vp_p.n11427 vp_p.n11424 16.403
R4594 vp_p.n11413 vp_p.n11410 16.403
R4595 vp_p.n11399 vp_p.n11396 16.403
R4596 vp_p.n11385 vp_p.n11382 16.403
R4597 vp_p.n11371 vp_p.n11368 16.403
R4598 vp_p.n11357 vp_p.n11354 16.403
R4599 vp_p.n11343 vp_p.n11340 16.403
R4600 vp_p.n11329 vp_p.n11326 16.403
R4601 vp_p.n11315 vp_p.n11312 16.403
R4602 vp_p.n11301 vp_p.n11298 16.403
R4603 vp_p.n11287 vp_p.n11284 16.403
R4604 vp_p.n11273 vp_p.n11270 16.403
R4605 vp_p.n11259 vp_p.n11256 16.403
R4606 vp_p.n11245 vp_p.n11242 16.403
R4607 vp_p.n11231 vp_p.n11228 16.403
R4608 vp_p.n11217 vp_p.n11214 16.403
R4609 vp_p.n11203 vp_p.n11200 16.403
R4610 vp_p.n11189 vp_p.n11186 16.403
R4611 vp_p.n11175 vp_p.n11172 16.403
R4612 vp_p.n11161 vp_p.n11158 16.403
R4613 vp_p.n11147 vp_p.n11144 16.403
R4614 vp_p.n11133 vp_p.n11130 16.403
R4615 vp_p.n11119 vp_p.n11116 16.403
R4616 vp_p.n11105 vp_p.n11102 16.403
R4617 vp_p.n11091 vp_p.n11088 16.403
R4618 vp_p.n11077 vp_p.n11074 16.403
R4619 vp_p.n11063 vp_p.n11060 16.403
R4620 vp_p.n11049 vp_p.n11046 16.403
R4621 vp_p.n11035 vp_p.n11032 16.403
R4622 vp_p.n11021 vp_p.n11018 16.403
R4623 vp_p.n11007 vp_p.n11004 16.403
R4624 vp_p.n10993 vp_p.n10990 16.403
R4625 vp_p.n10979 vp_p.n10976 16.403
R4626 vp_p.n10965 vp_p.n10962 16.403
R4627 vp_p.n10951 vp_p.n10948 16.403
R4628 vp_p.n10937 vp_p.n10934 16.403
R4629 vp_p.n10923 vp_p.n10920 16.403
R4630 vp_p.n10909 vp_p.n10906 16.403
R4631 vp_p.n10895 vp_p.n10892 16.403
R4632 vp_p.n10881 vp_p.n10878 16.403
R4633 vp_p.n10867 vp_p.n10864 16.403
R4634 vp_p.n10853 vp_p.n10850 16.403
R4635 vp_p.n10839 vp_p.n10836 16.403
R4636 vp_p.n10825 vp_p.n10822 16.403
R4637 vp_p.n10811 vp_p.n10808 16.403
R4638 vp_p.n10797 vp_p.n10794 16.403
R4639 vp_p.n10783 vp_p.n10780 16.403
R4640 vp_p.n10769 vp_p.n10766 16.403
R4641 vp_p.n10755 vp_p.n10752 16.403
R4642 vp_p.n10741 vp_p.n10738 16.403
R4643 vp_p.n10727 vp_p.n10724 16.403
R4644 vp_p.n10713 vp_p.n10710 16.403
R4645 vp_p.n10699 vp_p.n10696 16.403
R4646 vp_p.n10685 vp_p.n10682 16.403
R4647 vp_p.n10671 vp_p.n10668 16.403
R4648 vp_p.n10657 vp_p.n10654 16.403
R4649 vp_p.n17250 vp_p.n17247 16.403
R4650 vp_p.n17236 vp_p.n17233 16.403
R4651 vp_p.n17222 vp_p.n17219 16.403
R4652 vp_p.n17208 vp_p.n17205 16.403
R4653 vp_p.n17194 vp_p.n17191 16.403
R4654 vp_p.n17180 vp_p.n17177 16.403
R4655 vp_p.n17166 vp_p.n17163 16.403
R4656 vp_p.n17152 vp_p.n17149 16.403
R4657 vp_p.n17138 vp_p.n17135 16.403
R4658 vp_p.n17124 vp_p.n17121 16.403
R4659 vp_p.n17110 vp_p.n17107 16.403
R4660 vp_p.n17096 vp_p.n17093 16.403
R4661 vp_p.n17082 vp_p.n17079 16.403
R4662 vp_p.n17068 vp_p.n17065 16.403
R4663 vp_p.n17054 vp_p.n17051 16.403
R4664 vp_p.n17040 vp_p.n17037 16.403
R4665 vp_p.n17026 vp_p.n17023 16.403
R4666 vp_p.n17012 vp_p.n17009 16.403
R4667 vp_p.n16998 vp_p.n16995 16.403
R4668 vp_p.n16984 vp_p.n16981 16.403
R4669 vp_p.n16970 vp_p.n16967 16.403
R4670 vp_p.n16956 vp_p.n16953 16.403
R4671 vp_p.n16942 vp_p.n16939 16.403
R4672 vp_p.n16928 vp_p.n16925 16.403
R4673 vp_p.n16914 vp_p.n16911 16.403
R4674 vp_p.n16900 vp_p.n16897 16.403
R4675 vp_p.n16886 vp_p.n16883 16.403
R4676 vp_p.n16872 vp_p.n16869 16.403
R4677 vp_p.n16858 vp_p.n16855 16.403
R4678 vp_p.n16844 vp_p.n16841 16.403
R4679 vp_p.n16830 vp_p.n16827 16.403
R4680 vp_p.n16816 vp_p.n16813 16.403
R4681 vp_p.n16802 vp_p.n16799 16.403
R4682 vp_p.n16788 vp_p.n16785 16.403
R4683 vp_p.n16774 vp_p.n16771 16.403
R4684 vp_p.n16760 vp_p.n16757 16.403
R4685 vp_p.n16746 vp_p.n16743 16.403
R4686 vp_p.n16732 vp_p.n16729 16.403
R4687 vp_p.n16718 vp_p.n16715 16.403
R4688 vp_p.n16704 vp_p.n16701 16.403
R4689 vp_p.n16690 vp_p.n16687 16.403
R4690 vp_p.n16676 vp_p.n16673 16.403
R4691 vp_p.n16662 vp_p.n16659 16.403
R4692 vp_p.n16648 vp_p.n16645 16.403
R4693 vp_p.n16634 vp_p.n16631 16.403
R4694 vp_p.n16620 vp_p.n16617 16.403
R4695 vp_p.n16606 vp_p.n16603 16.403
R4696 vp_p.n16592 vp_p.n16589 16.403
R4697 vp_p.n16578 vp_p.n16575 16.403
R4698 vp_p.n16564 vp_p.n16561 16.403
R4699 vp_p.n16550 vp_p.n16547 16.403
R4700 vp_p.n16536 vp_p.n16533 16.403
R4701 vp_p.n16522 vp_p.n16519 16.403
R4702 vp_p.n16508 vp_p.n16505 16.403
R4703 vp_p.n16494 vp_p.n16491 16.403
R4704 vp_p.n16480 vp_p.n16477 16.403
R4705 vp_p.n16466 vp_p.n16463 16.403
R4706 vp_p.n16452 vp_p.n16449 16.403
R4707 vp_p.n16438 vp_p.n16435 16.403
R4708 vp_p.n16424 vp_p.n16421 16.403
R4709 vp_p.n16410 vp_p.n16407 16.403
R4710 vp_p.n16396 vp_p.n16393 16.403
R4711 vp_p.n16382 vp_p.n16379 16.403
R4712 vp_p.n16368 vp_p.n16365 16.403
R4713 vp_p.n16354 vp_p.n16351 16.403
R4714 vp_p.n16340 vp_p.n16337 16.403
R4715 vp_p.n16326 vp_p.n16323 16.403
R4716 vp_p.n10158 vp_p.n10155 16.403
R4717 vp_p.n10144 vp_p.n10141 16.403
R4718 vp_p.n10130 vp_p.n10127 16.403
R4719 vp_p.n10116 vp_p.n10113 16.403
R4720 vp_p.n10102 vp_p.n10099 16.403
R4721 vp_p.n10088 vp_p.n10085 16.403
R4722 vp_p.n10074 vp_p.n10071 16.403
R4723 vp_p.n10060 vp_p.n10057 16.403
R4724 vp_p.n10046 vp_p.n10043 16.403
R4725 vp_p.n10032 vp_p.n10029 16.403
R4726 vp_p.n10018 vp_p.n10015 16.403
R4727 vp_p.n10004 vp_p.n10001 16.403
R4728 vp_p.n9990 vp_p.n9987 16.403
R4729 vp_p.n9976 vp_p.n9973 16.403
R4730 vp_p.n9962 vp_p.n9959 16.403
R4731 vp_p.n9948 vp_p.n9945 16.403
R4732 vp_p.n9934 vp_p.n9931 16.403
R4733 vp_p.n9920 vp_p.n9917 16.403
R4734 vp_p.n9906 vp_p.n9903 16.403
R4735 vp_p.n9892 vp_p.n9889 16.403
R4736 vp_p.n9878 vp_p.n9875 16.403
R4737 vp_p.n9864 vp_p.n9861 16.403
R4738 vp_p.n9850 vp_p.n9847 16.403
R4739 vp_p.n9836 vp_p.n9833 16.403
R4740 vp_p.n9822 vp_p.n9819 16.403
R4741 vp_p.n9808 vp_p.n9805 16.403
R4742 vp_p.n9794 vp_p.n9791 16.403
R4743 vp_p.n9780 vp_p.n9777 16.403
R4744 vp_p.n9766 vp_p.n9763 16.403
R4745 vp_p.n9752 vp_p.n9749 16.403
R4746 vp_p.n9738 vp_p.n9735 16.403
R4747 vp_p.n9724 vp_p.n9721 16.403
R4748 vp_p.n9710 vp_p.n9707 16.403
R4749 vp_p.n9696 vp_p.n9693 16.403
R4750 vp_p.n9682 vp_p.n9679 16.403
R4751 vp_p.n9668 vp_p.n9665 16.403
R4752 vp_p.n9654 vp_p.n9651 16.403
R4753 vp_p.n9640 vp_p.n9637 16.403
R4754 vp_p.n9626 vp_p.n9623 16.403
R4755 vp_p.n9612 vp_p.n9609 16.403
R4756 vp_p.n9598 vp_p.n9595 16.403
R4757 vp_p.n9584 vp_p.n9581 16.403
R4758 vp_p.n9570 vp_p.n9567 16.403
R4759 vp_p.n9556 vp_p.n9553 16.403
R4760 vp_p.n9542 vp_p.n9539 16.403
R4761 vp_p.n9528 vp_p.n9525 16.403
R4762 vp_p.n9514 vp_p.n9511 16.403
R4763 vp_p.n9500 vp_p.n9497 16.403
R4764 vp_p.n9486 vp_p.n9483 16.403
R4765 vp_p.n9472 vp_p.n9469 16.403
R4766 vp_p.n9458 vp_p.n9455 16.403
R4767 vp_p.n9444 vp_p.n9441 16.403
R4768 vp_p.n9430 vp_p.n9427 16.403
R4769 vp_p.n9416 vp_p.n9413 16.403
R4770 vp_p.n9402 vp_p.n9399 16.403
R4771 vp_p.n9388 vp_p.n9385 16.403
R4772 vp_p.n9374 vp_p.n9371 16.403
R4773 vp_p.n9360 vp_p.n9357 16.403
R4774 vp_p.n9346 vp_p.n9343 16.403
R4775 vp_p.n9332 vp_p.n9329 16.403
R4776 vp_p.n9318 vp_p.n9315 16.403
R4777 vp_p.n9304 vp_p.n9301 16.403
R4778 vp_p.n9290 vp_p.n9287 16.403
R4779 vp_p.n9276 vp_p.n9273 16.403
R4780 vp_p.n9262 vp_p.n9259 16.403
R4781 vp_p.n9248 vp_p.n9245 16.403
R4782 vp_p.n9234 vp_p.n9231 16.403
R4783 vp_p.n9220 vp_p.n9217 16.403
R4784 vp_p.n18691 vp_p.n18688 16.403
R4785 vp_p.n18677 vp_p.n18674 16.403
R4786 vp_p.n18663 vp_p.n18660 16.403
R4787 vp_p.n18649 vp_p.n18646 16.403
R4788 vp_p.n18635 vp_p.n18632 16.403
R4789 vp_p.n18621 vp_p.n18618 16.403
R4790 vp_p.n18607 vp_p.n18604 16.403
R4791 vp_p.n18593 vp_p.n18590 16.403
R4792 vp_p.n18579 vp_p.n18576 16.403
R4793 vp_p.n18565 vp_p.n18562 16.403
R4794 vp_p.n18551 vp_p.n18548 16.403
R4795 vp_p.n18537 vp_p.n18534 16.403
R4796 vp_p.n18523 vp_p.n18520 16.403
R4797 vp_p.n18509 vp_p.n18506 16.403
R4798 vp_p.n18495 vp_p.n18492 16.403
R4799 vp_p.n18481 vp_p.n18478 16.403
R4800 vp_p.n18467 vp_p.n18464 16.403
R4801 vp_p.n18453 vp_p.n18450 16.403
R4802 vp_p.n18439 vp_p.n18436 16.403
R4803 vp_p.n18425 vp_p.n18422 16.403
R4804 vp_p.n18411 vp_p.n18408 16.403
R4805 vp_p.n18397 vp_p.n18394 16.403
R4806 vp_p.n18383 vp_p.n18380 16.403
R4807 vp_p.n18369 vp_p.n18366 16.403
R4808 vp_p.n18355 vp_p.n18352 16.403
R4809 vp_p.n18341 vp_p.n18338 16.403
R4810 vp_p.n18327 vp_p.n18324 16.403
R4811 vp_p.n18313 vp_p.n18310 16.403
R4812 vp_p.n18299 vp_p.n18296 16.403
R4813 vp_p.n18285 vp_p.n18282 16.403
R4814 vp_p.n18271 vp_p.n18268 16.403
R4815 vp_p.n18257 vp_p.n18254 16.403
R4816 vp_p.n18243 vp_p.n18240 16.403
R4817 vp_p.n18229 vp_p.n18226 16.403
R4818 vp_p.n18215 vp_p.n18212 16.403
R4819 vp_p.n18201 vp_p.n18198 16.403
R4820 vp_p.n18187 vp_p.n18184 16.403
R4821 vp_p.n18173 vp_p.n18170 16.403
R4822 vp_p.n18159 vp_p.n18156 16.403
R4823 vp_p.n18145 vp_p.n18142 16.403
R4824 vp_p.n18131 vp_p.n18128 16.403
R4825 vp_p.n18117 vp_p.n18114 16.403
R4826 vp_p.n18103 vp_p.n18100 16.403
R4827 vp_p.n18089 vp_p.n18086 16.403
R4828 vp_p.n18075 vp_p.n18072 16.403
R4829 vp_p.n18061 vp_p.n18058 16.403
R4830 vp_p.n18047 vp_p.n18044 16.403
R4831 vp_p.n18033 vp_p.n18030 16.403
R4832 vp_p.n18019 vp_p.n18016 16.403
R4833 vp_p.n18005 vp_p.n18002 16.403
R4834 vp_p.n17991 vp_p.n17988 16.403
R4835 vp_p.n17977 vp_p.n17974 16.403
R4836 vp_p.n17963 vp_p.n17960 16.403
R4837 vp_p.n17949 vp_p.n17946 16.403
R4838 vp_p.n17935 vp_p.n17932 16.403
R4839 vp_p.n17921 vp_p.n17918 16.403
R4840 vp_p.n17907 vp_p.n17904 16.403
R4841 vp_p.n17893 vp_p.n17890 16.403
R4842 vp_p.n17879 vp_p.n17876 16.403
R4843 vp_p.n17865 vp_p.n17862 16.403
R4844 vp_p.n17851 vp_p.n17848 16.403
R4845 vp_p.n17837 vp_p.n17834 16.403
R4846 vp_p.n17823 vp_p.n17820 16.403
R4847 vp_p.n17809 vp_p.n17806 16.403
R4848 vp_p.n17795 vp_p.n17792 16.403
R4849 vp_p.n17781 vp_p.n17778 16.403
R4850 vp_p.n17767 vp_p.n17764 16.403
R4851 vp_p.n17753 vp_p.n17750 16.403
R4852 vp_p.n1426 vp_p.n1423 16.403
R4853 vp_p.n1412 vp_p.n1409 16.403
R4854 vp_p.n1398 vp_p.n1395 16.403
R4855 vp_p.n1384 vp_p.n1381 16.403
R4856 vp_p.n1370 vp_p.n1367 16.403
R4857 vp_p.n1356 vp_p.n1353 16.403
R4858 vp_p.n1342 vp_p.n1339 16.403
R4859 vp_p.n1328 vp_p.n1325 16.403
R4860 vp_p.n1314 vp_p.n1311 16.403
R4861 vp_p.n1300 vp_p.n1297 16.403
R4862 vp_p.n1286 vp_p.n1283 16.403
R4863 vp_p.n1272 vp_p.n1269 16.403
R4864 vp_p.n1258 vp_p.n1255 16.403
R4865 vp_p.n1244 vp_p.n1241 16.403
R4866 vp_p.n1230 vp_p.n1227 16.403
R4867 vp_p.n1216 vp_p.n1213 16.403
R4868 vp_p.n1202 vp_p.n1199 16.403
R4869 vp_p.n1188 vp_p.n1185 16.403
R4870 vp_p.n1174 vp_p.n1171 16.403
R4871 vp_p.n1160 vp_p.n1157 16.403
R4872 vp_p.n1146 vp_p.n1143 16.403
R4873 vp_p.n1132 vp_p.n1129 16.403
R4874 vp_p.n1118 vp_p.n1115 16.403
R4875 vp_p.n1104 vp_p.n1101 16.403
R4876 vp_p.n1090 vp_p.n1087 16.403
R4877 vp_p.n1076 vp_p.n1073 16.403
R4878 vp_p.n1062 vp_p.n1059 16.403
R4879 vp_p.n1048 vp_p.n1045 16.403
R4880 vp_p.n1034 vp_p.n1031 16.403
R4881 vp_p.n1020 vp_p.n1017 16.403
R4882 vp_p.n1006 vp_p.n1003 16.403
R4883 vp_p.n992 vp_p.n989 16.403
R4884 vp_p.n978 vp_p.n975 16.403
R4885 vp_p.n964 vp_p.n961 16.403
R4886 vp_p.n950 vp_p.n947 16.403
R4887 vp_p.n936 vp_p.n933 16.403
R4888 vp_p.n922 vp_p.n919 16.403
R4889 vp_p.n908 vp_p.n905 16.403
R4890 vp_p.n894 vp_p.n891 16.403
R4891 vp_p.n880 vp_p.n877 16.403
R4892 vp_p.n866 vp_p.n863 16.403
R4893 vp_p.n852 vp_p.n849 16.403
R4894 vp_p.n838 vp_p.n835 16.403
R4895 vp_p.n824 vp_p.n821 16.403
R4896 vp_p.n810 vp_p.n807 16.403
R4897 vp_p.n796 vp_p.n793 16.403
R4898 vp_p.n782 vp_p.n779 16.403
R4899 vp_p.n768 vp_p.n765 16.403
R4900 vp_p.n754 vp_p.n751 16.403
R4901 vp_p.n740 vp_p.n737 16.403
R4902 vp_p.n726 vp_p.n723 16.403
R4903 vp_p.n712 vp_p.n709 16.403
R4904 vp_p.n698 vp_p.n695 16.403
R4905 vp_p.n684 vp_p.n681 16.403
R4906 vp_p.n670 vp_p.n667 16.403
R4907 vp_p.n656 vp_p.n653 16.403
R4908 vp_p.n642 vp_p.n639 16.403
R4909 vp_p.n628 vp_p.n625 16.403
R4910 vp_p.n614 vp_p.n611 16.403
R4911 vp_p.n600 vp_p.n597 16.403
R4912 vp_p.n586 vp_p.n583 16.403
R4913 vp_p.n572 vp_p.n569 16.403
R4914 vp_p.n558 vp_p.n555 16.403
R4915 vp_p.n544 vp_p.n541 16.403
R4916 vp_p.n530 vp_p.n527 16.403
R4917 vp_p.n516 vp_p.n513 16.403
R4918 vp_p.n502 vp_p.n499 16.403
R4919 vp_p.n488 vp_p.n485 16.403
R4920 vp_p.n474 vp_p.n471 16.403
R4921 vp_p.n20131 vp_p.n20128 16.403
R4922 vp_p.n20117 vp_p.n20114 16.403
R4923 vp_p.n20103 vp_p.n20100 16.403
R4924 vp_p.n20089 vp_p.n20086 16.403
R4925 vp_p.n20075 vp_p.n20072 16.403
R4926 vp_p.n20061 vp_p.n20058 16.403
R4927 vp_p.n20047 vp_p.n20044 16.403
R4928 vp_p.n20033 vp_p.n20030 16.403
R4929 vp_p.n20019 vp_p.n20016 16.403
R4930 vp_p.n20005 vp_p.n20002 16.403
R4931 vp_p.n19991 vp_p.n19988 16.403
R4932 vp_p.n19977 vp_p.n19974 16.403
R4933 vp_p.n19963 vp_p.n19960 16.403
R4934 vp_p.n19949 vp_p.n19946 16.403
R4935 vp_p.n19935 vp_p.n19932 16.403
R4936 vp_p.n19921 vp_p.n19918 16.403
R4937 vp_p.n19907 vp_p.n19904 16.403
R4938 vp_p.n19893 vp_p.n19890 16.403
R4939 vp_p.n19879 vp_p.n19876 16.403
R4940 vp_p.n19865 vp_p.n19862 16.403
R4941 vp_p.n19851 vp_p.n19848 16.403
R4942 vp_p.n19837 vp_p.n19834 16.403
R4943 vp_p.n19823 vp_p.n19820 16.403
R4944 vp_p.n19809 vp_p.n19806 16.403
R4945 vp_p.n19795 vp_p.n19792 16.403
R4946 vp_p.n19781 vp_p.n19778 16.403
R4947 vp_p.n19767 vp_p.n19764 16.403
R4948 vp_p.n19753 vp_p.n19750 16.403
R4949 vp_p.n19739 vp_p.n19736 16.403
R4950 vp_p.n19725 vp_p.n19722 16.403
R4951 vp_p.n19711 vp_p.n19708 16.403
R4952 vp_p.n19697 vp_p.n19694 16.403
R4953 vp_p.n19683 vp_p.n19680 16.403
R4954 vp_p.n19669 vp_p.n19666 16.403
R4955 vp_p.n19655 vp_p.n19652 16.403
R4956 vp_p.n19641 vp_p.n19638 16.403
R4957 vp_p.n19627 vp_p.n19624 16.403
R4958 vp_p.n19613 vp_p.n19610 16.403
R4959 vp_p.n19599 vp_p.n19596 16.403
R4960 vp_p.n19585 vp_p.n19582 16.403
R4961 vp_p.n19571 vp_p.n19568 16.403
R4962 vp_p.n19557 vp_p.n19554 16.403
R4963 vp_p.n19543 vp_p.n19540 16.403
R4964 vp_p.n19529 vp_p.n19526 16.403
R4965 vp_p.n19515 vp_p.n19512 16.403
R4966 vp_p.n19501 vp_p.n19498 16.403
R4967 vp_p.n19487 vp_p.n19484 16.403
R4968 vp_p.n19473 vp_p.n19470 16.403
R4969 vp_p.n19459 vp_p.n19456 16.403
R4970 vp_p.n19445 vp_p.n19442 16.403
R4971 vp_p.n19431 vp_p.n19428 16.403
R4972 vp_p.n19417 vp_p.n19414 16.403
R4973 vp_p.n19403 vp_p.n19400 16.403
R4974 vp_p.n19389 vp_p.n19386 16.403
R4975 vp_p.n19375 vp_p.n19372 16.403
R4976 vp_p.n19361 vp_p.n19358 16.403
R4977 vp_p.n19347 vp_p.n19344 16.403
R4978 vp_p.n19333 vp_p.n19330 16.403
R4979 vp_p.n19319 vp_p.n19316 16.403
R4980 vp_p.n19305 vp_p.n19302 16.403
R4981 vp_p.n19291 vp_p.n19288 16.403
R4982 vp_p.n19277 vp_p.n19274 16.403
R4983 vp_p.n19263 vp_p.n19260 16.403
R4984 vp_p.n19249 vp_p.n19246 16.403
R4985 vp_p.n19235 vp_p.n19232 16.403
R4986 vp_p.n19221 vp_p.n19218 16.403
R4987 vp_p.n19207 vp_p.n19204 16.403
R4988 vp_p.n19193 vp_p.n19190 16.403
R4989 vp_p.n19179 vp_p.n19176 16.403
R4990 vp_p.n2866 vp_p.n2863 16.403
R4991 vp_p.n2852 vp_p.n2849 16.403
R4992 vp_p.n2838 vp_p.n2835 16.403
R4993 vp_p.n2824 vp_p.n2821 16.403
R4994 vp_p.n2810 vp_p.n2807 16.403
R4995 vp_p.n2796 vp_p.n2793 16.403
R4996 vp_p.n2782 vp_p.n2779 16.403
R4997 vp_p.n2768 vp_p.n2765 16.403
R4998 vp_p.n2754 vp_p.n2751 16.403
R4999 vp_p.n2740 vp_p.n2737 16.403
R5000 vp_p.n2726 vp_p.n2723 16.403
R5001 vp_p.n2712 vp_p.n2709 16.403
R5002 vp_p.n2698 vp_p.n2695 16.403
R5003 vp_p.n2684 vp_p.n2681 16.403
R5004 vp_p.n2670 vp_p.n2667 16.403
R5005 vp_p.n2656 vp_p.n2653 16.403
R5006 vp_p.n2642 vp_p.n2639 16.403
R5007 vp_p.n2628 vp_p.n2625 16.403
R5008 vp_p.n2614 vp_p.n2611 16.403
R5009 vp_p.n2600 vp_p.n2597 16.403
R5010 vp_p.n2586 vp_p.n2583 16.403
R5011 vp_p.n2572 vp_p.n2569 16.403
R5012 vp_p.n2558 vp_p.n2555 16.403
R5013 vp_p.n2544 vp_p.n2541 16.403
R5014 vp_p.n2530 vp_p.n2527 16.403
R5015 vp_p.n2516 vp_p.n2513 16.403
R5016 vp_p.n2502 vp_p.n2499 16.403
R5017 vp_p.n2488 vp_p.n2485 16.403
R5018 vp_p.n2474 vp_p.n2471 16.403
R5019 vp_p.n2460 vp_p.n2457 16.403
R5020 vp_p.n2446 vp_p.n2443 16.403
R5021 vp_p.n2432 vp_p.n2429 16.403
R5022 vp_p.n2418 vp_p.n2415 16.403
R5023 vp_p.n2404 vp_p.n2401 16.403
R5024 vp_p.n2390 vp_p.n2387 16.403
R5025 vp_p.n2376 vp_p.n2373 16.403
R5026 vp_p.n2362 vp_p.n2359 16.403
R5027 vp_p.n2348 vp_p.n2345 16.403
R5028 vp_p.n2334 vp_p.n2331 16.403
R5029 vp_p.n2320 vp_p.n2317 16.403
R5030 vp_p.n2306 vp_p.n2303 16.403
R5031 vp_p.n2292 vp_p.n2289 16.403
R5032 vp_p.n2278 vp_p.n2275 16.403
R5033 vp_p.n2264 vp_p.n2261 16.403
R5034 vp_p.n2250 vp_p.n2247 16.403
R5035 vp_p.n2236 vp_p.n2233 16.403
R5036 vp_p.n2222 vp_p.n2219 16.403
R5037 vp_p.n2208 vp_p.n2205 16.403
R5038 vp_p.n2194 vp_p.n2191 16.403
R5039 vp_p.n2180 vp_p.n2177 16.403
R5040 vp_p.n2166 vp_p.n2163 16.403
R5041 vp_p.n2152 vp_p.n2149 16.403
R5042 vp_p.n2138 vp_p.n2135 16.403
R5043 vp_p.n2124 vp_p.n2121 16.403
R5044 vp_p.n2110 vp_p.n2107 16.403
R5045 vp_p.n2096 vp_p.n2093 16.403
R5046 vp_p.n2082 vp_p.n2079 16.403
R5047 vp_p.n2068 vp_p.n2065 16.403
R5048 vp_p.n2054 vp_p.n2051 16.403
R5049 vp_p.n2040 vp_p.n2037 16.403
R5050 vp_p.n2026 vp_p.n2023 16.403
R5051 vp_p.n2012 vp_p.n2009 16.403
R5052 vp_p.n1998 vp_p.n1995 16.403
R5053 vp_p.n1984 vp_p.n1981 16.403
R5054 vp_p.n1970 vp_p.n1967 16.403
R5055 vp_p.n1956 vp_p.n1953 16.403
R5056 vp_p.n1942 vp_p.n1939 16.403
R5057 vp_p.n1928 vp_p.n1925 16.403
R5058 vp_p.n1914 vp_p.n1911 16.403
R5059 vp_p.n1900 vp_p.n1897 16.403
R5060 vp_p.n21570 vp_p.n21567 16.403
R5061 vp_p.n21556 vp_p.n21553 16.403
R5062 vp_p.n21542 vp_p.n21539 16.403
R5063 vp_p.n21528 vp_p.n21525 16.403
R5064 vp_p.n21514 vp_p.n21511 16.403
R5065 vp_p.n21500 vp_p.n21497 16.403
R5066 vp_p.n21486 vp_p.n21483 16.403
R5067 vp_p.n21472 vp_p.n21469 16.403
R5068 vp_p.n21458 vp_p.n21455 16.403
R5069 vp_p.n21444 vp_p.n21441 16.403
R5070 vp_p.n21430 vp_p.n21427 16.403
R5071 vp_p.n21416 vp_p.n21413 16.403
R5072 vp_p.n21402 vp_p.n21399 16.403
R5073 vp_p.n21388 vp_p.n21385 16.403
R5074 vp_p.n21374 vp_p.n21371 16.403
R5075 vp_p.n21360 vp_p.n21357 16.403
R5076 vp_p.n21346 vp_p.n21343 16.403
R5077 vp_p.n21332 vp_p.n21329 16.403
R5078 vp_p.n21318 vp_p.n21315 16.403
R5079 vp_p.n21304 vp_p.n21301 16.403
R5080 vp_p.n21290 vp_p.n21287 16.403
R5081 vp_p.n21276 vp_p.n21273 16.403
R5082 vp_p.n21262 vp_p.n21259 16.403
R5083 vp_p.n21248 vp_p.n21245 16.403
R5084 vp_p.n21234 vp_p.n21231 16.403
R5085 vp_p.n21220 vp_p.n21217 16.403
R5086 vp_p.n21206 vp_p.n21203 16.403
R5087 vp_p.n21192 vp_p.n21189 16.403
R5088 vp_p.n21178 vp_p.n21175 16.403
R5089 vp_p.n21164 vp_p.n21161 16.403
R5090 vp_p.n21150 vp_p.n21147 16.403
R5091 vp_p.n21136 vp_p.n21133 16.403
R5092 vp_p.n21122 vp_p.n21119 16.403
R5093 vp_p.n21108 vp_p.n21105 16.403
R5094 vp_p.n21094 vp_p.n21091 16.403
R5095 vp_p.n21080 vp_p.n21077 16.403
R5096 vp_p.n21066 vp_p.n21063 16.403
R5097 vp_p.n21052 vp_p.n21049 16.403
R5098 vp_p.n21038 vp_p.n21035 16.403
R5099 vp_p.n21024 vp_p.n21021 16.403
R5100 vp_p.n21010 vp_p.n21007 16.403
R5101 vp_p.n20996 vp_p.n20993 16.403
R5102 vp_p.n20982 vp_p.n20979 16.403
R5103 vp_p.n20968 vp_p.n20965 16.403
R5104 vp_p.n20954 vp_p.n20951 16.403
R5105 vp_p.n20940 vp_p.n20937 16.403
R5106 vp_p.n20926 vp_p.n20923 16.403
R5107 vp_p.n20912 vp_p.n20909 16.403
R5108 vp_p.n20898 vp_p.n20895 16.403
R5109 vp_p.n20884 vp_p.n20881 16.403
R5110 vp_p.n20870 vp_p.n20867 16.403
R5111 vp_p.n20856 vp_p.n20853 16.403
R5112 vp_p.n20842 vp_p.n20839 16.403
R5113 vp_p.n20828 vp_p.n20825 16.403
R5114 vp_p.n20814 vp_p.n20811 16.403
R5115 vp_p.n20800 vp_p.n20797 16.403
R5116 vp_p.n20786 vp_p.n20783 16.403
R5117 vp_p.n20772 vp_p.n20769 16.403
R5118 vp_p.n20758 vp_p.n20755 16.403
R5119 vp_p.n20744 vp_p.n20741 16.403
R5120 vp_p.n20730 vp_p.n20727 16.403
R5121 vp_p.n20716 vp_p.n20713 16.403
R5122 vp_p.n20702 vp_p.n20699 16.403
R5123 vp_p.n20688 vp_p.n20685 16.403
R5124 vp_p.n20674 vp_p.n20671 16.403
R5125 vp_p.n20660 vp_p.n20657 16.403
R5126 vp_p.n20646 vp_p.n20643 16.403
R5127 vp_p.n20632 vp_p.n20629 16.403
R5128 vp_p.n20618 vp_p.n20615 16.403
R5129 vp_p.n20604 vp_p.n20601 16.403
R5130 vp_p.n4305 vp_p.n4302 16.403
R5131 vp_p.n4291 vp_p.n4288 16.403
R5132 vp_p.n4277 vp_p.n4274 16.403
R5133 vp_p.n4263 vp_p.n4260 16.403
R5134 vp_p.n4249 vp_p.n4246 16.403
R5135 vp_p.n4235 vp_p.n4232 16.403
R5136 vp_p.n4221 vp_p.n4218 16.403
R5137 vp_p.n4207 vp_p.n4204 16.403
R5138 vp_p.n4193 vp_p.n4190 16.403
R5139 vp_p.n4179 vp_p.n4176 16.403
R5140 vp_p.n4165 vp_p.n4162 16.403
R5141 vp_p.n4151 vp_p.n4148 16.403
R5142 vp_p.n4137 vp_p.n4134 16.403
R5143 vp_p.n4123 vp_p.n4120 16.403
R5144 vp_p.n4109 vp_p.n4106 16.403
R5145 vp_p.n4095 vp_p.n4092 16.403
R5146 vp_p.n4081 vp_p.n4078 16.403
R5147 vp_p.n4067 vp_p.n4064 16.403
R5148 vp_p.n4053 vp_p.n4050 16.403
R5149 vp_p.n4039 vp_p.n4036 16.403
R5150 vp_p.n4025 vp_p.n4022 16.403
R5151 vp_p.n4011 vp_p.n4008 16.403
R5152 vp_p.n3997 vp_p.n3994 16.403
R5153 vp_p.n3983 vp_p.n3980 16.403
R5154 vp_p.n3969 vp_p.n3966 16.403
R5155 vp_p.n3955 vp_p.n3952 16.403
R5156 vp_p.n3941 vp_p.n3938 16.403
R5157 vp_p.n3927 vp_p.n3924 16.403
R5158 vp_p.n3913 vp_p.n3910 16.403
R5159 vp_p.n3899 vp_p.n3896 16.403
R5160 vp_p.n3885 vp_p.n3882 16.403
R5161 vp_p.n3871 vp_p.n3868 16.403
R5162 vp_p.n3857 vp_p.n3854 16.403
R5163 vp_p.n3843 vp_p.n3840 16.403
R5164 vp_p.n3829 vp_p.n3826 16.403
R5165 vp_p.n3815 vp_p.n3812 16.403
R5166 vp_p.n3801 vp_p.n3798 16.403
R5167 vp_p.n3787 vp_p.n3784 16.403
R5168 vp_p.n3773 vp_p.n3770 16.403
R5169 vp_p.n3759 vp_p.n3756 16.403
R5170 vp_p.n3745 vp_p.n3742 16.403
R5171 vp_p.n3731 vp_p.n3728 16.403
R5172 vp_p.n3717 vp_p.n3714 16.403
R5173 vp_p.n3703 vp_p.n3700 16.403
R5174 vp_p.n3689 vp_p.n3686 16.403
R5175 vp_p.n3675 vp_p.n3672 16.403
R5176 vp_p.n3661 vp_p.n3658 16.403
R5177 vp_p.n3647 vp_p.n3644 16.403
R5178 vp_p.n3633 vp_p.n3630 16.403
R5179 vp_p.n3619 vp_p.n3616 16.403
R5180 vp_p.n3605 vp_p.n3602 16.403
R5181 vp_p.n3591 vp_p.n3588 16.403
R5182 vp_p.n3577 vp_p.n3574 16.403
R5183 vp_p.n3563 vp_p.n3560 16.403
R5184 vp_p.n3549 vp_p.n3546 16.403
R5185 vp_p.n3535 vp_p.n3532 16.403
R5186 vp_p.n3521 vp_p.n3518 16.403
R5187 vp_p.n3507 vp_p.n3504 16.403
R5188 vp_p.n3493 vp_p.n3490 16.403
R5189 vp_p.n3479 vp_p.n3476 16.403
R5190 vp_p.n3465 vp_p.n3462 16.403
R5191 vp_p.n3451 vp_p.n3448 16.403
R5192 vp_p.n3437 vp_p.n3434 16.403
R5193 vp_p.n3423 vp_p.n3420 16.403
R5194 vp_p.n3409 vp_p.n3406 16.403
R5195 vp_p.n3395 vp_p.n3392 16.403
R5196 vp_p.n3381 vp_p.n3378 16.403
R5197 vp_p.n3367 vp_p.n3364 16.403
R5198 vp_p.n3353 vp_p.n3350 16.403
R5199 vp_p.n3339 vp_p.n3336 16.403
R5200 vp_p.n3325 vp_p.n3322 16.403
R5201 vp_p.n23008 vp_p.n23005 16.403
R5202 vp_p.n22994 vp_p.n22991 16.403
R5203 vp_p.n22980 vp_p.n22977 16.403
R5204 vp_p.n22966 vp_p.n22963 16.403
R5205 vp_p.n22952 vp_p.n22949 16.403
R5206 vp_p.n22938 vp_p.n22935 16.403
R5207 vp_p.n22924 vp_p.n22921 16.403
R5208 vp_p.n22910 vp_p.n22907 16.403
R5209 vp_p.n22896 vp_p.n22893 16.403
R5210 vp_p.n22882 vp_p.n22879 16.403
R5211 vp_p.n22868 vp_p.n22865 16.403
R5212 vp_p.n22854 vp_p.n22851 16.403
R5213 vp_p.n22840 vp_p.n22837 16.403
R5214 vp_p.n22826 vp_p.n22823 16.403
R5215 vp_p.n22812 vp_p.n22809 16.403
R5216 vp_p.n22798 vp_p.n22795 16.403
R5217 vp_p.n22784 vp_p.n22781 16.403
R5218 vp_p.n22770 vp_p.n22767 16.403
R5219 vp_p.n22756 vp_p.n22753 16.403
R5220 vp_p.n22742 vp_p.n22739 16.403
R5221 vp_p.n22728 vp_p.n22725 16.403
R5222 vp_p.n22714 vp_p.n22711 16.403
R5223 vp_p.n22700 vp_p.n22697 16.403
R5224 vp_p.n22686 vp_p.n22683 16.403
R5225 vp_p.n22672 vp_p.n22669 16.403
R5226 vp_p.n22658 vp_p.n22655 16.403
R5227 vp_p.n22644 vp_p.n22641 16.403
R5228 vp_p.n22630 vp_p.n22627 16.403
R5229 vp_p.n22616 vp_p.n22613 16.403
R5230 vp_p.n22602 vp_p.n22599 16.403
R5231 vp_p.n22588 vp_p.n22585 16.403
R5232 vp_p.n22574 vp_p.n22571 16.403
R5233 vp_p.n22560 vp_p.n22557 16.403
R5234 vp_p.n22546 vp_p.n22543 16.403
R5235 vp_p.n22532 vp_p.n22529 16.403
R5236 vp_p.n22518 vp_p.n22515 16.403
R5237 vp_p.n22504 vp_p.n22501 16.403
R5238 vp_p.n22490 vp_p.n22487 16.403
R5239 vp_p.n22476 vp_p.n22473 16.403
R5240 vp_p.n22462 vp_p.n22459 16.403
R5241 vp_p.n22448 vp_p.n22445 16.403
R5242 vp_p.n22434 vp_p.n22431 16.403
R5243 vp_p.n22420 vp_p.n22417 16.403
R5244 vp_p.n22406 vp_p.n22403 16.403
R5245 vp_p.n22392 vp_p.n22389 16.403
R5246 vp_p.n22378 vp_p.n22375 16.403
R5247 vp_p.n22364 vp_p.n22361 16.403
R5248 vp_p.n22350 vp_p.n22347 16.403
R5249 vp_p.n22336 vp_p.n22333 16.403
R5250 vp_p.n22322 vp_p.n22319 16.403
R5251 vp_p.n22308 vp_p.n22305 16.403
R5252 vp_p.n22294 vp_p.n22291 16.403
R5253 vp_p.n22280 vp_p.n22277 16.403
R5254 vp_p.n22266 vp_p.n22263 16.403
R5255 vp_p.n22252 vp_p.n22249 16.403
R5256 vp_p.n22238 vp_p.n22235 16.403
R5257 vp_p.n22224 vp_p.n22221 16.403
R5258 vp_p.n22210 vp_p.n22207 16.403
R5259 vp_p.n22196 vp_p.n22193 16.403
R5260 vp_p.n22182 vp_p.n22179 16.403
R5261 vp_p.n22168 vp_p.n22165 16.403
R5262 vp_p.n22154 vp_p.n22151 16.403
R5263 vp_p.n22140 vp_p.n22137 16.403
R5264 vp_p.n22126 vp_p.n22123 16.403
R5265 vp_p.n22112 vp_p.n22109 16.403
R5266 vp_p.n22098 vp_p.n22095 16.403
R5267 vp_p.n22084 vp_p.n22081 16.403
R5268 vp_p.n22070 vp_p.n22067 16.403
R5269 vp_p.n22056 vp_p.n22053 16.403
R5270 vp_p.n22042 vp_p.n22039 16.403
R5271 vp_p.n22028 vp_p.n22025 16.403
R5272 vp_p.n5743 vp_p.n5740 16.403
R5273 vp_p.n5729 vp_p.n5726 16.403
R5274 vp_p.n5715 vp_p.n5712 16.403
R5275 vp_p.n5701 vp_p.n5698 16.403
R5276 vp_p.n5687 vp_p.n5684 16.403
R5277 vp_p.n5673 vp_p.n5670 16.403
R5278 vp_p.n5659 vp_p.n5656 16.403
R5279 vp_p.n5645 vp_p.n5642 16.403
R5280 vp_p.n5631 vp_p.n5628 16.403
R5281 vp_p.n5617 vp_p.n5614 16.403
R5282 vp_p.n5603 vp_p.n5600 16.403
R5283 vp_p.n5589 vp_p.n5586 16.403
R5284 vp_p.n5575 vp_p.n5572 16.403
R5285 vp_p.n5561 vp_p.n5558 16.403
R5286 vp_p.n5547 vp_p.n5544 16.403
R5287 vp_p.n5533 vp_p.n5530 16.403
R5288 vp_p.n5519 vp_p.n5516 16.403
R5289 vp_p.n5505 vp_p.n5502 16.403
R5290 vp_p.n5491 vp_p.n5488 16.403
R5291 vp_p.n5477 vp_p.n5474 16.403
R5292 vp_p.n5463 vp_p.n5460 16.403
R5293 vp_p.n5449 vp_p.n5446 16.403
R5294 vp_p.n5435 vp_p.n5432 16.403
R5295 vp_p.n5421 vp_p.n5418 16.403
R5296 vp_p.n5407 vp_p.n5404 16.403
R5297 vp_p.n5393 vp_p.n5390 16.403
R5298 vp_p.n5379 vp_p.n5376 16.403
R5299 vp_p.n5365 vp_p.n5362 16.403
R5300 vp_p.n5351 vp_p.n5348 16.403
R5301 vp_p.n5337 vp_p.n5334 16.403
R5302 vp_p.n5323 vp_p.n5320 16.403
R5303 vp_p.n5309 vp_p.n5306 16.403
R5304 vp_p.n5295 vp_p.n5292 16.403
R5305 vp_p.n5281 vp_p.n5278 16.403
R5306 vp_p.n5267 vp_p.n5264 16.403
R5307 vp_p.n5253 vp_p.n5250 16.403
R5308 vp_p.n5239 vp_p.n5236 16.403
R5309 vp_p.n5225 vp_p.n5222 16.403
R5310 vp_p.n5211 vp_p.n5208 16.403
R5311 vp_p.n5197 vp_p.n5194 16.403
R5312 vp_p.n5183 vp_p.n5180 16.403
R5313 vp_p.n5169 vp_p.n5166 16.403
R5314 vp_p.n5155 vp_p.n5152 16.403
R5315 vp_p.n5141 vp_p.n5138 16.403
R5316 vp_p.n5127 vp_p.n5124 16.403
R5317 vp_p.n5113 vp_p.n5110 16.403
R5318 vp_p.n5099 vp_p.n5096 16.403
R5319 vp_p.n5085 vp_p.n5082 16.403
R5320 vp_p.n5071 vp_p.n5068 16.403
R5321 vp_p.n5057 vp_p.n5054 16.403
R5322 vp_p.n5043 vp_p.n5040 16.403
R5323 vp_p.n5029 vp_p.n5026 16.403
R5324 vp_p.n5015 vp_p.n5012 16.403
R5325 vp_p.n5001 vp_p.n4998 16.403
R5326 vp_p.n4987 vp_p.n4984 16.403
R5327 vp_p.n4973 vp_p.n4970 16.403
R5328 vp_p.n4959 vp_p.n4956 16.403
R5329 vp_p.n4945 vp_p.n4942 16.403
R5330 vp_p.n4931 vp_p.n4928 16.403
R5331 vp_p.n4917 vp_p.n4914 16.403
R5332 vp_p.n4903 vp_p.n4900 16.403
R5333 vp_p.n4889 vp_p.n4886 16.403
R5334 vp_p.n4875 vp_p.n4872 16.403
R5335 vp_p.n4861 vp_p.n4858 16.403
R5336 vp_p.n4847 vp_p.n4844 16.403
R5337 vp_p.n4833 vp_p.n4830 16.403
R5338 vp_p.n4819 vp_p.n4816 16.403
R5339 vp_p.n4805 vp_p.n4802 16.403
R5340 vp_p.n4791 vp_p.n4788 16.403
R5341 vp_p.n4777 vp_p.n4774 16.403
R5342 vp_p.n4763 vp_p.n4760 16.403
R5343 vp_p.n4749 vp_p.n4746 16.403
R5344 vp_p.n24445 vp_p.n24442 16.403
R5345 vp_p.n24431 vp_p.n24428 16.403
R5346 vp_p.n24417 vp_p.n24414 16.403
R5347 vp_p.n24403 vp_p.n24400 16.403
R5348 vp_p.n24389 vp_p.n24386 16.403
R5349 vp_p.n24375 vp_p.n24372 16.403
R5350 vp_p.n24361 vp_p.n24358 16.403
R5351 vp_p.n24347 vp_p.n24344 16.403
R5352 vp_p.n24333 vp_p.n24330 16.403
R5353 vp_p.n24319 vp_p.n24316 16.403
R5354 vp_p.n24305 vp_p.n24302 16.403
R5355 vp_p.n24291 vp_p.n24288 16.403
R5356 vp_p.n24277 vp_p.n24274 16.403
R5357 vp_p.n24263 vp_p.n24260 16.403
R5358 vp_p.n24249 vp_p.n24246 16.403
R5359 vp_p.n24235 vp_p.n24232 16.403
R5360 vp_p.n24221 vp_p.n24218 16.403
R5361 vp_p.n24207 vp_p.n24204 16.403
R5362 vp_p.n24193 vp_p.n24190 16.403
R5363 vp_p.n24179 vp_p.n24176 16.403
R5364 vp_p.n24165 vp_p.n24162 16.403
R5365 vp_p.n24151 vp_p.n24148 16.403
R5366 vp_p.n24137 vp_p.n24134 16.403
R5367 vp_p.n24123 vp_p.n24120 16.403
R5368 vp_p.n24109 vp_p.n24106 16.403
R5369 vp_p.n24095 vp_p.n24092 16.403
R5370 vp_p.n24081 vp_p.n24078 16.403
R5371 vp_p.n24067 vp_p.n24064 16.403
R5372 vp_p.n24053 vp_p.n24050 16.403
R5373 vp_p.n24039 vp_p.n24036 16.403
R5374 vp_p.n24025 vp_p.n24022 16.403
R5375 vp_p.n24011 vp_p.n24008 16.403
R5376 vp_p.n23997 vp_p.n23994 16.403
R5377 vp_p.n23983 vp_p.n23980 16.403
R5378 vp_p.n23969 vp_p.n23966 16.403
R5379 vp_p.n23955 vp_p.n23952 16.403
R5380 vp_p.n23941 vp_p.n23938 16.403
R5381 vp_p.n23927 vp_p.n23924 16.403
R5382 vp_p.n23913 vp_p.n23910 16.403
R5383 vp_p.n23899 vp_p.n23896 16.403
R5384 vp_p.n23885 vp_p.n23882 16.403
R5385 vp_p.n23871 vp_p.n23868 16.403
R5386 vp_p.n23857 vp_p.n23854 16.403
R5387 vp_p.n23843 vp_p.n23840 16.403
R5388 vp_p.n23829 vp_p.n23826 16.403
R5389 vp_p.n23815 vp_p.n23812 16.403
R5390 vp_p.n23801 vp_p.n23798 16.403
R5391 vp_p.n23787 vp_p.n23784 16.403
R5392 vp_p.n23773 vp_p.n23770 16.403
R5393 vp_p.n23759 vp_p.n23756 16.403
R5394 vp_p.n23745 vp_p.n23742 16.403
R5395 vp_p.n23731 vp_p.n23728 16.403
R5396 vp_p.n23717 vp_p.n23714 16.403
R5397 vp_p.n23703 vp_p.n23700 16.403
R5398 vp_p.n23689 vp_p.n23686 16.403
R5399 vp_p.n23675 vp_p.n23672 16.403
R5400 vp_p.n23661 vp_p.n23658 16.403
R5401 vp_p.n23647 vp_p.n23644 16.403
R5402 vp_p.n23633 vp_p.n23630 16.403
R5403 vp_p.n23619 vp_p.n23616 16.403
R5404 vp_p.n23605 vp_p.n23602 16.403
R5405 vp_p.n23591 vp_p.n23588 16.403
R5406 vp_p.n23577 vp_p.n23574 16.403
R5407 vp_p.n23563 vp_p.n23560 16.403
R5408 vp_p.n23549 vp_p.n23546 16.403
R5409 vp_p.n23535 vp_p.n23532 16.403
R5410 vp_p.n23521 vp_p.n23518 16.403
R5411 vp_p.n23507 vp_p.n23504 16.403
R5412 vp_p.n23493 vp_p.n23490 16.403
R5413 vp_p.n23479 vp_p.n23476 16.403
R5414 vp_p.n23465 vp_p.n23462 16.403
R5415 vp_p.n23451 vp_p.n23448 16.403
R5416 vp_p.n7180 vp_p.n7177 16.403
R5417 vp_p.n7166 vp_p.n7163 16.403
R5418 vp_p.n7152 vp_p.n7149 16.403
R5419 vp_p.n7138 vp_p.n7135 16.403
R5420 vp_p.n7124 vp_p.n7121 16.403
R5421 vp_p.n7110 vp_p.n7107 16.403
R5422 vp_p.n7096 vp_p.n7093 16.403
R5423 vp_p.n7082 vp_p.n7079 16.403
R5424 vp_p.n7068 vp_p.n7065 16.403
R5425 vp_p.n7054 vp_p.n7051 16.403
R5426 vp_p.n7040 vp_p.n7037 16.403
R5427 vp_p.n7026 vp_p.n7023 16.403
R5428 vp_p.n7012 vp_p.n7009 16.403
R5429 vp_p.n6998 vp_p.n6995 16.403
R5430 vp_p.n6984 vp_p.n6981 16.403
R5431 vp_p.n6970 vp_p.n6967 16.403
R5432 vp_p.n6956 vp_p.n6953 16.403
R5433 vp_p.n6942 vp_p.n6939 16.403
R5434 vp_p.n6928 vp_p.n6925 16.403
R5435 vp_p.n6914 vp_p.n6911 16.403
R5436 vp_p.n6900 vp_p.n6897 16.403
R5437 vp_p.n6886 vp_p.n6883 16.403
R5438 vp_p.n6872 vp_p.n6869 16.403
R5439 vp_p.n6858 vp_p.n6855 16.403
R5440 vp_p.n6844 vp_p.n6841 16.403
R5441 vp_p.n6830 vp_p.n6827 16.403
R5442 vp_p.n6816 vp_p.n6813 16.403
R5443 vp_p.n6802 vp_p.n6799 16.403
R5444 vp_p.n6788 vp_p.n6785 16.403
R5445 vp_p.n6774 vp_p.n6771 16.403
R5446 vp_p.n6760 vp_p.n6757 16.403
R5447 vp_p.n6746 vp_p.n6743 16.403
R5448 vp_p.n6732 vp_p.n6729 16.403
R5449 vp_p.n6718 vp_p.n6715 16.403
R5450 vp_p.n6704 vp_p.n6701 16.403
R5451 vp_p.n6690 vp_p.n6687 16.403
R5452 vp_p.n6676 vp_p.n6673 16.403
R5453 vp_p.n6662 vp_p.n6659 16.403
R5454 vp_p.n6648 vp_p.n6645 16.403
R5455 vp_p.n6634 vp_p.n6631 16.403
R5456 vp_p.n6620 vp_p.n6617 16.403
R5457 vp_p.n6606 vp_p.n6603 16.403
R5458 vp_p.n6592 vp_p.n6589 16.403
R5459 vp_p.n6578 vp_p.n6575 16.403
R5460 vp_p.n6564 vp_p.n6561 16.403
R5461 vp_p.n6550 vp_p.n6547 16.403
R5462 vp_p.n6536 vp_p.n6533 16.403
R5463 vp_p.n6522 vp_p.n6519 16.403
R5464 vp_p.n6508 vp_p.n6505 16.403
R5465 vp_p.n6494 vp_p.n6491 16.403
R5466 vp_p.n6480 vp_p.n6477 16.403
R5467 vp_p.n6466 vp_p.n6463 16.403
R5468 vp_p.n6452 vp_p.n6449 16.403
R5469 vp_p.n6438 vp_p.n6435 16.403
R5470 vp_p.n6424 vp_p.n6421 16.403
R5471 vp_p.n6410 vp_p.n6407 16.403
R5472 vp_p.n6396 vp_p.n6393 16.403
R5473 vp_p.n6382 vp_p.n6379 16.403
R5474 vp_p.n6368 vp_p.n6365 16.403
R5475 vp_p.n6354 vp_p.n6351 16.403
R5476 vp_p.n6340 vp_p.n6337 16.403
R5477 vp_p.n6326 vp_p.n6323 16.403
R5478 vp_p.n6312 vp_p.n6309 16.403
R5479 vp_p.n6298 vp_p.n6295 16.403
R5480 vp_p.n6284 vp_p.n6281 16.403
R5481 vp_p.n6270 vp_p.n6267 16.403
R5482 vp_p.n6256 vp_p.n6253 16.403
R5483 vp_p.n6242 vp_p.n6239 16.403
R5484 vp_p.n6228 vp_p.n6225 16.403
R5485 vp_p.n6214 vp_p.n6211 16.403
R5486 vp_p.n6200 vp_p.n6197 16.403
R5487 vp_p.n6186 vp_p.n6183 16.403
R5488 vp_p.n6172 vp_p.n6169 16.403
R5489 vp_p.n25881 vp_p.n25878 16.403
R5490 vp_p.n25867 vp_p.n25864 16.403
R5491 vp_p.n25853 vp_p.n25850 16.403
R5492 vp_p.n25839 vp_p.n25836 16.403
R5493 vp_p.n25825 vp_p.n25822 16.403
R5494 vp_p.n25811 vp_p.n25808 16.403
R5495 vp_p.n25797 vp_p.n25794 16.403
R5496 vp_p.n25783 vp_p.n25780 16.403
R5497 vp_p.n25769 vp_p.n25766 16.403
R5498 vp_p.n25755 vp_p.n25752 16.403
R5499 vp_p.n25741 vp_p.n25738 16.403
R5500 vp_p.n25727 vp_p.n25724 16.403
R5501 vp_p.n25713 vp_p.n25710 16.403
R5502 vp_p.n25699 vp_p.n25696 16.403
R5503 vp_p.n25685 vp_p.n25682 16.403
R5504 vp_p.n25671 vp_p.n25668 16.403
R5505 vp_p.n25657 vp_p.n25654 16.403
R5506 vp_p.n25643 vp_p.n25640 16.403
R5507 vp_p.n25629 vp_p.n25626 16.403
R5508 vp_p.n25615 vp_p.n25612 16.403
R5509 vp_p.n25601 vp_p.n25598 16.403
R5510 vp_p.n25587 vp_p.n25584 16.403
R5511 vp_p.n25573 vp_p.n25570 16.403
R5512 vp_p.n25559 vp_p.n25556 16.403
R5513 vp_p.n25545 vp_p.n25542 16.403
R5514 vp_p.n25531 vp_p.n25528 16.403
R5515 vp_p.n25517 vp_p.n25514 16.403
R5516 vp_p.n25503 vp_p.n25500 16.403
R5517 vp_p.n25489 vp_p.n25486 16.403
R5518 vp_p.n25475 vp_p.n25472 16.403
R5519 vp_p.n25461 vp_p.n25458 16.403
R5520 vp_p.n25447 vp_p.n25444 16.403
R5521 vp_p.n25433 vp_p.n25430 16.403
R5522 vp_p.n25419 vp_p.n25416 16.403
R5523 vp_p.n25405 vp_p.n25402 16.403
R5524 vp_p.n25391 vp_p.n25388 16.403
R5525 vp_p.n25377 vp_p.n25374 16.403
R5526 vp_p.n25363 vp_p.n25360 16.403
R5527 vp_p.n25349 vp_p.n25346 16.403
R5528 vp_p.n25335 vp_p.n25332 16.403
R5529 vp_p.n25321 vp_p.n25318 16.403
R5530 vp_p.n25307 vp_p.n25304 16.403
R5531 vp_p.n25293 vp_p.n25290 16.403
R5532 vp_p.n25279 vp_p.n25276 16.403
R5533 vp_p.n25265 vp_p.n25262 16.403
R5534 vp_p.n25251 vp_p.n25248 16.403
R5535 vp_p.n25237 vp_p.n25234 16.403
R5536 vp_p.n25223 vp_p.n25220 16.403
R5537 vp_p.n25209 vp_p.n25206 16.403
R5538 vp_p.n25195 vp_p.n25192 16.403
R5539 vp_p.n25181 vp_p.n25178 16.403
R5540 vp_p.n25167 vp_p.n25164 16.403
R5541 vp_p.n25153 vp_p.n25150 16.403
R5542 vp_p.n25139 vp_p.n25136 16.403
R5543 vp_p.n25125 vp_p.n25122 16.403
R5544 vp_p.n25111 vp_p.n25108 16.403
R5545 vp_p.n25097 vp_p.n25094 16.403
R5546 vp_p.n25083 vp_p.n25080 16.403
R5547 vp_p.n25069 vp_p.n25066 16.403
R5548 vp_p.n25055 vp_p.n25052 16.403
R5549 vp_p.n25041 vp_p.n25038 16.403
R5550 vp_p.n25027 vp_p.n25024 16.403
R5551 vp_p.n25013 vp_p.n25010 16.403
R5552 vp_p.n24999 vp_p.n24996 16.403
R5553 vp_p.n24985 vp_p.n24982 16.403
R5554 vp_p.n24971 vp_p.n24968 16.403
R5555 vp_p.n24957 vp_p.n24954 16.403
R5556 vp_p.n24943 vp_p.n24940 16.403
R5557 vp_p.n24929 vp_p.n24926 16.403
R5558 vp_p.n24915 vp_p.n24912 16.403
R5559 vp_p.n24901 vp_p.n24898 16.403
R5560 vp_p.n24887 vp_p.n24884 16.403
R5561 vp_p.n24873 vp_p.n24870 16.403
R5562 vp_p.n7594 vp_p.n7591 16.403
R5563 vp_p.n7608 vp_p.n7605 16.403
R5564 vp_p.n7622 vp_p.n7619 16.403
R5565 vp_p.n7636 vp_p.n7633 16.403
R5566 vp_p.n7650 vp_p.n7647 16.403
R5567 vp_p.n7664 vp_p.n7661 16.403
R5568 vp_p.n7678 vp_p.n7675 16.403
R5569 vp_p.n7692 vp_p.n7689 16.403
R5570 vp_p.n7706 vp_p.n7703 16.403
R5571 vp_p.n7720 vp_p.n7717 16.403
R5572 vp_p.n7734 vp_p.n7731 16.403
R5573 vp_p.n7748 vp_p.n7745 16.403
R5574 vp_p.n7762 vp_p.n7759 16.403
R5575 vp_p.n7776 vp_p.n7773 16.403
R5576 vp_p.n7790 vp_p.n7787 16.403
R5577 vp_p.n7804 vp_p.n7801 16.403
R5578 vp_p.n7818 vp_p.n7815 16.403
R5579 vp_p.n7832 vp_p.n7829 16.403
R5580 vp_p.n7846 vp_p.n7843 16.403
R5581 vp_p.n7860 vp_p.n7857 16.403
R5582 vp_p.n7874 vp_p.n7871 16.403
R5583 vp_p.n7888 vp_p.n7885 16.403
R5584 vp_p.n7902 vp_p.n7899 16.403
R5585 vp_p.n7916 vp_p.n7913 16.403
R5586 vp_p.n7930 vp_p.n7927 16.403
R5587 vp_p.n7944 vp_p.n7941 16.403
R5588 vp_p.n7958 vp_p.n7955 16.403
R5589 vp_p.n7972 vp_p.n7969 16.403
R5590 vp_p.n7986 vp_p.n7983 16.403
R5591 vp_p.n8000 vp_p.n7997 16.403
R5592 vp_p.n8014 vp_p.n8011 16.403
R5593 vp_p.n8028 vp_p.n8025 16.403
R5594 vp_p.n8042 vp_p.n8039 16.403
R5595 vp_p.n8056 vp_p.n8053 16.403
R5596 vp_p.n8070 vp_p.n8067 16.403
R5597 vp_p.n8084 vp_p.n8081 16.403
R5598 vp_p.n8098 vp_p.n8095 16.403
R5599 vp_p.n8112 vp_p.n8109 16.403
R5600 vp_p.n8126 vp_p.n8123 16.403
R5601 vp_p.n8140 vp_p.n8137 16.403
R5602 vp_p.n8154 vp_p.n8151 16.403
R5603 vp_p.n8168 vp_p.n8165 16.403
R5604 vp_p.n8182 vp_p.n8179 16.403
R5605 vp_p.n8196 vp_p.n8193 16.403
R5606 vp_p.n8210 vp_p.n8207 16.403
R5607 vp_p.n8224 vp_p.n8221 16.403
R5608 vp_p.n8238 vp_p.n8235 16.403
R5609 vp_p.n8252 vp_p.n8249 16.403
R5610 vp_p.n8266 vp_p.n8263 16.403
R5611 vp_p.n8280 vp_p.n8277 16.403
R5612 vp_p.n8294 vp_p.n8291 16.403
R5613 vp_p.n8308 vp_p.n8305 16.403
R5614 vp_p.n8322 vp_p.n8319 16.403
R5615 vp_p.n8336 vp_p.n8333 16.403
R5616 vp_p.n8350 vp_p.n8347 16.403
R5617 vp_p.n8364 vp_p.n8361 16.403
R5618 vp_p.n8378 vp_p.n8375 16.403
R5619 vp_p.n8392 vp_p.n8389 16.403
R5620 vp_p.n8406 vp_p.n8403 16.403
R5621 vp_p.n8420 vp_p.n8417 16.403
R5622 vp_p.n8434 vp_p.n8431 16.403
R5623 vp_p.n8448 vp_p.n8445 16.403
R5624 vp_p.n8462 vp_p.n8459 16.403
R5625 vp_p.n8476 vp_p.n8473 16.403
R5626 vp_p.n8490 vp_p.n8487 16.403
R5627 vp_p.n8504 vp_p.n8501 16.403
R5628 vp_p.n8518 vp_p.n8515 16.403
R5629 vp_p.n8532 vp_p.n8529 16.403
R5630 vp_p.n8546 vp_p.n8543 16.403
R5631 vp_p.n8560 vp_p.n8557 16.403
R5632 vp_p.n8574 vp_p.n8571 16.403
R5633 vp_p.n8588 vp_p.n8585 16.403
R5634 vp_p.n8602 vp_p.n8599 16.403
R5635 vp_p.n8616 vp_p.n8613 16.403
R5636 vp_p.n26298 vp_p.n26295 16.403
R5637 vp_p.n26312 vp_p.n26309 16.403
R5638 vp_p.n26326 vp_p.n26323 16.403
R5639 vp_p.n26340 vp_p.n26337 16.403
R5640 vp_p.n26354 vp_p.n26351 16.403
R5641 vp_p.n26368 vp_p.n26365 16.403
R5642 vp_p.n26382 vp_p.n26379 16.403
R5643 vp_p.n26396 vp_p.n26393 16.403
R5644 vp_p.n26410 vp_p.n26407 16.403
R5645 vp_p.n26424 vp_p.n26421 16.403
R5646 vp_p.n26438 vp_p.n26435 16.403
R5647 vp_p.n26452 vp_p.n26449 16.403
R5648 vp_p.n26466 vp_p.n26463 16.403
R5649 vp_p.n26480 vp_p.n26477 16.403
R5650 vp_p.n26494 vp_p.n26491 16.403
R5651 vp_p.n26508 vp_p.n26505 16.403
R5652 vp_p.n26522 vp_p.n26519 16.403
R5653 vp_p.n26536 vp_p.n26533 16.403
R5654 vp_p.n26550 vp_p.n26547 16.403
R5655 vp_p.n26564 vp_p.n26561 16.403
R5656 vp_p.n26578 vp_p.n26575 16.403
R5657 vp_p.n26592 vp_p.n26589 16.403
R5658 vp_p.n26606 vp_p.n26603 16.403
R5659 vp_p.n26620 vp_p.n26617 16.403
R5660 vp_p.n26634 vp_p.n26631 16.403
R5661 vp_p.n26648 vp_p.n26645 16.403
R5662 vp_p.n26662 vp_p.n26659 16.403
R5663 vp_p.n26676 vp_p.n26673 16.403
R5664 vp_p.n26690 vp_p.n26687 16.403
R5665 vp_p.n26704 vp_p.n26701 16.403
R5666 vp_p.n26718 vp_p.n26715 16.403
R5667 vp_p.n26732 vp_p.n26729 16.403
R5668 vp_p.n26746 vp_p.n26743 16.403
R5669 vp_p.n26760 vp_p.n26757 16.403
R5670 vp_p.n26774 vp_p.n26771 16.403
R5671 vp_p.n26788 vp_p.n26785 16.403
R5672 vp_p.n26802 vp_p.n26799 16.403
R5673 vp_p.n26816 vp_p.n26813 16.403
R5674 vp_p.n26830 vp_p.n26827 16.403
R5675 vp_p.n26844 vp_p.n26841 16.403
R5676 vp_p.n26858 vp_p.n26855 16.403
R5677 vp_p.n26872 vp_p.n26869 16.403
R5678 vp_p.n26886 vp_p.n26883 16.403
R5679 vp_p.n26900 vp_p.n26897 16.403
R5680 vp_p.n26914 vp_p.n26911 16.403
R5681 vp_p.n26928 vp_p.n26925 16.403
R5682 vp_p.n26942 vp_p.n26939 16.403
R5683 vp_p.n26956 vp_p.n26953 16.403
R5684 vp_p.n26970 vp_p.n26967 16.403
R5685 vp_p.n26984 vp_p.n26981 16.403
R5686 vp_p.n26998 vp_p.n26995 16.403
R5687 vp_p.n27012 vp_p.n27009 16.403
R5688 vp_p.n27026 vp_p.n27023 16.403
R5689 vp_p.n27040 vp_p.n27037 16.403
R5690 vp_p.n27054 vp_p.n27051 16.403
R5691 vp_p.n27068 vp_p.n27065 16.403
R5692 vp_p.n27082 vp_p.n27079 16.403
R5693 vp_p.n27096 vp_p.n27093 16.403
R5694 vp_p.n27110 vp_p.n27107 16.403
R5695 vp_p.n27124 vp_p.n27121 16.403
R5696 vp_p.n27138 vp_p.n27135 16.403
R5697 vp_p.n27152 vp_p.n27149 16.403
R5698 vp_p.n27166 vp_p.n27163 16.403
R5699 vp_p.n27180 vp_p.n27177 16.403
R5700 vp_p.n27194 vp_p.n27191 16.403
R5701 vp_p.n27208 vp_p.n27205 16.403
R5702 vp_p.n27222 vp_p.n27219 16.403
R5703 vp_p.n27236 vp_p.n27233 16.403
R5704 vp_p.n27250 vp_p.n27247 16.403
R5705 vp_p.n27264 vp_p.n27261 16.403
R5706 vp_p.n27278 vp_p.n27275 16.403
R5707 vp_p.n27292 vp_p.n27289 16.403
R5708 vp_p.n27306 vp_p.n27303 16.403
R5709 vp_p.n27320 vp_p.n27317 16.403
R5710 vp_p.n26284 vp_p.n26281 16.402
R5711 vp_p.n13182 vp_p.n13181 16.399
R5712 vp_p.n13187 vp_p.n13186 16.399
R5713 vp_p.n13192 vp_p.n13191 16.399
R5714 vp_p.n13197 vp_p.n13196 16.399
R5715 vp_p.n13202 vp_p.n13201 16.399
R5716 vp_p.n13207 vp_p.n13206 16.399
R5717 vp_p.n13212 vp_p.n13211 16.399
R5718 vp_p.n13217 vp_p.n13216 16.399
R5719 vp_p.n13222 vp_p.n13221 16.399
R5720 vp_p.n13227 vp_p.n13226 16.399
R5721 vp_p.n13232 vp_p.n13231 16.399
R5722 vp_p.n13237 vp_p.n13236 16.399
R5723 vp_p.n13242 vp_p.n13241 16.399
R5724 vp_p.n13247 vp_p.n13246 16.399
R5725 vp_p.n13252 vp_p.n13251 16.399
R5726 vp_p.n13257 vp_p.n13256 16.399
R5727 vp_p.n13262 vp_p.n13261 16.399
R5728 vp_p.n13267 vp_p.n13266 16.399
R5729 vp_p.n13272 vp_p.n13271 16.399
R5730 vp_p.n13277 vp_p.n13276 16.399
R5731 vp_p.n13282 vp_p.n13281 16.399
R5732 vp_p.n13287 vp_p.n13286 16.399
R5733 vp_p.n13292 vp_p.n13291 16.399
R5734 vp_p.n13297 vp_p.n13296 16.399
R5735 vp_p.n13302 vp_p.n13301 16.399
R5736 vp_p.n13307 vp_p.n13306 16.399
R5737 vp_p.n13312 vp_p.n13311 16.399
R5738 vp_p.n13317 vp_p.n13316 16.399
R5739 vp_p.n13322 vp_p.n13321 16.399
R5740 vp_p.n13327 vp_p.n13326 16.399
R5741 vp_p.n13332 vp_p.n13331 16.399
R5742 vp_p.n13337 vp_p.n13336 16.399
R5743 vp_p.n13342 vp_p.n13341 16.399
R5744 vp_p.n13347 vp_p.n13346 16.399
R5745 vp_p.n13352 vp_p.n13351 16.399
R5746 vp_p.n13357 vp_p.n13356 16.399
R5747 vp_p.n13362 vp_p.n13361 16.399
R5748 vp_p.n13367 vp_p.n13366 16.399
R5749 vp_p.n13372 vp_p.n13371 16.399
R5750 vp_p.n13377 vp_p.n13376 16.399
R5751 vp_p.n13382 vp_p.n13381 16.399
R5752 vp_p.n13387 vp_p.n13386 16.399
R5753 vp_p.n13392 vp_p.n13391 16.399
R5754 vp_p.n13397 vp_p.n13396 16.399
R5755 vp_p.n13402 vp_p.n13401 16.399
R5756 vp_p.n13407 vp_p.n13406 16.399
R5757 vp_p.n13412 vp_p.n13411 16.399
R5758 vp_p.n13417 vp_p.n13416 16.399
R5759 vp_p.n13422 vp_p.n13421 16.399
R5760 vp_p.n13427 vp_p.n13426 16.399
R5761 vp_p.n13432 vp_p.n13431 16.399
R5762 vp_p.n13437 vp_p.n13436 16.399
R5763 vp_p.n13442 vp_p.n13441 16.399
R5764 vp_p.n13447 vp_p.n13446 16.399
R5765 vp_p.n13452 vp_p.n13451 16.399
R5766 vp_p.n13457 vp_p.n13456 16.399
R5767 vp_p.n13462 vp_p.n13461 16.399
R5768 vp_p.n13467 vp_p.n13466 16.399
R5769 vp_p.n13472 vp_p.n13471 16.399
R5770 vp_p.n13477 vp_p.n13476 16.399
R5771 vp_p.n13482 vp_p.n13481 16.399
R5772 vp_p.n13487 vp_p.n13486 16.399
R5773 vp_p.n13492 vp_p.n13491 16.399
R5774 vp_p.n13497 vp_p.n13496 16.399
R5775 vp_p.n13502 vp_p.n13501 16.399
R5776 vp_p.n13507 vp_p.n13506 16.399
R5777 vp_p.n13512 vp_p.n13511 16.399
R5778 vp_p.n13517 vp_p.n13516 16.399
R5779 vp_p.n13522 vp_p.n13521 16.399
R5780 vp_p.n13527 vp_p.n13526 16.399
R5781 vp_p.n13532 vp_p.n13531 16.399
R5782 vp_p.n13537 vp_p.n13536 16.399
R5783 vp_p.n13542 vp_p.n13541 16.399
R5784 vp_p.n13547 vp_p.n13546 16.399
R5785 vp_p.n13552 vp_p.n13551 16.399
R5786 vp_p.n13557 vp_p.n13556 16.399
R5787 vp_p.n13562 vp_p.n13561 16.399
R5788 vp_p.n13567 vp_p.n13566 16.399
R5789 vp_p.n13572 vp_p.n13571 16.399
R5790 vp_p.n13577 vp_p.n13576 16.399
R5791 vp_p.n13582 vp_p.n13581 16.399
R5792 vp_p.n13587 vp_p.n13586 16.399
R5793 vp_p.n13592 vp_p.n13591 16.399
R5794 vp_p.n13597 vp_p.n13596 16.399
R5795 vp_p.n13602 vp_p.n13601 16.399
R5796 vp_p.n13607 vp_p.n13606 16.399
R5797 vp_p.n13612 vp_p.n13611 16.399
R5798 vp_p.n13617 vp_p.n13616 16.399
R5799 vp_p.n13622 vp_p.n13621 16.399
R5800 vp_p.n13627 vp_p.n13626 16.399
R5801 vp_p.n13632 vp_p.n13631 16.399
R5802 vp_p.n13637 vp_p.n13636 16.399
R5803 vp_p.n13642 vp_p.n13641 16.399
R5804 vp_p.n13647 vp_p.n13646 16.399
R5805 vp_p.n13652 vp_p.n13651 16.399
R5806 vp_p.n13657 vp_p.n13656 16.399
R5807 vp_p.n13662 vp_p.n13661 16.399
R5808 vp_p.n13667 vp_p.n13666 16.399
R5809 vp_p.n13672 vp_p.n13671 16.399
R5810 vp_p.n13677 vp_p.n13676 16.399
R5811 vp_p.n13682 vp_p.n13681 16.399
R5812 vp_p.n13687 vp_p.n13686 16.399
R5813 vp_p.n13692 vp_p.n13691 16.399
R5814 vp_p.n13697 vp_p.n13696 16.399
R5815 vp_p.n13702 vp_p.n13701 16.399
R5816 vp_p.n13707 vp_p.n13706 16.399
R5817 vp_p.n13712 vp_p.n13711 16.399
R5818 vp_p.n13717 vp_p.n13716 16.399
R5819 vp_p.n13722 vp_p.n13721 16.399
R5820 vp_p.n13727 vp_p.n13726 16.399
R5821 vp_p.n13732 vp_p.n13731 16.399
R5822 vp_p.n13737 vp_p.n13736 16.399
R5823 vp_p.n13742 vp_p.n13741 16.399
R5824 vp_p.n13747 vp_p.n13746 16.399
R5825 vp_p.n13752 vp_p.n13751 16.399
R5826 vp_p.n13757 vp_p.n13756 16.399
R5827 vp_p.n13762 vp_p.n13761 16.399
R5828 vp_p.n13767 vp_p.n13766 16.399
R5829 vp_p.n13772 vp_p.n13771 16.399
R5830 vp_p.n13777 vp_p.n13776 16.399
R5831 vp_p.n13782 vp_p.n13781 16.399
R5832 vp_p.n13787 vp_p.n13786 16.399
R5833 vp_p.n13792 vp_p.n13791 16.399
R5834 vp_p.n13797 vp_p.n13796 16.399
R5835 vp_p.n13802 vp_p.n13801 16.399
R5836 vp_p.n13807 vp_p.n13806 16.399
R5837 vp_p.n13812 vp_p.n13811 16.399
R5838 vp_p.n13817 vp_p.n13816 16.399
R5839 vp_p.n13822 vp_p.n13821 16.399
R5840 vp_p.n13827 vp_p.n13826 16.399
R5841 vp_p.n13832 vp_p.n13831 16.399
R5842 vp_p.n11743 vp_p.n11742 16.399
R5843 vp_p.n11748 vp_p.n11747 16.399
R5844 vp_p.n11753 vp_p.n11752 16.399
R5845 vp_p.n11758 vp_p.n11757 16.399
R5846 vp_p.n11763 vp_p.n11762 16.399
R5847 vp_p.n11768 vp_p.n11767 16.399
R5848 vp_p.n11773 vp_p.n11772 16.399
R5849 vp_p.n11778 vp_p.n11777 16.399
R5850 vp_p.n11783 vp_p.n11782 16.399
R5851 vp_p.n11788 vp_p.n11787 16.399
R5852 vp_p.n11793 vp_p.n11792 16.399
R5853 vp_p.n11798 vp_p.n11797 16.399
R5854 vp_p.n11803 vp_p.n11802 16.399
R5855 vp_p.n11808 vp_p.n11807 16.399
R5856 vp_p.n11813 vp_p.n11812 16.399
R5857 vp_p.n11818 vp_p.n11817 16.399
R5858 vp_p.n11823 vp_p.n11822 16.399
R5859 vp_p.n11828 vp_p.n11827 16.399
R5860 vp_p.n11833 vp_p.n11832 16.399
R5861 vp_p.n11838 vp_p.n11837 16.399
R5862 vp_p.n11843 vp_p.n11842 16.399
R5863 vp_p.n11848 vp_p.n11847 16.399
R5864 vp_p.n11853 vp_p.n11852 16.399
R5865 vp_p.n11858 vp_p.n11857 16.399
R5866 vp_p.n11863 vp_p.n11862 16.399
R5867 vp_p.n11868 vp_p.n11867 16.399
R5868 vp_p.n11873 vp_p.n11872 16.399
R5869 vp_p.n11878 vp_p.n11877 16.399
R5870 vp_p.n11883 vp_p.n11882 16.399
R5871 vp_p.n11888 vp_p.n11887 16.399
R5872 vp_p.n11893 vp_p.n11892 16.399
R5873 vp_p.n11898 vp_p.n11897 16.399
R5874 vp_p.n11903 vp_p.n11902 16.399
R5875 vp_p.n11908 vp_p.n11907 16.399
R5876 vp_p.n11913 vp_p.n11912 16.399
R5877 vp_p.n11918 vp_p.n11917 16.399
R5878 vp_p.n11923 vp_p.n11922 16.399
R5879 vp_p.n11928 vp_p.n11927 16.399
R5880 vp_p.n11933 vp_p.n11932 16.399
R5881 vp_p.n11938 vp_p.n11937 16.399
R5882 vp_p.n11943 vp_p.n11942 16.399
R5883 vp_p.n11948 vp_p.n11947 16.399
R5884 vp_p.n11953 vp_p.n11952 16.399
R5885 vp_p.n11958 vp_p.n11957 16.399
R5886 vp_p.n11963 vp_p.n11962 16.399
R5887 vp_p.n11968 vp_p.n11967 16.399
R5888 vp_p.n11973 vp_p.n11972 16.399
R5889 vp_p.n11978 vp_p.n11977 16.399
R5890 vp_p.n11983 vp_p.n11982 16.399
R5891 vp_p.n11988 vp_p.n11987 16.399
R5892 vp_p.n11993 vp_p.n11992 16.399
R5893 vp_p.n11998 vp_p.n11997 16.399
R5894 vp_p.n12003 vp_p.n12002 16.399
R5895 vp_p.n12008 vp_p.n12007 16.399
R5896 vp_p.n12013 vp_p.n12012 16.399
R5897 vp_p.n12018 vp_p.n12017 16.399
R5898 vp_p.n12023 vp_p.n12022 16.399
R5899 vp_p.n12028 vp_p.n12027 16.399
R5900 vp_p.n12033 vp_p.n12032 16.399
R5901 vp_p.n12038 vp_p.n12037 16.399
R5902 vp_p.n12043 vp_p.n12042 16.399
R5903 vp_p.n12048 vp_p.n12047 16.399
R5904 vp_p.n12053 vp_p.n12052 16.399
R5905 vp_p.n12058 vp_p.n12057 16.399
R5906 vp_p.n12063 vp_p.n12062 16.399
R5907 vp_p.n12068 vp_p.n12067 16.399
R5908 vp_p.n14541 vp_p.n14540 16.399
R5909 vp_p.n14546 vp_p.n14545 16.399
R5910 vp_p.n14551 vp_p.n14550 16.399
R5911 vp_p.n14556 vp_p.n14555 16.399
R5912 vp_p.n14561 vp_p.n14560 16.399
R5913 vp_p.n14566 vp_p.n14565 16.399
R5914 vp_p.n14571 vp_p.n14570 16.399
R5915 vp_p.n14576 vp_p.n14575 16.399
R5916 vp_p.n14581 vp_p.n14580 16.399
R5917 vp_p.n14586 vp_p.n14585 16.399
R5918 vp_p.n14591 vp_p.n14590 16.399
R5919 vp_p.n14596 vp_p.n14595 16.399
R5920 vp_p.n14601 vp_p.n14600 16.399
R5921 vp_p.n14606 vp_p.n14605 16.399
R5922 vp_p.n14611 vp_p.n14610 16.399
R5923 vp_p.n14616 vp_p.n14615 16.399
R5924 vp_p.n14621 vp_p.n14620 16.399
R5925 vp_p.n14626 vp_p.n14625 16.399
R5926 vp_p.n14631 vp_p.n14630 16.399
R5927 vp_p.n14636 vp_p.n14635 16.399
R5928 vp_p.n14641 vp_p.n14640 16.399
R5929 vp_p.n14646 vp_p.n14645 16.399
R5930 vp_p.n14651 vp_p.n14650 16.399
R5931 vp_p.n14656 vp_p.n14655 16.399
R5932 vp_p.n14661 vp_p.n14660 16.399
R5933 vp_p.n14666 vp_p.n14665 16.399
R5934 vp_p.n14671 vp_p.n14670 16.399
R5935 vp_p.n14676 vp_p.n14675 16.399
R5936 vp_p.n14681 vp_p.n14680 16.399
R5937 vp_p.n14686 vp_p.n14685 16.399
R5938 vp_p.n14691 vp_p.n14690 16.399
R5939 vp_p.n14696 vp_p.n14695 16.399
R5940 vp_p.n14701 vp_p.n14700 16.399
R5941 vp_p.n14706 vp_p.n14705 16.399
R5942 vp_p.n14711 vp_p.n14710 16.399
R5943 vp_p.n14716 vp_p.n14715 16.399
R5944 vp_p.n14721 vp_p.n14720 16.399
R5945 vp_p.n14726 vp_p.n14725 16.399
R5946 vp_p.n14731 vp_p.n14730 16.399
R5947 vp_p.n14736 vp_p.n14735 16.399
R5948 vp_p.n14741 vp_p.n14740 16.399
R5949 vp_p.n14746 vp_p.n14745 16.399
R5950 vp_p.n14751 vp_p.n14750 16.399
R5951 vp_p.n14756 vp_p.n14755 16.399
R5952 vp_p.n14761 vp_p.n14760 16.399
R5953 vp_p.n14766 vp_p.n14765 16.399
R5954 vp_p.n14771 vp_p.n14770 16.399
R5955 vp_p.n14776 vp_p.n14775 16.399
R5956 vp_p.n14781 vp_p.n14780 16.399
R5957 vp_p.n14786 vp_p.n14785 16.399
R5958 vp_p.n14791 vp_p.n14790 16.399
R5959 vp_p.n14796 vp_p.n14795 16.399
R5960 vp_p.n14801 vp_p.n14800 16.399
R5961 vp_p.n14806 vp_p.n14805 16.399
R5962 vp_p.n14811 vp_p.n14810 16.399
R5963 vp_p.n14816 vp_p.n14815 16.399
R5964 vp_p.n14821 vp_p.n14820 16.399
R5965 vp_p.n14826 vp_p.n14825 16.399
R5966 vp_p.n14831 vp_p.n14830 16.399
R5967 vp_p.n14836 vp_p.n14835 16.399
R5968 vp_p.n14841 vp_p.n14840 16.399
R5969 vp_p.n14846 vp_p.n14845 16.399
R5970 vp_p.n14851 vp_p.n14850 16.399
R5971 vp_p.n14856 vp_p.n14855 16.399
R5972 vp_p.n14861 vp_p.n14860 16.399
R5973 vp_p.n14866 vp_p.n14865 16.399
R5974 vp_p.n14871 vp_p.n14870 16.399
R5975 vp_p.n10300 vp_p.n10299 16.399
R5976 vp_p.n10305 vp_p.n10304 16.399
R5977 vp_p.n10310 vp_p.n10309 16.399
R5978 vp_p.n10315 vp_p.n10314 16.399
R5979 vp_p.n10320 vp_p.n10319 16.399
R5980 vp_p.n10325 vp_p.n10324 16.399
R5981 vp_p.n10330 vp_p.n10329 16.399
R5982 vp_p.n10335 vp_p.n10334 16.399
R5983 vp_p.n10340 vp_p.n10339 16.399
R5984 vp_p.n10345 vp_p.n10344 16.399
R5985 vp_p.n10350 vp_p.n10349 16.399
R5986 vp_p.n10355 vp_p.n10354 16.399
R5987 vp_p.n10360 vp_p.n10359 16.399
R5988 vp_p.n10365 vp_p.n10364 16.399
R5989 vp_p.n10370 vp_p.n10369 16.399
R5990 vp_p.n10375 vp_p.n10374 16.399
R5991 vp_p.n10380 vp_p.n10379 16.399
R5992 vp_p.n10385 vp_p.n10384 16.399
R5993 vp_p.n10390 vp_p.n10389 16.399
R5994 vp_p.n10395 vp_p.n10394 16.399
R5995 vp_p.n10400 vp_p.n10399 16.399
R5996 vp_p.n10405 vp_p.n10404 16.399
R5997 vp_p.n10410 vp_p.n10409 16.399
R5998 vp_p.n10415 vp_p.n10414 16.399
R5999 vp_p.n10420 vp_p.n10419 16.399
R6000 vp_p.n10425 vp_p.n10424 16.399
R6001 vp_p.n10430 vp_p.n10429 16.399
R6002 vp_p.n10435 vp_p.n10434 16.399
R6003 vp_p.n10440 vp_p.n10439 16.399
R6004 vp_p.n10445 vp_p.n10444 16.399
R6005 vp_p.n10450 vp_p.n10449 16.399
R6006 vp_p.n10455 vp_p.n10454 16.399
R6007 vp_p.n10460 vp_p.n10459 16.399
R6008 vp_p.n10465 vp_p.n10464 16.399
R6009 vp_p.n10470 vp_p.n10469 16.399
R6010 vp_p.n10475 vp_p.n10474 16.399
R6011 vp_p.n10480 vp_p.n10479 16.399
R6012 vp_p.n10485 vp_p.n10484 16.399
R6013 vp_p.n10490 vp_p.n10489 16.399
R6014 vp_p.n10495 vp_p.n10494 16.399
R6015 vp_p.n10500 vp_p.n10499 16.399
R6016 vp_p.n10505 vp_p.n10504 16.399
R6017 vp_p.n10510 vp_p.n10509 16.399
R6018 vp_p.n10515 vp_p.n10514 16.399
R6019 vp_p.n10520 vp_p.n10519 16.399
R6020 vp_p.n10525 vp_p.n10524 16.399
R6021 vp_p.n10530 vp_p.n10529 16.399
R6022 vp_p.n10535 vp_p.n10534 16.399
R6023 vp_p.n10540 vp_p.n10539 16.399
R6024 vp_p.n10545 vp_p.n10544 16.399
R6025 vp_p.n10550 vp_p.n10549 16.399
R6026 vp_p.n10555 vp_p.n10554 16.399
R6027 vp_p.n10560 vp_p.n10559 16.399
R6028 vp_p.n10565 vp_p.n10564 16.399
R6029 vp_p.n10570 vp_p.n10569 16.399
R6030 vp_p.n10575 vp_p.n10574 16.399
R6031 vp_p.n10580 vp_p.n10579 16.399
R6032 vp_p.n10585 vp_p.n10584 16.399
R6033 vp_p.n10590 vp_p.n10589 16.399
R6034 vp_p.n10595 vp_p.n10594 16.399
R6035 vp_p.n10600 vp_p.n10599 16.399
R6036 vp_p.n10605 vp_p.n10604 16.399
R6037 vp_p.n10610 vp_p.n10609 16.399
R6038 vp_p.n10615 vp_p.n10614 16.399
R6039 vp_p.n10620 vp_p.n10619 16.399
R6040 vp_p.n10625 vp_p.n10624 16.399
R6041 vp_p.n10630 vp_p.n10629 16.399
R6042 vp_p.n15964 vp_p.n15963 16.399
R6043 vp_p.n15969 vp_p.n15968 16.399
R6044 vp_p.n15974 vp_p.n15973 16.399
R6045 vp_p.n15979 vp_p.n15978 16.399
R6046 vp_p.n15984 vp_p.n15983 16.399
R6047 vp_p.n15989 vp_p.n15988 16.399
R6048 vp_p.n15994 vp_p.n15993 16.399
R6049 vp_p.n15999 vp_p.n15998 16.399
R6050 vp_p.n16004 vp_p.n16003 16.399
R6051 vp_p.n16009 vp_p.n16008 16.399
R6052 vp_p.n16014 vp_p.n16013 16.399
R6053 vp_p.n16019 vp_p.n16018 16.399
R6054 vp_p.n16024 vp_p.n16023 16.399
R6055 vp_p.n16029 vp_p.n16028 16.399
R6056 vp_p.n16034 vp_p.n16033 16.399
R6057 vp_p.n16039 vp_p.n16038 16.399
R6058 vp_p.n16044 vp_p.n16043 16.399
R6059 vp_p.n16049 vp_p.n16048 16.399
R6060 vp_p.n16054 vp_p.n16053 16.399
R6061 vp_p.n16059 vp_p.n16058 16.399
R6062 vp_p.n16064 vp_p.n16063 16.399
R6063 vp_p.n16069 vp_p.n16068 16.399
R6064 vp_p.n16074 vp_p.n16073 16.399
R6065 vp_p.n16079 vp_p.n16078 16.399
R6066 vp_p.n16084 vp_p.n16083 16.399
R6067 vp_p.n16089 vp_p.n16088 16.399
R6068 vp_p.n16094 vp_p.n16093 16.399
R6069 vp_p.n16099 vp_p.n16098 16.399
R6070 vp_p.n16104 vp_p.n16103 16.399
R6071 vp_p.n16109 vp_p.n16108 16.399
R6072 vp_p.n16114 vp_p.n16113 16.399
R6073 vp_p.n16119 vp_p.n16118 16.399
R6074 vp_p.n16124 vp_p.n16123 16.399
R6075 vp_p.n16129 vp_p.n16128 16.399
R6076 vp_p.n16134 vp_p.n16133 16.399
R6077 vp_p.n16139 vp_p.n16138 16.399
R6078 vp_p.n16144 vp_p.n16143 16.399
R6079 vp_p.n16149 vp_p.n16148 16.399
R6080 vp_p.n16154 vp_p.n16153 16.399
R6081 vp_p.n16159 vp_p.n16158 16.399
R6082 vp_p.n16164 vp_p.n16163 16.399
R6083 vp_p.n16169 vp_p.n16168 16.399
R6084 vp_p.n16174 vp_p.n16173 16.399
R6085 vp_p.n16179 vp_p.n16178 16.399
R6086 vp_p.n16184 vp_p.n16183 16.399
R6087 vp_p.n16189 vp_p.n16188 16.399
R6088 vp_p.n16194 vp_p.n16193 16.399
R6089 vp_p.n16199 vp_p.n16198 16.399
R6090 vp_p.n16204 vp_p.n16203 16.399
R6091 vp_p.n16209 vp_p.n16208 16.399
R6092 vp_p.n16214 vp_p.n16213 16.399
R6093 vp_p.n16219 vp_p.n16218 16.399
R6094 vp_p.n16224 vp_p.n16223 16.399
R6095 vp_p.n16229 vp_p.n16228 16.399
R6096 vp_p.n16234 vp_p.n16233 16.399
R6097 vp_p.n16239 vp_p.n16238 16.399
R6098 vp_p.n16244 vp_p.n16243 16.399
R6099 vp_p.n16249 vp_p.n16248 16.399
R6100 vp_p.n16254 vp_p.n16253 16.399
R6101 vp_p.n16259 vp_p.n16258 16.399
R6102 vp_p.n16264 vp_p.n16263 16.399
R6103 vp_p.n16269 vp_p.n16268 16.399
R6104 vp_p.n16274 vp_p.n16273 16.399
R6105 vp_p.n16279 vp_p.n16278 16.399
R6106 vp_p.n16284 vp_p.n16283 16.399
R6107 vp_p.n16289 vp_p.n16288 16.399
R6108 vp_p.n16294 vp_p.n16293 16.399
R6109 vp_p.n16299 vp_p.n16298 16.399
R6110 vp_p.n8793 vp_p.n8792 16.399
R6111 vp_p.n8798 vp_p.n8797 16.399
R6112 vp_p.n8803 vp_p.n8802 16.399
R6113 vp_p.n8808 vp_p.n8807 16.399
R6114 vp_p.n8813 vp_p.n8812 16.399
R6115 vp_p.n8818 vp_p.n8817 16.399
R6116 vp_p.n8823 vp_p.n8822 16.399
R6117 vp_p.n8828 vp_p.n8827 16.399
R6118 vp_p.n8833 vp_p.n8832 16.399
R6119 vp_p.n8838 vp_p.n8837 16.399
R6120 vp_p.n8843 vp_p.n8842 16.399
R6121 vp_p.n8848 vp_p.n8847 16.399
R6122 vp_p.n8853 vp_p.n8852 16.399
R6123 vp_p.n8858 vp_p.n8857 16.399
R6124 vp_p.n8863 vp_p.n8862 16.399
R6125 vp_p.n8868 vp_p.n8867 16.399
R6126 vp_p.n8873 vp_p.n8872 16.399
R6127 vp_p.n8878 vp_p.n8877 16.399
R6128 vp_p.n8883 vp_p.n8882 16.399
R6129 vp_p.n8888 vp_p.n8887 16.399
R6130 vp_p.n8893 vp_p.n8892 16.399
R6131 vp_p.n8898 vp_p.n8897 16.399
R6132 vp_p.n8903 vp_p.n8902 16.399
R6133 vp_p.n8908 vp_p.n8907 16.399
R6134 vp_p.n8913 vp_p.n8912 16.399
R6135 vp_p.n8918 vp_p.n8917 16.399
R6136 vp_p.n8923 vp_p.n8922 16.399
R6137 vp_p.n8928 vp_p.n8927 16.399
R6138 vp_p.n8933 vp_p.n8932 16.399
R6139 vp_p.n8938 vp_p.n8937 16.399
R6140 vp_p.n8943 vp_p.n8942 16.399
R6141 vp_p.n8948 vp_p.n8947 16.399
R6142 vp_p.n8953 vp_p.n8952 16.399
R6143 vp_p.n8958 vp_p.n8957 16.399
R6144 vp_p.n8963 vp_p.n8962 16.399
R6145 vp_p.n8968 vp_p.n8967 16.399
R6146 vp_p.n8973 vp_p.n8972 16.399
R6147 vp_p.n8978 vp_p.n8977 16.399
R6148 vp_p.n8983 vp_p.n8982 16.399
R6149 vp_p.n8988 vp_p.n8987 16.399
R6150 vp_p.n8993 vp_p.n8992 16.399
R6151 vp_p.n8998 vp_p.n8997 16.399
R6152 vp_p.n9003 vp_p.n9002 16.399
R6153 vp_p.n9008 vp_p.n9007 16.399
R6154 vp_p.n9013 vp_p.n9012 16.399
R6155 vp_p.n9018 vp_p.n9017 16.399
R6156 vp_p.n9023 vp_p.n9022 16.399
R6157 vp_p.n9028 vp_p.n9027 16.399
R6158 vp_p.n9033 vp_p.n9032 16.399
R6159 vp_p.n9038 vp_p.n9037 16.399
R6160 vp_p.n9043 vp_p.n9042 16.399
R6161 vp_p.n9048 vp_p.n9047 16.399
R6162 vp_p.n9053 vp_p.n9052 16.399
R6163 vp_p.n9058 vp_p.n9057 16.399
R6164 vp_p.n9063 vp_p.n9062 16.399
R6165 vp_p.n9068 vp_p.n9067 16.399
R6166 vp_p.n9073 vp_p.n9072 16.399
R6167 vp_p.n9078 vp_p.n9077 16.399
R6168 vp_p.n9083 vp_p.n9082 16.399
R6169 vp_p.n9088 vp_p.n9087 16.399
R6170 vp_p.n9093 vp_p.n9092 16.399
R6171 vp_p.n9098 vp_p.n9097 16.399
R6172 vp_p.n9103 vp_p.n9102 16.399
R6173 vp_p.n9108 vp_p.n9107 16.399
R6174 vp_p.n9113 vp_p.n9112 16.399
R6175 vp_p.n9118 vp_p.n9117 16.399
R6176 vp_p.n9123 vp_p.n9122 16.399
R6177 vp_p.n9128 vp_p.n9127 16.399
R6178 vp_p.n17386 vp_p.n17385 16.399
R6179 vp_p.n17391 vp_p.n17390 16.399
R6180 vp_p.n17396 vp_p.n17395 16.399
R6181 vp_p.n17401 vp_p.n17400 16.399
R6182 vp_p.n17406 vp_p.n17405 16.399
R6183 vp_p.n17411 vp_p.n17410 16.399
R6184 vp_p.n17416 vp_p.n17415 16.399
R6185 vp_p.n17421 vp_p.n17420 16.399
R6186 vp_p.n17426 vp_p.n17425 16.399
R6187 vp_p.n17431 vp_p.n17430 16.399
R6188 vp_p.n17436 vp_p.n17435 16.399
R6189 vp_p.n17441 vp_p.n17440 16.399
R6190 vp_p.n17446 vp_p.n17445 16.399
R6191 vp_p.n17451 vp_p.n17450 16.399
R6192 vp_p.n17456 vp_p.n17455 16.399
R6193 vp_p.n17461 vp_p.n17460 16.399
R6194 vp_p.n17466 vp_p.n17465 16.399
R6195 vp_p.n17471 vp_p.n17470 16.399
R6196 vp_p.n17476 vp_p.n17475 16.399
R6197 vp_p.n17481 vp_p.n17480 16.399
R6198 vp_p.n17486 vp_p.n17485 16.399
R6199 vp_p.n17491 vp_p.n17490 16.399
R6200 vp_p.n17496 vp_p.n17495 16.399
R6201 vp_p.n17501 vp_p.n17500 16.399
R6202 vp_p.n17506 vp_p.n17505 16.399
R6203 vp_p.n17511 vp_p.n17510 16.399
R6204 vp_p.n17516 vp_p.n17515 16.399
R6205 vp_p.n17521 vp_p.n17520 16.399
R6206 vp_p.n17526 vp_p.n17525 16.399
R6207 vp_p.n17531 vp_p.n17530 16.399
R6208 vp_p.n17536 vp_p.n17535 16.399
R6209 vp_p.n17541 vp_p.n17540 16.399
R6210 vp_p.n17546 vp_p.n17545 16.399
R6211 vp_p.n17551 vp_p.n17550 16.399
R6212 vp_p.n17556 vp_p.n17555 16.399
R6213 vp_p.n17561 vp_p.n17560 16.399
R6214 vp_p.n17566 vp_p.n17565 16.399
R6215 vp_p.n17571 vp_p.n17570 16.399
R6216 vp_p.n17576 vp_p.n17575 16.399
R6217 vp_p.n17581 vp_p.n17580 16.399
R6218 vp_p.n17586 vp_p.n17585 16.399
R6219 vp_p.n17591 vp_p.n17590 16.399
R6220 vp_p.n17596 vp_p.n17595 16.399
R6221 vp_p.n17601 vp_p.n17600 16.399
R6222 vp_p.n17606 vp_p.n17605 16.399
R6223 vp_p.n17611 vp_p.n17610 16.399
R6224 vp_p.n17616 vp_p.n17615 16.399
R6225 vp_p.n17621 vp_p.n17620 16.399
R6226 vp_p.n17626 vp_p.n17625 16.399
R6227 vp_p.n17631 vp_p.n17630 16.399
R6228 vp_p.n17636 vp_p.n17635 16.399
R6229 vp_p.n17641 vp_p.n17640 16.399
R6230 vp_p.n17646 vp_p.n17645 16.399
R6231 vp_p.n17651 vp_p.n17650 16.399
R6232 vp_p.n17656 vp_p.n17655 16.399
R6233 vp_p.n17661 vp_p.n17660 16.399
R6234 vp_p.n17666 vp_p.n17665 16.399
R6235 vp_p.n17671 vp_p.n17670 16.399
R6236 vp_p.n17676 vp_p.n17675 16.399
R6237 vp_p.n17681 vp_p.n17680 16.399
R6238 vp_p.n17686 vp_p.n17685 16.399
R6239 vp_p.n17691 vp_p.n17690 16.399
R6240 vp_p.n17696 vp_p.n17695 16.399
R6241 vp_p.n17701 vp_p.n17700 16.399
R6242 vp_p.n17706 vp_p.n17705 16.399
R6243 vp_p.n17711 vp_p.n17710 16.399
R6244 vp_p.n17716 vp_p.n17715 16.399
R6245 vp_p.n17721 vp_p.n17720 16.399
R6246 vp_p.n17726 vp_p.n17725 16.399
R6247 vp_p.n49 vp_p.n48 16.399
R6248 vp_p.n54 vp_p.n53 16.399
R6249 vp_p.n59 vp_p.n58 16.399
R6250 vp_p.n64 vp_p.n63 16.399
R6251 vp_p.n69 vp_p.n68 16.399
R6252 vp_p.n74 vp_p.n73 16.399
R6253 vp_p.n79 vp_p.n78 16.399
R6254 vp_p.n84 vp_p.n83 16.399
R6255 vp_p.n89 vp_p.n88 16.399
R6256 vp_p.n94 vp_p.n93 16.399
R6257 vp_p.n99 vp_p.n98 16.399
R6258 vp_p.n104 vp_p.n103 16.399
R6259 vp_p.n109 vp_p.n108 16.399
R6260 vp_p.n114 vp_p.n113 16.399
R6261 vp_p.n119 vp_p.n118 16.399
R6262 vp_p.n124 vp_p.n123 16.399
R6263 vp_p.n129 vp_p.n128 16.399
R6264 vp_p.n134 vp_p.n133 16.399
R6265 vp_p.n139 vp_p.n138 16.399
R6266 vp_p.n144 vp_p.n143 16.399
R6267 vp_p.n149 vp_p.n148 16.399
R6268 vp_p.n154 vp_p.n153 16.399
R6269 vp_p.n159 vp_p.n158 16.399
R6270 vp_p.n164 vp_p.n163 16.399
R6271 vp_p.n169 vp_p.n168 16.399
R6272 vp_p.n174 vp_p.n173 16.399
R6273 vp_p.n179 vp_p.n178 16.399
R6274 vp_p.n184 vp_p.n183 16.399
R6275 vp_p.n189 vp_p.n188 16.399
R6276 vp_p.n194 vp_p.n193 16.399
R6277 vp_p.n199 vp_p.n198 16.399
R6278 vp_p.n204 vp_p.n203 16.399
R6279 vp_p.n209 vp_p.n208 16.399
R6280 vp_p.n214 vp_p.n213 16.399
R6281 vp_p.n219 vp_p.n218 16.399
R6282 vp_p.n224 vp_p.n223 16.399
R6283 vp_p.n229 vp_p.n228 16.399
R6284 vp_p.n234 vp_p.n233 16.399
R6285 vp_p.n239 vp_p.n238 16.399
R6286 vp_p.n244 vp_p.n243 16.399
R6287 vp_p.n249 vp_p.n248 16.399
R6288 vp_p.n254 vp_p.n253 16.399
R6289 vp_p.n259 vp_p.n258 16.399
R6290 vp_p.n264 vp_p.n263 16.399
R6291 vp_p.n269 vp_p.n268 16.399
R6292 vp_p.n274 vp_p.n273 16.399
R6293 vp_p.n279 vp_p.n278 16.399
R6294 vp_p.n284 vp_p.n283 16.399
R6295 vp_p.n289 vp_p.n288 16.399
R6296 vp_p.n294 vp_p.n293 16.399
R6297 vp_p.n299 vp_p.n298 16.399
R6298 vp_p.n304 vp_p.n303 16.399
R6299 vp_p.n309 vp_p.n308 16.399
R6300 vp_p.n314 vp_p.n313 16.399
R6301 vp_p.n319 vp_p.n318 16.399
R6302 vp_p.n324 vp_p.n323 16.399
R6303 vp_p.n329 vp_p.n328 16.399
R6304 vp_p.n334 vp_p.n333 16.399
R6305 vp_p.n339 vp_p.n338 16.399
R6306 vp_p.n344 vp_p.n343 16.399
R6307 vp_p.n349 vp_p.n348 16.399
R6308 vp_p.n354 vp_p.n353 16.399
R6309 vp_p.n359 vp_p.n358 16.399
R6310 vp_p.n364 vp_p.n363 16.399
R6311 vp_p.n369 vp_p.n368 16.399
R6312 vp_p.n374 vp_p.n373 16.399
R6313 vp_p.n379 vp_p.n378 16.399
R6314 vp_p.n384 vp_p.n383 16.399
R6315 vp_p.n389 vp_p.n388 16.399
R6316 vp_p.n18807 vp_p.n18806 16.399
R6317 vp_p.n18812 vp_p.n18811 16.399
R6318 vp_p.n18817 vp_p.n18816 16.399
R6319 vp_p.n18822 vp_p.n18821 16.399
R6320 vp_p.n18827 vp_p.n18826 16.399
R6321 vp_p.n18832 vp_p.n18831 16.399
R6322 vp_p.n18837 vp_p.n18836 16.399
R6323 vp_p.n18842 vp_p.n18841 16.399
R6324 vp_p.n18847 vp_p.n18846 16.399
R6325 vp_p.n18852 vp_p.n18851 16.399
R6326 vp_p.n18857 vp_p.n18856 16.399
R6327 vp_p.n18862 vp_p.n18861 16.399
R6328 vp_p.n18867 vp_p.n18866 16.399
R6329 vp_p.n18872 vp_p.n18871 16.399
R6330 vp_p.n18877 vp_p.n18876 16.399
R6331 vp_p.n18882 vp_p.n18881 16.399
R6332 vp_p.n18887 vp_p.n18886 16.399
R6333 vp_p.n18892 vp_p.n18891 16.399
R6334 vp_p.n18897 vp_p.n18896 16.399
R6335 vp_p.n18902 vp_p.n18901 16.399
R6336 vp_p.n18907 vp_p.n18906 16.399
R6337 vp_p.n18912 vp_p.n18911 16.399
R6338 vp_p.n18917 vp_p.n18916 16.399
R6339 vp_p.n18922 vp_p.n18921 16.399
R6340 vp_p.n18927 vp_p.n18926 16.399
R6341 vp_p.n18932 vp_p.n18931 16.399
R6342 vp_p.n18937 vp_p.n18936 16.399
R6343 vp_p.n18942 vp_p.n18941 16.399
R6344 vp_p.n18947 vp_p.n18946 16.399
R6345 vp_p.n18952 vp_p.n18951 16.399
R6346 vp_p.n18957 vp_p.n18956 16.399
R6347 vp_p.n18962 vp_p.n18961 16.399
R6348 vp_p.n18967 vp_p.n18966 16.399
R6349 vp_p.n18972 vp_p.n18971 16.399
R6350 vp_p.n18977 vp_p.n18976 16.399
R6351 vp_p.n18982 vp_p.n18981 16.399
R6352 vp_p.n18987 vp_p.n18986 16.399
R6353 vp_p.n18992 vp_p.n18991 16.399
R6354 vp_p.n18997 vp_p.n18996 16.399
R6355 vp_p.n19002 vp_p.n19001 16.399
R6356 vp_p.n19007 vp_p.n19006 16.399
R6357 vp_p.n19012 vp_p.n19011 16.399
R6358 vp_p.n19017 vp_p.n19016 16.399
R6359 vp_p.n19022 vp_p.n19021 16.399
R6360 vp_p.n19027 vp_p.n19026 16.399
R6361 vp_p.n19032 vp_p.n19031 16.399
R6362 vp_p.n19037 vp_p.n19036 16.399
R6363 vp_p.n19042 vp_p.n19041 16.399
R6364 vp_p.n19047 vp_p.n19046 16.399
R6365 vp_p.n19052 vp_p.n19051 16.399
R6366 vp_p.n19057 vp_p.n19056 16.399
R6367 vp_p.n19062 vp_p.n19061 16.399
R6368 vp_p.n19067 vp_p.n19066 16.399
R6369 vp_p.n19072 vp_p.n19071 16.399
R6370 vp_p.n19077 vp_p.n19076 16.399
R6371 vp_p.n19082 vp_p.n19081 16.399
R6372 vp_p.n19087 vp_p.n19086 16.399
R6373 vp_p.n19092 vp_p.n19091 16.399
R6374 vp_p.n19097 vp_p.n19096 16.399
R6375 vp_p.n19102 vp_p.n19101 16.399
R6376 vp_p.n19107 vp_p.n19106 16.399
R6377 vp_p.n19112 vp_p.n19111 16.399
R6378 vp_p.n19117 vp_p.n19116 16.399
R6379 vp_p.n19122 vp_p.n19121 16.399
R6380 vp_p.n19127 vp_p.n19126 16.399
R6381 vp_p.n19132 vp_p.n19131 16.399
R6382 vp_p.n19137 vp_p.n19136 16.399
R6383 vp_p.n19142 vp_p.n19141 16.399
R6384 vp_p.n19147 vp_p.n19146 16.399
R6385 vp_p.n19152 vp_p.n19151 16.399
R6386 vp_p.n1528 vp_p.n1527 16.399
R6387 vp_p.n1533 vp_p.n1532 16.399
R6388 vp_p.n1538 vp_p.n1537 16.399
R6389 vp_p.n1543 vp_p.n1542 16.399
R6390 vp_p.n1548 vp_p.n1547 16.399
R6391 vp_p.n1553 vp_p.n1552 16.399
R6392 vp_p.n1558 vp_p.n1557 16.399
R6393 vp_p.n1563 vp_p.n1562 16.399
R6394 vp_p.n1568 vp_p.n1567 16.399
R6395 vp_p.n1573 vp_p.n1572 16.399
R6396 vp_p.n1578 vp_p.n1577 16.399
R6397 vp_p.n1583 vp_p.n1582 16.399
R6398 vp_p.n1588 vp_p.n1587 16.399
R6399 vp_p.n1593 vp_p.n1592 16.399
R6400 vp_p.n1598 vp_p.n1597 16.399
R6401 vp_p.n1603 vp_p.n1602 16.399
R6402 vp_p.n1608 vp_p.n1607 16.399
R6403 vp_p.n1613 vp_p.n1612 16.399
R6404 vp_p.n1618 vp_p.n1617 16.399
R6405 vp_p.n1623 vp_p.n1622 16.399
R6406 vp_p.n1628 vp_p.n1627 16.399
R6407 vp_p.n1633 vp_p.n1632 16.399
R6408 vp_p.n1638 vp_p.n1637 16.399
R6409 vp_p.n1643 vp_p.n1642 16.399
R6410 vp_p.n1648 vp_p.n1647 16.399
R6411 vp_p.n1653 vp_p.n1652 16.399
R6412 vp_p.n1658 vp_p.n1657 16.399
R6413 vp_p.n1663 vp_p.n1662 16.399
R6414 vp_p.n1668 vp_p.n1667 16.399
R6415 vp_p.n1673 vp_p.n1672 16.399
R6416 vp_p.n1678 vp_p.n1677 16.399
R6417 vp_p.n1683 vp_p.n1682 16.399
R6418 vp_p.n1688 vp_p.n1687 16.399
R6419 vp_p.n1693 vp_p.n1692 16.399
R6420 vp_p.n1698 vp_p.n1697 16.399
R6421 vp_p.n1703 vp_p.n1702 16.399
R6422 vp_p.n1708 vp_p.n1707 16.399
R6423 vp_p.n1713 vp_p.n1712 16.399
R6424 vp_p.n1718 vp_p.n1717 16.399
R6425 vp_p.n1723 vp_p.n1722 16.399
R6426 vp_p.n1728 vp_p.n1727 16.399
R6427 vp_p.n1733 vp_p.n1732 16.399
R6428 vp_p.n1738 vp_p.n1737 16.399
R6429 vp_p.n1743 vp_p.n1742 16.399
R6430 vp_p.n1748 vp_p.n1747 16.399
R6431 vp_p.n1753 vp_p.n1752 16.399
R6432 vp_p.n1758 vp_p.n1757 16.399
R6433 vp_p.n1763 vp_p.n1762 16.399
R6434 vp_p.n1768 vp_p.n1767 16.399
R6435 vp_p.n1773 vp_p.n1772 16.399
R6436 vp_p.n1778 vp_p.n1777 16.399
R6437 vp_p.n1783 vp_p.n1782 16.399
R6438 vp_p.n1788 vp_p.n1787 16.399
R6439 vp_p.n1793 vp_p.n1792 16.399
R6440 vp_p.n1798 vp_p.n1797 16.399
R6441 vp_p.n1803 vp_p.n1802 16.399
R6442 vp_p.n1808 vp_p.n1807 16.399
R6443 vp_p.n1813 vp_p.n1812 16.399
R6444 vp_p.n1818 vp_p.n1817 16.399
R6445 vp_p.n1823 vp_p.n1822 16.399
R6446 vp_p.n1828 vp_p.n1827 16.399
R6447 vp_p.n1833 vp_p.n1832 16.399
R6448 vp_p.n1838 vp_p.n1837 16.399
R6449 vp_p.n1843 vp_p.n1842 16.399
R6450 vp_p.n1848 vp_p.n1847 16.399
R6451 vp_p.n1853 vp_p.n1852 16.399
R6452 vp_p.n1858 vp_p.n1857 16.399
R6453 vp_p.n1863 vp_p.n1862 16.399
R6454 vp_p.n1868 vp_p.n1867 16.399
R6455 vp_p.n1873 vp_p.n1872 16.399
R6456 vp_p.n20227 vp_p.n20226 16.399
R6457 vp_p.n20232 vp_p.n20231 16.399
R6458 vp_p.n20237 vp_p.n20236 16.399
R6459 vp_p.n20242 vp_p.n20241 16.399
R6460 vp_p.n20247 vp_p.n20246 16.399
R6461 vp_p.n20252 vp_p.n20251 16.399
R6462 vp_p.n20257 vp_p.n20256 16.399
R6463 vp_p.n20262 vp_p.n20261 16.399
R6464 vp_p.n20267 vp_p.n20266 16.399
R6465 vp_p.n20272 vp_p.n20271 16.399
R6466 vp_p.n20277 vp_p.n20276 16.399
R6467 vp_p.n20282 vp_p.n20281 16.399
R6468 vp_p.n20287 vp_p.n20286 16.399
R6469 vp_p.n20292 vp_p.n20291 16.399
R6470 vp_p.n20297 vp_p.n20296 16.399
R6471 vp_p.n20302 vp_p.n20301 16.399
R6472 vp_p.n20307 vp_p.n20306 16.399
R6473 vp_p.n20312 vp_p.n20311 16.399
R6474 vp_p.n20317 vp_p.n20316 16.399
R6475 vp_p.n20322 vp_p.n20321 16.399
R6476 vp_p.n20327 vp_p.n20326 16.399
R6477 vp_p.n20332 vp_p.n20331 16.399
R6478 vp_p.n20337 vp_p.n20336 16.399
R6479 vp_p.n20342 vp_p.n20341 16.399
R6480 vp_p.n20347 vp_p.n20346 16.399
R6481 vp_p.n20352 vp_p.n20351 16.399
R6482 vp_p.n20357 vp_p.n20356 16.399
R6483 vp_p.n20362 vp_p.n20361 16.399
R6484 vp_p.n20367 vp_p.n20366 16.399
R6485 vp_p.n20372 vp_p.n20371 16.399
R6486 vp_p.n20377 vp_p.n20376 16.399
R6487 vp_p.n20382 vp_p.n20381 16.399
R6488 vp_p.n20387 vp_p.n20386 16.399
R6489 vp_p.n20392 vp_p.n20391 16.399
R6490 vp_p.n20397 vp_p.n20396 16.399
R6491 vp_p.n20402 vp_p.n20401 16.399
R6492 vp_p.n20407 vp_p.n20406 16.399
R6493 vp_p.n20412 vp_p.n20411 16.399
R6494 vp_p.n20417 vp_p.n20416 16.399
R6495 vp_p.n20422 vp_p.n20421 16.399
R6496 vp_p.n20427 vp_p.n20426 16.399
R6497 vp_p.n20432 vp_p.n20431 16.399
R6498 vp_p.n20437 vp_p.n20436 16.399
R6499 vp_p.n20442 vp_p.n20441 16.399
R6500 vp_p.n20447 vp_p.n20446 16.399
R6501 vp_p.n20452 vp_p.n20451 16.399
R6502 vp_p.n20457 vp_p.n20456 16.399
R6503 vp_p.n20462 vp_p.n20461 16.399
R6504 vp_p.n20467 vp_p.n20466 16.399
R6505 vp_p.n20472 vp_p.n20471 16.399
R6506 vp_p.n20477 vp_p.n20476 16.399
R6507 vp_p.n20482 vp_p.n20481 16.399
R6508 vp_p.n20487 vp_p.n20486 16.399
R6509 vp_p.n20492 vp_p.n20491 16.399
R6510 vp_p.n20497 vp_p.n20496 16.399
R6511 vp_p.n20502 vp_p.n20501 16.399
R6512 vp_p.n20507 vp_p.n20506 16.399
R6513 vp_p.n20512 vp_p.n20511 16.399
R6514 vp_p.n20517 vp_p.n20516 16.399
R6515 vp_p.n20522 vp_p.n20521 16.399
R6516 vp_p.n20527 vp_p.n20526 16.399
R6517 vp_p.n20532 vp_p.n20531 16.399
R6518 vp_p.n20537 vp_p.n20536 16.399
R6519 vp_p.n20542 vp_p.n20541 16.399
R6520 vp_p.n20547 vp_p.n20546 16.399
R6521 vp_p.n20552 vp_p.n20551 16.399
R6522 vp_p.n20557 vp_p.n20556 16.399
R6523 vp_p.n20562 vp_p.n20561 16.399
R6524 vp_p.n20567 vp_p.n20566 16.399
R6525 vp_p.n20572 vp_p.n20571 16.399
R6526 vp_p.n20577 vp_p.n20576 16.399
R6527 vp_p.n2948 vp_p.n2947 16.399
R6528 vp_p.n2953 vp_p.n2952 16.399
R6529 vp_p.n2958 vp_p.n2957 16.399
R6530 vp_p.n2963 vp_p.n2962 16.399
R6531 vp_p.n2968 vp_p.n2967 16.399
R6532 vp_p.n2973 vp_p.n2972 16.399
R6533 vp_p.n2978 vp_p.n2977 16.399
R6534 vp_p.n2983 vp_p.n2982 16.399
R6535 vp_p.n2988 vp_p.n2987 16.399
R6536 vp_p.n2993 vp_p.n2992 16.399
R6537 vp_p.n2998 vp_p.n2997 16.399
R6538 vp_p.n3003 vp_p.n3002 16.399
R6539 vp_p.n3008 vp_p.n3007 16.399
R6540 vp_p.n3013 vp_p.n3012 16.399
R6541 vp_p.n3018 vp_p.n3017 16.399
R6542 vp_p.n3023 vp_p.n3022 16.399
R6543 vp_p.n3028 vp_p.n3027 16.399
R6544 vp_p.n3033 vp_p.n3032 16.399
R6545 vp_p.n3038 vp_p.n3037 16.399
R6546 vp_p.n3043 vp_p.n3042 16.399
R6547 vp_p.n3048 vp_p.n3047 16.399
R6548 vp_p.n3053 vp_p.n3052 16.399
R6549 vp_p.n3058 vp_p.n3057 16.399
R6550 vp_p.n3063 vp_p.n3062 16.399
R6551 vp_p.n3068 vp_p.n3067 16.399
R6552 vp_p.n3073 vp_p.n3072 16.399
R6553 vp_p.n3078 vp_p.n3077 16.399
R6554 vp_p.n3083 vp_p.n3082 16.399
R6555 vp_p.n3088 vp_p.n3087 16.399
R6556 vp_p.n3093 vp_p.n3092 16.399
R6557 vp_p.n3098 vp_p.n3097 16.399
R6558 vp_p.n3103 vp_p.n3102 16.399
R6559 vp_p.n3108 vp_p.n3107 16.399
R6560 vp_p.n3113 vp_p.n3112 16.399
R6561 vp_p.n3118 vp_p.n3117 16.399
R6562 vp_p.n3123 vp_p.n3122 16.399
R6563 vp_p.n3128 vp_p.n3127 16.399
R6564 vp_p.n3133 vp_p.n3132 16.399
R6565 vp_p.n3138 vp_p.n3137 16.399
R6566 vp_p.n3143 vp_p.n3142 16.399
R6567 vp_p.n3148 vp_p.n3147 16.399
R6568 vp_p.n3153 vp_p.n3152 16.399
R6569 vp_p.n3158 vp_p.n3157 16.399
R6570 vp_p.n3163 vp_p.n3162 16.399
R6571 vp_p.n3168 vp_p.n3167 16.399
R6572 vp_p.n3173 vp_p.n3172 16.399
R6573 vp_p.n3178 vp_p.n3177 16.399
R6574 vp_p.n3183 vp_p.n3182 16.399
R6575 vp_p.n3188 vp_p.n3187 16.399
R6576 vp_p.n3193 vp_p.n3192 16.399
R6577 vp_p.n3198 vp_p.n3197 16.399
R6578 vp_p.n3203 vp_p.n3202 16.399
R6579 vp_p.n3208 vp_p.n3207 16.399
R6580 vp_p.n3213 vp_p.n3212 16.399
R6581 vp_p.n3218 vp_p.n3217 16.399
R6582 vp_p.n3223 vp_p.n3222 16.399
R6583 vp_p.n3228 vp_p.n3227 16.399
R6584 vp_p.n3233 vp_p.n3232 16.399
R6585 vp_p.n3238 vp_p.n3237 16.399
R6586 vp_p.n3243 vp_p.n3242 16.399
R6587 vp_p.n3248 vp_p.n3247 16.399
R6588 vp_p.n3253 vp_p.n3252 16.399
R6589 vp_p.n3258 vp_p.n3257 16.399
R6590 vp_p.n3263 vp_p.n3262 16.399
R6591 vp_p.n3268 vp_p.n3267 16.399
R6592 vp_p.n3273 vp_p.n3272 16.399
R6593 vp_p.n3278 vp_p.n3277 16.399
R6594 vp_p.n3283 vp_p.n3282 16.399
R6595 vp_p.n3288 vp_p.n3287 16.399
R6596 vp_p.n3293 vp_p.n3292 16.399
R6597 vp_p.n3298 vp_p.n3297 16.399
R6598 vp_p.n21646 vp_p.n21645 16.399
R6599 vp_p.n21651 vp_p.n21650 16.399
R6600 vp_p.n21656 vp_p.n21655 16.399
R6601 vp_p.n21661 vp_p.n21660 16.399
R6602 vp_p.n21666 vp_p.n21665 16.399
R6603 vp_p.n21671 vp_p.n21670 16.399
R6604 vp_p.n21676 vp_p.n21675 16.399
R6605 vp_p.n21681 vp_p.n21680 16.399
R6606 vp_p.n21686 vp_p.n21685 16.399
R6607 vp_p.n21691 vp_p.n21690 16.399
R6608 vp_p.n21696 vp_p.n21695 16.399
R6609 vp_p.n21701 vp_p.n21700 16.399
R6610 vp_p.n21706 vp_p.n21705 16.399
R6611 vp_p.n21711 vp_p.n21710 16.399
R6612 vp_p.n21716 vp_p.n21715 16.399
R6613 vp_p.n21721 vp_p.n21720 16.399
R6614 vp_p.n21726 vp_p.n21725 16.399
R6615 vp_p.n21731 vp_p.n21730 16.399
R6616 vp_p.n21736 vp_p.n21735 16.399
R6617 vp_p.n21741 vp_p.n21740 16.399
R6618 vp_p.n21746 vp_p.n21745 16.399
R6619 vp_p.n21751 vp_p.n21750 16.399
R6620 vp_p.n21756 vp_p.n21755 16.399
R6621 vp_p.n21761 vp_p.n21760 16.399
R6622 vp_p.n21766 vp_p.n21765 16.399
R6623 vp_p.n21771 vp_p.n21770 16.399
R6624 vp_p.n21776 vp_p.n21775 16.399
R6625 vp_p.n21781 vp_p.n21780 16.399
R6626 vp_p.n21786 vp_p.n21785 16.399
R6627 vp_p.n21791 vp_p.n21790 16.399
R6628 vp_p.n21796 vp_p.n21795 16.399
R6629 vp_p.n21801 vp_p.n21800 16.399
R6630 vp_p.n21806 vp_p.n21805 16.399
R6631 vp_p.n21811 vp_p.n21810 16.399
R6632 vp_p.n21816 vp_p.n21815 16.399
R6633 vp_p.n21821 vp_p.n21820 16.399
R6634 vp_p.n21826 vp_p.n21825 16.399
R6635 vp_p.n21831 vp_p.n21830 16.399
R6636 vp_p.n21836 vp_p.n21835 16.399
R6637 vp_p.n21841 vp_p.n21840 16.399
R6638 vp_p.n21846 vp_p.n21845 16.399
R6639 vp_p.n21851 vp_p.n21850 16.399
R6640 vp_p.n21856 vp_p.n21855 16.399
R6641 vp_p.n21861 vp_p.n21860 16.399
R6642 vp_p.n21866 vp_p.n21865 16.399
R6643 vp_p.n21871 vp_p.n21870 16.399
R6644 vp_p.n21876 vp_p.n21875 16.399
R6645 vp_p.n21881 vp_p.n21880 16.399
R6646 vp_p.n21886 vp_p.n21885 16.399
R6647 vp_p.n21891 vp_p.n21890 16.399
R6648 vp_p.n21896 vp_p.n21895 16.399
R6649 vp_p.n21901 vp_p.n21900 16.399
R6650 vp_p.n21906 vp_p.n21905 16.399
R6651 vp_p.n21911 vp_p.n21910 16.399
R6652 vp_p.n21916 vp_p.n21915 16.399
R6653 vp_p.n21921 vp_p.n21920 16.399
R6654 vp_p.n21926 vp_p.n21925 16.399
R6655 vp_p.n21931 vp_p.n21930 16.399
R6656 vp_p.n21936 vp_p.n21935 16.399
R6657 vp_p.n21941 vp_p.n21940 16.399
R6658 vp_p.n21946 vp_p.n21945 16.399
R6659 vp_p.n21951 vp_p.n21950 16.399
R6660 vp_p.n21956 vp_p.n21955 16.399
R6661 vp_p.n21961 vp_p.n21960 16.399
R6662 vp_p.n21966 vp_p.n21965 16.399
R6663 vp_p.n21971 vp_p.n21970 16.399
R6664 vp_p.n21976 vp_p.n21975 16.399
R6665 vp_p.n21981 vp_p.n21980 16.399
R6666 vp_p.n21986 vp_p.n21985 16.399
R6667 vp_p.n21991 vp_p.n21990 16.399
R6668 vp_p.n21996 vp_p.n21995 16.399
R6669 vp_p.n22001 vp_p.n22000 16.399
R6670 vp_p.n4367 vp_p.n4366 16.399
R6671 vp_p.n4372 vp_p.n4371 16.399
R6672 vp_p.n4377 vp_p.n4376 16.399
R6673 vp_p.n4382 vp_p.n4381 16.399
R6674 vp_p.n4387 vp_p.n4386 16.399
R6675 vp_p.n4392 vp_p.n4391 16.399
R6676 vp_p.n4397 vp_p.n4396 16.399
R6677 vp_p.n4402 vp_p.n4401 16.399
R6678 vp_p.n4407 vp_p.n4406 16.399
R6679 vp_p.n4412 vp_p.n4411 16.399
R6680 vp_p.n4417 vp_p.n4416 16.399
R6681 vp_p.n4422 vp_p.n4421 16.399
R6682 vp_p.n4427 vp_p.n4426 16.399
R6683 vp_p.n4432 vp_p.n4431 16.399
R6684 vp_p.n4437 vp_p.n4436 16.399
R6685 vp_p.n4442 vp_p.n4441 16.399
R6686 vp_p.n4447 vp_p.n4446 16.399
R6687 vp_p.n4452 vp_p.n4451 16.399
R6688 vp_p.n4457 vp_p.n4456 16.399
R6689 vp_p.n4462 vp_p.n4461 16.399
R6690 vp_p.n4467 vp_p.n4466 16.399
R6691 vp_p.n4472 vp_p.n4471 16.399
R6692 vp_p.n4477 vp_p.n4476 16.399
R6693 vp_p.n4482 vp_p.n4481 16.399
R6694 vp_p.n4487 vp_p.n4486 16.399
R6695 vp_p.n4492 vp_p.n4491 16.399
R6696 vp_p.n4497 vp_p.n4496 16.399
R6697 vp_p.n4502 vp_p.n4501 16.399
R6698 vp_p.n4507 vp_p.n4506 16.399
R6699 vp_p.n4512 vp_p.n4511 16.399
R6700 vp_p.n4517 vp_p.n4516 16.399
R6701 vp_p.n4522 vp_p.n4521 16.399
R6702 vp_p.n4527 vp_p.n4526 16.399
R6703 vp_p.n4532 vp_p.n4531 16.399
R6704 vp_p.n4537 vp_p.n4536 16.399
R6705 vp_p.n4542 vp_p.n4541 16.399
R6706 vp_p.n4547 vp_p.n4546 16.399
R6707 vp_p.n4552 vp_p.n4551 16.399
R6708 vp_p.n4557 vp_p.n4556 16.399
R6709 vp_p.n4562 vp_p.n4561 16.399
R6710 vp_p.n4567 vp_p.n4566 16.399
R6711 vp_p.n4572 vp_p.n4571 16.399
R6712 vp_p.n4577 vp_p.n4576 16.399
R6713 vp_p.n4582 vp_p.n4581 16.399
R6714 vp_p.n4587 vp_p.n4586 16.399
R6715 vp_p.n4592 vp_p.n4591 16.399
R6716 vp_p.n4597 vp_p.n4596 16.399
R6717 vp_p.n4602 vp_p.n4601 16.399
R6718 vp_p.n4607 vp_p.n4606 16.399
R6719 vp_p.n4612 vp_p.n4611 16.399
R6720 vp_p.n4617 vp_p.n4616 16.399
R6721 vp_p.n4622 vp_p.n4621 16.399
R6722 vp_p.n4627 vp_p.n4626 16.399
R6723 vp_p.n4632 vp_p.n4631 16.399
R6724 vp_p.n4637 vp_p.n4636 16.399
R6725 vp_p.n4642 vp_p.n4641 16.399
R6726 vp_p.n4647 vp_p.n4646 16.399
R6727 vp_p.n4652 vp_p.n4651 16.399
R6728 vp_p.n4657 vp_p.n4656 16.399
R6729 vp_p.n4662 vp_p.n4661 16.399
R6730 vp_p.n4667 vp_p.n4666 16.399
R6731 vp_p.n4672 vp_p.n4671 16.399
R6732 vp_p.n4677 vp_p.n4676 16.399
R6733 vp_p.n4682 vp_p.n4681 16.399
R6734 vp_p.n4687 vp_p.n4686 16.399
R6735 vp_p.n4692 vp_p.n4691 16.399
R6736 vp_p.n4697 vp_p.n4696 16.399
R6737 vp_p.n4702 vp_p.n4701 16.399
R6738 vp_p.n4707 vp_p.n4706 16.399
R6739 vp_p.n4712 vp_p.n4711 16.399
R6740 vp_p.n4717 vp_p.n4716 16.399
R6741 vp_p.n4722 vp_p.n4721 16.399
R6742 vp_p.n23064 vp_p.n23063 16.399
R6743 vp_p.n23069 vp_p.n23068 16.399
R6744 vp_p.n23074 vp_p.n23073 16.399
R6745 vp_p.n23079 vp_p.n23078 16.399
R6746 vp_p.n23084 vp_p.n23083 16.399
R6747 vp_p.n23089 vp_p.n23088 16.399
R6748 vp_p.n23094 vp_p.n23093 16.399
R6749 vp_p.n23099 vp_p.n23098 16.399
R6750 vp_p.n23104 vp_p.n23103 16.399
R6751 vp_p.n23109 vp_p.n23108 16.399
R6752 vp_p.n23114 vp_p.n23113 16.399
R6753 vp_p.n23119 vp_p.n23118 16.399
R6754 vp_p.n23124 vp_p.n23123 16.399
R6755 vp_p.n23129 vp_p.n23128 16.399
R6756 vp_p.n23134 vp_p.n23133 16.399
R6757 vp_p.n23139 vp_p.n23138 16.399
R6758 vp_p.n23144 vp_p.n23143 16.399
R6759 vp_p.n23149 vp_p.n23148 16.399
R6760 vp_p.n23154 vp_p.n23153 16.399
R6761 vp_p.n23159 vp_p.n23158 16.399
R6762 vp_p.n23164 vp_p.n23163 16.399
R6763 vp_p.n23169 vp_p.n23168 16.399
R6764 vp_p.n23174 vp_p.n23173 16.399
R6765 vp_p.n23179 vp_p.n23178 16.399
R6766 vp_p.n23184 vp_p.n23183 16.399
R6767 vp_p.n23189 vp_p.n23188 16.399
R6768 vp_p.n23194 vp_p.n23193 16.399
R6769 vp_p.n23199 vp_p.n23198 16.399
R6770 vp_p.n23204 vp_p.n23203 16.399
R6771 vp_p.n23209 vp_p.n23208 16.399
R6772 vp_p.n23214 vp_p.n23213 16.399
R6773 vp_p.n23219 vp_p.n23218 16.399
R6774 vp_p.n23224 vp_p.n23223 16.399
R6775 vp_p.n23229 vp_p.n23228 16.399
R6776 vp_p.n23234 vp_p.n23233 16.399
R6777 vp_p.n23239 vp_p.n23238 16.399
R6778 vp_p.n23244 vp_p.n23243 16.399
R6779 vp_p.n23249 vp_p.n23248 16.399
R6780 vp_p.n23254 vp_p.n23253 16.399
R6781 vp_p.n23259 vp_p.n23258 16.399
R6782 vp_p.n23264 vp_p.n23263 16.399
R6783 vp_p.n23269 vp_p.n23268 16.399
R6784 vp_p.n23274 vp_p.n23273 16.399
R6785 vp_p.n23279 vp_p.n23278 16.399
R6786 vp_p.n23284 vp_p.n23283 16.399
R6787 vp_p.n23289 vp_p.n23288 16.399
R6788 vp_p.n23294 vp_p.n23293 16.399
R6789 vp_p.n23299 vp_p.n23298 16.399
R6790 vp_p.n23304 vp_p.n23303 16.399
R6791 vp_p.n23309 vp_p.n23308 16.399
R6792 vp_p.n23314 vp_p.n23313 16.399
R6793 vp_p.n23319 vp_p.n23318 16.399
R6794 vp_p.n23324 vp_p.n23323 16.399
R6795 vp_p.n23329 vp_p.n23328 16.399
R6796 vp_p.n23334 vp_p.n23333 16.399
R6797 vp_p.n23339 vp_p.n23338 16.399
R6798 vp_p.n23344 vp_p.n23343 16.399
R6799 vp_p.n23349 vp_p.n23348 16.399
R6800 vp_p.n23354 vp_p.n23353 16.399
R6801 vp_p.n23359 vp_p.n23358 16.399
R6802 vp_p.n23364 vp_p.n23363 16.399
R6803 vp_p.n23369 vp_p.n23368 16.399
R6804 vp_p.n23374 vp_p.n23373 16.399
R6805 vp_p.n23379 vp_p.n23378 16.399
R6806 vp_p.n23384 vp_p.n23383 16.399
R6807 vp_p.n23389 vp_p.n23388 16.399
R6808 vp_p.n23394 vp_p.n23393 16.399
R6809 vp_p.n23399 vp_p.n23398 16.399
R6810 vp_p.n23404 vp_p.n23403 16.399
R6811 vp_p.n23409 vp_p.n23408 16.399
R6812 vp_p.n23414 vp_p.n23413 16.399
R6813 vp_p.n23419 vp_p.n23418 16.399
R6814 vp_p.n23424 vp_p.n23423 16.399
R6815 vp_p.n5785 vp_p.n5784 16.399
R6816 vp_p.n5790 vp_p.n5789 16.399
R6817 vp_p.n5795 vp_p.n5794 16.399
R6818 vp_p.n5800 vp_p.n5799 16.399
R6819 vp_p.n5805 vp_p.n5804 16.399
R6820 vp_p.n5810 vp_p.n5809 16.399
R6821 vp_p.n5815 vp_p.n5814 16.399
R6822 vp_p.n5820 vp_p.n5819 16.399
R6823 vp_p.n5825 vp_p.n5824 16.399
R6824 vp_p.n5830 vp_p.n5829 16.399
R6825 vp_p.n5835 vp_p.n5834 16.399
R6826 vp_p.n5840 vp_p.n5839 16.399
R6827 vp_p.n5845 vp_p.n5844 16.399
R6828 vp_p.n5850 vp_p.n5849 16.399
R6829 vp_p.n5855 vp_p.n5854 16.399
R6830 vp_p.n5860 vp_p.n5859 16.399
R6831 vp_p.n5865 vp_p.n5864 16.399
R6832 vp_p.n5870 vp_p.n5869 16.399
R6833 vp_p.n5875 vp_p.n5874 16.399
R6834 vp_p.n5880 vp_p.n5879 16.399
R6835 vp_p.n5885 vp_p.n5884 16.399
R6836 vp_p.n5890 vp_p.n5889 16.399
R6837 vp_p.n5895 vp_p.n5894 16.399
R6838 vp_p.n5900 vp_p.n5899 16.399
R6839 vp_p.n5905 vp_p.n5904 16.399
R6840 vp_p.n5910 vp_p.n5909 16.399
R6841 vp_p.n5915 vp_p.n5914 16.399
R6842 vp_p.n5920 vp_p.n5919 16.399
R6843 vp_p.n5925 vp_p.n5924 16.399
R6844 vp_p.n5930 vp_p.n5929 16.399
R6845 vp_p.n5935 vp_p.n5934 16.399
R6846 vp_p.n5940 vp_p.n5939 16.399
R6847 vp_p.n5945 vp_p.n5944 16.399
R6848 vp_p.n5950 vp_p.n5949 16.399
R6849 vp_p.n5955 vp_p.n5954 16.399
R6850 vp_p.n5960 vp_p.n5959 16.399
R6851 vp_p.n5965 vp_p.n5964 16.399
R6852 vp_p.n5970 vp_p.n5969 16.399
R6853 vp_p.n5975 vp_p.n5974 16.399
R6854 vp_p.n5980 vp_p.n5979 16.399
R6855 vp_p.n5985 vp_p.n5984 16.399
R6856 vp_p.n5990 vp_p.n5989 16.399
R6857 vp_p.n5995 vp_p.n5994 16.399
R6858 vp_p.n6000 vp_p.n5999 16.399
R6859 vp_p.n6005 vp_p.n6004 16.399
R6860 vp_p.n6010 vp_p.n6009 16.399
R6861 vp_p.n6015 vp_p.n6014 16.399
R6862 vp_p.n6020 vp_p.n6019 16.399
R6863 vp_p.n6025 vp_p.n6024 16.399
R6864 vp_p.n6030 vp_p.n6029 16.399
R6865 vp_p.n6035 vp_p.n6034 16.399
R6866 vp_p.n6040 vp_p.n6039 16.399
R6867 vp_p.n6045 vp_p.n6044 16.399
R6868 vp_p.n6050 vp_p.n6049 16.399
R6869 vp_p.n6055 vp_p.n6054 16.399
R6870 vp_p.n6060 vp_p.n6059 16.399
R6871 vp_p.n6065 vp_p.n6064 16.399
R6872 vp_p.n6070 vp_p.n6069 16.399
R6873 vp_p.n6075 vp_p.n6074 16.399
R6874 vp_p.n6080 vp_p.n6079 16.399
R6875 vp_p.n6085 vp_p.n6084 16.399
R6876 vp_p.n6090 vp_p.n6089 16.399
R6877 vp_p.n6095 vp_p.n6094 16.399
R6878 vp_p.n6100 vp_p.n6099 16.399
R6879 vp_p.n6105 vp_p.n6104 16.399
R6880 vp_p.n6110 vp_p.n6109 16.399
R6881 vp_p.n6115 vp_p.n6114 16.399
R6882 vp_p.n6120 vp_p.n6119 16.399
R6883 vp_p.n6125 vp_p.n6124 16.399
R6884 vp_p.n6130 vp_p.n6129 16.399
R6885 vp_p.n6135 vp_p.n6134 16.399
R6886 vp_p.n6140 vp_p.n6139 16.399
R6887 vp_p.n6145 vp_p.n6144 16.399
R6888 vp_p.n24481 vp_p.n24480 16.399
R6889 vp_p.n24486 vp_p.n24485 16.399
R6890 vp_p.n24491 vp_p.n24490 16.399
R6891 vp_p.n24496 vp_p.n24495 16.399
R6892 vp_p.n24501 vp_p.n24500 16.399
R6893 vp_p.n24506 vp_p.n24505 16.399
R6894 vp_p.n24511 vp_p.n24510 16.399
R6895 vp_p.n24516 vp_p.n24515 16.399
R6896 vp_p.n24521 vp_p.n24520 16.399
R6897 vp_p.n24526 vp_p.n24525 16.399
R6898 vp_p.n24531 vp_p.n24530 16.399
R6899 vp_p.n24536 vp_p.n24535 16.399
R6900 vp_p.n24541 vp_p.n24540 16.399
R6901 vp_p.n24546 vp_p.n24545 16.399
R6902 vp_p.n24551 vp_p.n24550 16.399
R6903 vp_p.n24556 vp_p.n24555 16.399
R6904 vp_p.n24561 vp_p.n24560 16.399
R6905 vp_p.n24566 vp_p.n24565 16.399
R6906 vp_p.n24571 vp_p.n24570 16.399
R6907 vp_p.n24576 vp_p.n24575 16.399
R6908 vp_p.n24581 vp_p.n24580 16.399
R6909 vp_p.n24586 vp_p.n24585 16.399
R6910 vp_p.n24591 vp_p.n24590 16.399
R6911 vp_p.n24596 vp_p.n24595 16.399
R6912 vp_p.n24601 vp_p.n24600 16.399
R6913 vp_p.n24606 vp_p.n24605 16.399
R6914 vp_p.n24611 vp_p.n24610 16.399
R6915 vp_p.n24616 vp_p.n24615 16.399
R6916 vp_p.n24621 vp_p.n24620 16.399
R6917 vp_p.n24626 vp_p.n24625 16.399
R6918 vp_p.n24631 vp_p.n24630 16.399
R6919 vp_p.n24636 vp_p.n24635 16.399
R6920 vp_p.n24641 vp_p.n24640 16.399
R6921 vp_p.n24646 vp_p.n24645 16.399
R6922 vp_p.n24651 vp_p.n24650 16.399
R6923 vp_p.n24656 vp_p.n24655 16.399
R6924 vp_p.n24661 vp_p.n24660 16.399
R6925 vp_p.n24666 vp_p.n24665 16.399
R6926 vp_p.n24671 vp_p.n24670 16.399
R6927 vp_p.n24676 vp_p.n24675 16.399
R6928 vp_p.n24681 vp_p.n24680 16.399
R6929 vp_p.n24686 vp_p.n24685 16.399
R6930 vp_p.n24691 vp_p.n24690 16.399
R6931 vp_p.n24696 vp_p.n24695 16.399
R6932 vp_p.n24701 vp_p.n24700 16.399
R6933 vp_p.n24706 vp_p.n24705 16.399
R6934 vp_p.n24711 vp_p.n24710 16.399
R6935 vp_p.n24716 vp_p.n24715 16.399
R6936 vp_p.n24721 vp_p.n24720 16.399
R6937 vp_p.n24726 vp_p.n24725 16.399
R6938 vp_p.n24731 vp_p.n24730 16.399
R6939 vp_p.n24736 vp_p.n24735 16.399
R6940 vp_p.n24741 vp_p.n24740 16.399
R6941 vp_p.n24746 vp_p.n24745 16.399
R6942 vp_p.n24751 vp_p.n24750 16.399
R6943 vp_p.n24756 vp_p.n24755 16.399
R6944 vp_p.n24761 vp_p.n24760 16.399
R6945 vp_p.n24766 vp_p.n24765 16.399
R6946 vp_p.n24771 vp_p.n24770 16.399
R6947 vp_p.n24776 vp_p.n24775 16.399
R6948 vp_p.n24781 vp_p.n24780 16.399
R6949 vp_p.n24786 vp_p.n24785 16.399
R6950 vp_p.n24791 vp_p.n24790 16.399
R6951 vp_p.n24796 vp_p.n24795 16.399
R6952 vp_p.n24801 vp_p.n24800 16.399
R6953 vp_p.n24806 vp_p.n24805 16.399
R6954 vp_p.n24811 vp_p.n24810 16.399
R6955 vp_p.n24816 vp_p.n24815 16.399
R6956 vp_p.n24821 vp_p.n24820 16.399
R6957 vp_p.n24826 vp_p.n24825 16.399
R6958 vp_p.n24831 vp_p.n24830 16.399
R6959 vp_p.n24836 vp_p.n24835 16.399
R6960 vp_p.n24841 vp_p.n24840 16.399
R6961 vp_p.n24846 vp_p.n24845 16.399
R6962 vp_p.n7567 vp_p.n7566 16.399
R6963 vp_p.n7562 vp_p.n7561 16.399
R6964 vp_p.n7557 vp_p.n7556 16.399
R6965 vp_p.n7552 vp_p.n7551 16.399
R6966 vp_p.n7547 vp_p.n7546 16.399
R6967 vp_p.n7542 vp_p.n7541 16.399
R6968 vp_p.n7537 vp_p.n7536 16.399
R6969 vp_p.n7532 vp_p.n7531 16.399
R6970 vp_p.n7527 vp_p.n7526 16.399
R6971 vp_p.n7522 vp_p.n7521 16.399
R6972 vp_p.n7517 vp_p.n7516 16.399
R6973 vp_p.n7512 vp_p.n7511 16.399
R6974 vp_p.n7507 vp_p.n7506 16.399
R6975 vp_p.n7502 vp_p.n7501 16.399
R6976 vp_p.n7497 vp_p.n7496 16.399
R6977 vp_p.n7492 vp_p.n7491 16.399
R6978 vp_p.n7487 vp_p.n7486 16.399
R6979 vp_p.n7482 vp_p.n7481 16.399
R6980 vp_p.n7477 vp_p.n7476 16.399
R6981 vp_p.n7472 vp_p.n7471 16.399
R6982 vp_p.n7467 vp_p.n7466 16.399
R6983 vp_p.n7462 vp_p.n7461 16.399
R6984 vp_p.n7457 vp_p.n7456 16.399
R6985 vp_p.n7452 vp_p.n7451 16.399
R6986 vp_p.n7447 vp_p.n7446 16.399
R6987 vp_p.n7442 vp_p.n7441 16.399
R6988 vp_p.n7437 vp_p.n7436 16.399
R6989 vp_p.n7432 vp_p.n7431 16.399
R6990 vp_p.n7427 vp_p.n7426 16.399
R6991 vp_p.n7422 vp_p.n7421 16.399
R6992 vp_p.n7417 vp_p.n7416 16.399
R6993 vp_p.n7412 vp_p.n7411 16.399
R6994 vp_p.n7407 vp_p.n7406 16.399
R6995 vp_p.n7402 vp_p.n7401 16.399
R6996 vp_p.n7397 vp_p.n7396 16.399
R6997 vp_p.n7392 vp_p.n7391 16.399
R6998 vp_p.n7387 vp_p.n7386 16.399
R6999 vp_p.n7382 vp_p.n7381 16.399
R7000 vp_p.n7377 vp_p.n7376 16.399
R7001 vp_p.n7372 vp_p.n7371 16.399
R7002 vp_p.n7367 vp_p.n7366 16.399
R7003 vp_p.n7362 vp_p.n7361 16.399
R7004 vp_p.n7357 vp_p.n7356 16.399
R7005 vp_p.n7352 vp_p.n7351 16.399
R7006 vp_p.n7347 vp_p.n7346 16.399
R7007 vp_p.n7342 vp_p.n7341 16.399
R7008 vp_p.n7337 vp_p.n7336 16.399
R7009 vp_p.n7332 vp_p.n7331 16.399
R7010 vp_p.n7327 vp_p.n7326 16.399
R7011 vp_p.n7322 vp_p.n7321 16.399
R7012 vp_p.n7317 vp_p.n7316 16.399
R7013 vp_p.n7312 vp_p.n7311 16.399
R7014 vp_p.n7307 vp_p.n7306 16.399
R7015 vp_p.n7302 vp_p.n7301 16.399
R7016 vp_p.n7297 vp_p.n7296 16.399
R7017 vp_p.n7292 vp_p.n7291 16.399
R7018 vp_p.n7287 vp_p.n7286 16.399
R7019 vp_p.n7282 vp_p.n7281 16.399
R7020 vp_p.n7277 vp_p.n7276 16.399
R7021 vp_p.n7272 vp_p.n7271 16.399
R7022 vp_p.n7267 vp_p.n7266 16.399
R7023 vp_p.n7262 vp_p.n7261 16.399
R7024 vp_p.n7257 vp_p.n7256 16.399
R7025 vp_p.n7252 vp_p.n7251 16.399
R7026 vp_p.n7247 vp_p.n7246 16.399
R7027 vp_p.n7242 vp_p.n7241 16.399
R7028 vp_p.n7237 vp_p.n7236 16.399
R7029 vp_p.n7232 vp_p.n7231 16.399
R7030 vp_p.n7227 vp_p.n7226 16.399
R7031 vp_p.n7222 vp_p.n7221 16.399
R7032 vp_p.n7217 vp_p.n7216 16.399
R7033 vp_p.n7212 vp_p.n7211 16.399
R7034 vp_p.n7207 vp_p.n7206 16.399
R7035 vp_p.n26277 vp_p.n26276 16.399
R7036 vp_p.n26272 vp_p.n26271 16.399
R7037 vp_p.n26267 vp_p.n26266 16.399
R7038 vp_p.n26262 vp_p.n26261 16.399
R7039 vp_p.n26257 vp_p.n26256 16.399
R7040 vp_p.n26252 vp_p.n26251 16.399
R7041 vp_p.n26247 vp_p.n26246 16.399
R7042 vp_p.n26242 vp_p.n26241 16.399
R7043 vp_p.n26237 vp_p.n26236 16.399
R7044 vp_p.n26232 vp_p.n26231 16.399
R7045 vp_p.n26227 vp_p.n26226 16.399
R7046 vp_p.n26222 vp_p.n26221 16.399
R7047 vp_p.n26217 vp_p.n26216 16.399
R7048 vp_p.n26212 vp_p.n26211 16.399
R7049 vp_p.n26207 vp_p.n26206 16.399
R7050 vp_p.n26202 vp_p.n26201 16.399
R7051 vp_p.n26197 vp_p.n26196 16.399
R7052 vp_p.n26192 vp_p.n26191 16.399
R7053 vp_p.n26187 vp_p.n26186 16.399
R7054 vp_p.n26182 vp_p.n26181 16.399
R7055 vp_p.n26177 vp_p.n26176 16.399
R7056 vp_p.n26172 vp_p.n26171 16.399
R7057 vp_p.n26167 vp_p.n26166 16.399
R7058 vp_p.n26162 vp_p.n26161 16.399
R7059 vp_p.n26157 vp_p.n26156 16.399
R7060 vp_p.n26152 vp_p.n26151 16.399
R7061 vp_p.n26147 vp_p.n26146 16.399
R7062 vp_p.n26142 vp_p.n26141 16.399
R7063 vp_p.n26137 vp_p.n26136 16.399
R7064 vp_p.n26132 vp_p.n26131 16.399
R7065 vp_p.n26127 vp_p.n26126 16.399
R7066 vp_p.n26122 vp_p.n26121 16.399
R7067 vp_p.n26117 vp_p.n26116 16.399
R7068 vp_p.n26112 vp_p.n26111 16.399
R7069 vp_p.n26107 vp_p.n26106 16.399
R7070 vp_p.n26102 vp_p.n26101 16.399
R7071 vp_p.n26097 vp_p.n26096 16.399
R7072 vp_p.n26092 vp_p.n26091 16.399
R7073 vp_p.n26087 vp_p.n26086 16.399
R7074 vp_p.n26082 vp_p.n26081 16.399
R7075 vp_p.n26077 vp_p.n26076 16.399
R7076 vp_p.n26072 vp_p.n26071 16.399
R7077 vp_p.n26067 vp_p.n26066 16.399
R7078 vp_p.n26062 vp_p.n26061 16.399
R7079 vp_p.n26057 vp_p.n26056 16.399
R7080 vp_p.n26052 vp_p.n26051 16.399
R7081 vp_p.n26047 vp_p.n26046 16.399
R7082 vp_p.n26042 vp_p.n26041 16.399
R7083 vp_p.n26037 vp_p.n26036 16.399
R7084 vp_p.n26032 vp_p.n26031 16.399
R7085 vp_p.n26027 vp_p.n26026 16.399
R7086 vp_p.n26022 vp_p.n26021 16.399
R7087 vp_p.n26017 vp_p.n26016 16.399
R7088 vp_p.n26012 vp_p.n26011 16.399
R7089 vp_p.n26007 vp_p.n26006 16.399
R7090 vp_p.n26002 vp_p.n26001 16.399
R7091 vp_p.n25997 vp_p.n25996 16.399
R7092 vp_p.n25992 vp_p.n25991 16.399
R7093 vp_p.n25987 vp_p.n25986 16.399
R7094 vp_p.n25982 vp_p.n25981 16.399
R7095 vp_p.n25977 vp_p.n25976 16.399
R7096 vp_p.n25972 vp_p.n25971 16.399
R7097 vp_p.n25967 vp_p.n25966 16.399
R7098 vp_p.n25962 vp_p.n25961 16.399
R7099 vp_p.n25957 vp_p.n25956 16.399
R7100 vp_p.n25952 vp_p.n25951 16.399
R7101 vp_p.n25947 vp_p.n25946 16.399
R7102 vp_p.n25942 vp_p.n25941 16.399
R7103 vp_p.n25937 vp_p.n25936 16.399
R7104 vp_p.n25932 vp_p.n25931 16.399
R7105 vp_p.n25927 vp_p.n25926 16.399
R7106 vp_p.n25922 vp_p.n25921 16.399
R7107 vp_p.n25917 vp_p.n25916 16.399
R7108 vp_p.n25912 vp_p.n25911 16.399
R7109 vp_p.n25907 vp_p.n25906 16.399
R7110 vp_p.n26284 vp_p.n26283 16.399
R7111 vp_p.n7207 vp_p.n7204 14.806
R7112 vp_p.n5790 vp_p.n5787 14.806
R7113 vp_p.n7212 vp_p.n7209 14.806
R7114 vp_p.n4372 vp_p.n4369 14.806
R7115 vp_p.n5795 vp_p.n5792 14.806
R7116 vp_p.n7217 vp_p.n7214 14.806
R7117 vp_p.n2953 vp_p.n2950 14.806
R7118 vp_p.n4377 vp_p.n4374 14.806
R7119 vp_p.n5800 vp_p.n5797 14.806
R7120 vp_p.n7222 vp_p.n7219 14.806
R7121 vp_p.n1533 vp_p.n1530 14.806
R7122 vp_p.n2958 vp_p.n2955 14.806
R7123 vp_p.n4382 vp_p.n4379 14.806
R7124 vp_p.n5805 vp_p.n5802 14.806
R7125 vp_p.n7227 vp_p.n7224 14.806
R7126 vp_p.n54 vp_p.n51 14.806
R7127 vp_p.n1538 vp_p.n1535 14.806
R7128 vp_p.n2963 vp_p.n2960 14.806
R7129 vp_p.n4387 vp_p.n4384 14.806
R7130 vp_p.n5810 vp_p.n5807 14.806
R7131 vp_p.n7232 vp_p.n7229 14.806
R7132 vp_p.n8798 vp_p.n8795 14.806
R7133 vp_p.n59 vp_p.n56 14.806
R7134 vp_p.n1543 vp_p.n1540 14.806
R7135 vp_p.n2968 vp_p.n2965 14.806
R7136 vp_p.n4392 vp_p.n4389 14.806
R7137 vp_p.n5815 vp_p.n5812 14.806
R7138 vp_p.n7237 vp_p.n7234 14.806
R7139 vp_p.n10305 vp_p.n10302 14.806
R7140 vp_p.n8803 vp_p.n8800 14.806
R7141 vp_p.n64 vp_p.n61 14.806
R7142 vp_p.n1548 vp_p.n1545 14.806
R7143 vp_p.n2973 vp_p.n2970 14.806
R7144 vp_p.n4397 vp_p.n4394 14.806
R7145 vp_p.n5820 vp_p.n5817 14.806
R7146 vp_p.n7242 vp_p.n7239 14.806
R7147 vp_p.n13832 vp_p.n13829 14.806
R7148 vp_p.n12068 vp_p.n12065 14.806
R7149 vp_p.n10630 vp_p.n10627 14.806
R7150 vp_p.n9128 vp_p.n9125 14.806
R7151 vp_p.n389 vp_p.n386 14.806
R7152 vp_p.n1873 vp_p.n1870 14.806
R7153 vp_p.n3298 vp_p.n3295 14.806
R7154 vp_p.n4722 vp_p.n4719 14.806
R7155 vp_p.n6145 vp_p.n6142 14.806
R7156 vp_p.n7567 vp_p.n7564 14.806
R7157 vp_p.n14871 vp_p.n14868 14.806
R7158 vp_p.n16299 vp_p.n16296 14.806
R7159 vp_p.n17726 vp_p.n17723 14.806
R7160 vp_p.n19152 vp_p.n19149 14.806
R7161 vp_p.n20577 vp_p.n20574 14.806
R7162 vp_p.n22001 vp_p.n21998 14.806
R7163 vp_p.n23424 vp_p.n23421 14.806
R7164 vp_p.n24846 vp_p.n24843 14.806
R7165 vp_p.n26272 vp_p.n26269 14.806
R7166 vp_p.n13827 vp_p.n13824 14.806
R7167 vp_p.n13822 vp_p.n13819 14.806
R7168 vp_p.n12063 vp_p.n12060 14.806
R7169 vp_p.n10625 vp_p.n10622 14.806
R7170 vp_p.n9123 vp_p.n9120 14.806
R7171 vp_p.n384 vp_p.n381 14.806
R7172 vp_p.n1868 vp_p.n1865 14.806
R7173 vp_p.n3293 vp_p.n3290 14.806
R7174 vp_p.n4717 vp_p.n4714 14.806
R7175 vp_p.n6140 vp_p.n6137 14.806
R7176 vp_p.n7562 vp_p.n7559 14.806
R7177 vp_p.n14866 vp_p.n14863 14.806
R7178 vp_p.n16294 vp_p.n16291 14.806
R7179 vp_p.n17721 vp_p.n17718 14.806
R7180 vp_p.n19147 vp_p.n19144 14.806
R7181 vp_p.n20572 vp_p.n20569 14.806
R7182 vp_p.n21996 vp_p.n21993 14.806
R7183 vp_p.n23419 vp_p.n23416 14.806
R7184 vp_p.n24841 vp_p.n24838 14.806
R7185 vp_p.n26267 vp_p.n26264 14.806
R7186 vp_p.n13817 vp_p.n13814 14.806
R7187 vp_p.n13812 vp_p.n13809 14.806
R7188 vp_p.n12058 vp_p.n12055 14.806
R7189 vp_p.n10620 vp_p.n10617 14.806
R7190 vp_p.n9118 vp_p.n9115 14.806
R7191 vp_p.n379 vp_p.n376 14.806
R7192 vp_p.n1863 vp_p.n1860 14.806
R7193 vp_p.n3288 vp_p.n3285 14.806
R7194 vp_p.n4712 vp_p.n4709 14.806
R7195 vp_p.n6135 vp_p.n6132 14.806
R7196 vp_p.n7557 vp_p.n7554 14.806
R7197 vp_p.n14861 vp_p.n14858 14.806
R7198 vp_p.n16289 vp_p.n16286 14.806
R7199 vp_p.n17716 vp_p.n17713 14.806
R7200 vp_p.n19142 vp_p.n19139 14.806
R7201 vp_p.n20567 vp_p.n20564 14.806
R7202 vp_p.n21991 vp_p.n21988 14.806
R7203 vp_p.n23414 vp_p.n23411 14.806
R7204 vp_p.n24836 vp_p.n24833 14.806
R7205 vp_p.n26262 vp_p.n26259 14.806
R7206 vp_p.n13807 vp_p.n13804 14.806
R7207 vp_p.n13802 vp_p.n13799 14.806
R7208 vp_p.n12053 vp_p.n12050 14.806
R7209 vp_p.n10615 vp_p.n10612 14.806
R7210 vp_p.n9113 vp_p.n9110 14.806
R7211 vp_p.n374 vp_p.n371 14.806
R7212 vp_p.n1858 vp_p.n1855 14.806
R7213 vp_p.n3283 vp_p.n3280 14.806
R7214 vp_p.n4707 vp_p.n4704 14.806
R7215 vp_p.n6130 vp_p.n6127 14.806
R7216 vp_p.n7552 vp_p.n7549 14.806
R7217 vp_p.n14856 vp_p.n14853 14.806
R7218 vp_p.n16284 vp_p.n16281 14.806
R7219 vp_p.n17711 vp_p.n17708 14.806
R7220 vp_p.n19137 vp_p.n19134 14.806
R7221 vp_p.n20562 vp_p.n20559 14.806
R7222 vp_p.n21986 vp_p.n21983 14.806
R7223 vp_p.n23409 vp_p.n23406 14.806
R7224 vp_p.n24831 vp_p.n24828 14.806
R7225 vp_p.n26257 vp_p.n26254 14.806
R7226 vp_p.n13797 vp_p.n13794 14.806
R7227 vp_p.n13792 vp_p.n13789 14.806
R7228 vp_p.n12048 vp_p.n12045 14.806
R7229 vp_p.n10610 vp_p.n10607 14.806
R7230 vp_p.n9108 vp_p.n9105 14.806
R7231 vp_p.n369 vp_p.n366 14.806
R7232 vp_p.n1853 vp_p.n1850 14.806
R7233 vp_p.n3278 vp_p.n3275 14.806
R7234 vp_p.n4702 vp_p.n4699 14.806
R7235 vp_p.n6125 vp_p.n6122 14.806
R7236 vp_p.n7547 vp_p.n7544 14.806
R7237 vp_p.n14851 vp_p.n14848 14.806
R7238 vp_p.n16279 vp_p.n16276 14.806
R7239 vp_p.n17706 vp_p.n17703 14.806
R7240 vp_p.n19132 vp_p.n19129 14.806
R7241 vp_p.n20557 vp_p.n20554 14.806
R7242 vp_p.n21981 vp_p.n21978 14.806
R7243 vp_p.n23404 vp_p.n23401 14.806
R7244 vp_p.n24826 vp_p.n24823 14.806
R7245 vp_p.n26252 vp_p.n26249 14.806
R7246 vp_p.n13787 vp_p.n13784 14.806
R7247 vp_p.n13782 vp_p.n13779 14.806
R7248 vp_p.n12043 vp_p.n12040 14.806
R7249 vp_p.n10605 vp_p.n10602 14.806
R7250 vp_p.n9103 vp_p.n9100 14.806
R7251 vp_p.n364 vp_p.n361 14.806
R7252 vp_p.n1848 vp_p.n1845 14.806
R7253 vp_p.n3273 vp_p.n3270 14.806
R7254 vp_p.n4697 vp_p.n4694 14.806
R7255 vp_p.n6120 vp_p.n6117 14.806
R7256 vp_p.n7542 vp_p.n7539 14.806
R7257 vp_p.n14846 vp_p.n14843 14.806
R7258 vp_p.n16274 vp_p.n16271 14.806
R7259 vp_p.n17701 vp_p.n17698 14.806
R7260 vp_p.n19127 vp_p.n19124 14.806
R7261 vp_p.n20552 vp_p.n20549 14.806
R7262 vp_p.n21976 vp_p.n21973 14.806
R7263 vp_p.n23399 vp_p.n23396 14.806
R7264 vp_p.n24821 vp_p.n24818 14.806
R7265 vp_p.n26247 vp_p.n26244 14.806
R7266 vp_p.n13777 vp_p.n13774 14.806
R7267 vp_p.n13772 vp_p.n13769 14.806
R7268 vp_p.n12038 vp_p.n12035 14.806
R7269 vp_p.n10600 vp_p.n10597 14.806
R7270 vp_p.n9098 vp_p.n9095 14.806
R7271 vp_p.n359 vp_p.n356 14.806
R7272 vp_p.n1843 vp_p.n1840 14.806
R7273 vp_p.n3268 vp_p.n3265 14.806
R7274 vp_p.n4692 vp_p.n4689 14.806
R7275 vp_p.n6115 vp_p.n6112 14.806
R7276 vp_p.n7537 vp_p.n7534 14.806
R7277 vp_p.n14841 vp_p.n14838 14.806
R7278 vp_p.n16269 vp_p.n16266 14.806
R7279 vp_p.n17696 vp_p.n17693 14.806
R7280 vp_p.n19122 vp_p.n19119 14.806
R7281 vp_p.n20547 vp_p.n20544 14.806
R7282 vp_p.n21971 vp_p.n21968 14.806
R7283 vp_p.n23394 vp_p.n23391 14.806
R7284 vp_p.n24816 vp_p.n24813 14.806
R7285 vp_p.n26242 vp_p.n26239 14.806
R7286 vp_p.n13767 vp_p.n13764 14.806
R7287 vp_p.n13762 vp_p.n13759 14.806
R7288 vp_p.n12033 vp_p.n12030 14.806
R7289 vp_p.n10595 vp_p.n10592 14.806
R7290 vp_p.n9093 vp_p.n9090 14.806
R7291 vp_p.n354 vp_p.n351 14.806
R7292 vp_p.n1838 vp_p.n1835 14.806
R7293 vp_p.n3263 vp_p.n3260 14.806
R7294 vp_p.n4687 vp_p.n4684 14.806
R7295 vp_p.n6110 vp_p.n6107 14.806
R7296 vp_p.n7532 vp_p.n7529 14.806
R7297 vp_p.n14836 vp_p.n14833 14.806
R7298 vp_p.n16264 vp_p.n16261 14.806
R7299 vp_p.n17691 vp_p.n17688 14.806
R7300 vp_p.n19117 vp_p.n19114 14.806
R7301 vp_p.n20542 vp_p.n20539 14.806
R7302 vp_p.n21966 vp_p.n21963 14.806
R7303 vp_p.n23389 vp_p.n23386 14.806
R7304 vp_p.n24811 vp_p.n24808 14.806
R7305 vp_p.n26237 vp_p.n26234 14.806
R7306 vp_p.n13757 vp_p.n13754 14.806
R7307 vp_p.n13752 vp_p.n13749 14.806
R7308 vp_p.n12028 vp_p.n12025 14.806
R7309 vp_p.n10590 vp_p.n10587 14.806
R7310 vp_p.n9088 vp_p.n9085 14.806
R7311 vp_p.n349 vp_p.n346 14.806
R7312 vp_p.n1833 vp_p.n1830 14.806
R7313 vp_p.n3258 vp_p.n3255 14.806
R7314 vp_p.n4682 vp_p.n4679 14.806
R7315 vp_p.n6105 vp_p.n6102 14.806
R7316 vp_p.n7527 vp_p.n7524 14.806
R7317 vp_p.n14831 vp_p.n14828 14.806
R7318 vp_p.n16259 vp_p.n16256 14.806
R7319 vp_p.n17686 vp_p.n17683 14.806
R7320 vp_p.n19112 vp_p.n19109 14.806
R7321 vp_p.n20537 vp_p.n20534 14.806
R7322 vp_p.n21961 vp_p.n21958 14.806
R7323 vp_p.n23384 vp_p.n23381 14.806
R7324 vp_p.n24806 vp_p.n24803 14.806
R7325 vp_p.n26232 vp_p.n26229 14.806
R7326 vp_p.n13747 vp_p.n13744 14.806
R7327 vp_p.n13742 vp_p.n13739 14.806
R7328 vp_p.n12023 vp_p.n12020 14.806
R7329 vp_p.n10585 vp_p.n10582 14.806
R7330 vp_p.n9083 vp_p.n9080 14.806
R7331 vp_p.n344 vp_p.n341 14.806
R7332 vp_p.n1828 vp_p.n1825 14.806
R7333 vp_p.n3253 vp_p.n3250 14.806
R7334 vp_p.n4677 vp_p.n4674 14.806
R7335 vp_p.n6100 vp_p.n6097 14.806
R7336 vp_p.n7522 vp_p.n7519 14.806
R7337 vp_p.n14826 vp_p.n14823 14.806
R7338 vp_p.n16254 vp_p.n16251 14.806
R7339 vp_p.n17681 vp_p.n17678 14.806
R7340 vp_p.n19107 vp_p.n19104 14.806
R7341 vp_p.n20532 vp_p.n20529 14.806
R7342 vp_p.n21956 vp_p.n21953 14.806
R7343 vp_p.n23379 vp_p.n23376 14.806
R7344 vp_p.n24801 vp_p.n24798 14.806
R7345 vp_p.n26227 vp_p.n26224 14.806
R7346 vp_p.n13737 vp_p.n13734 14.806
R7347 vp_p.n13732 vp_p.n13729 14.806
R7348 vp_p.n12018 vp_p.n12015 14.806
R7349 vp_p.n10580 vp_p.n10577 14.806
R7350 vp_p.n9078 vp_p.n9075 14.806
R7351 vp_p.n339 vp_p.n336 14.806
R7352 vp_p.n1823 vp_p.n1820 14.806
R7353 vp_p.n3248 vp_p.n3245 14.806
R7354 vp_p.n4672 vp_p.n4669 14.806
R7355 vp_p.n6095 vp_p.n6092 14.806
R7356 vp_p.n7517 vp_p.n7514 14.806
R7357 vp_p.n14821 vp_p.n14818 14.806
R7358 vp_p.n16249 vp_p.n16246 14.806
R7359 vp_p.n17676 vp_p.n17673 14.806
R7360 vp_p.n19102 vp_p.n19099 14.806
R7361 vp_p.n20527 vp_p.n20524 14.806
R7362 vp_p.n21951 vp_p.n21948 14.806
R7363 vp_p.n23374 vp_p.n23371 14.806
R7364 vp_p.n24796 vp_p.n24793 14.806
R7365 vp_p.n26222 vp_p.n26219 14.806
R7366 vp_p.n13727 vp_p.n13724 14.806
R7367 vp_p.n13722 vp_p.n13719 14.806
R7368 vp_p.n12013 vp_p.n12010 14.806
R7369 vp_p.n10575 vp_p.n10572 14.806
R7370 vp_p.n9073 vp_p.n9070 14.806
R7371 vp_p.n334 vp_p.n331 14.806
R7372 vp_p.n1818 vp_p.n1815 14.806
R7373 vp_p.n3243 vp_p.n3240 14.806
R7374 vp_p.n4667 vp_p.n4664 14.806
R7375 vp_p.n6090 vp_p.n6087 14.806
R7376 vp_p.n7512 vp_p.n7509 14.806
R7377 vp_p.n14816 vp_p.n14813 14.806
R7378 vp_p.n16244 vp_p.n16241 14.806
R7379 vp_p.n17671 vp_p.n17668 14.806
R7380 vp_p.n19097 vp_p.n19094 14.806
R7381 vp_p.n20522 vp_p.n20519 14.806
R7382 vp_p.n21946 vp_p.n21943 14.806
R7383 vp_p.n23369 vp_p.n23366 14.806
R7384 vp_p.n24791 vp_p.n24788 14.806
R7385 vp_p.n26217 vp_p.n26214 14.806
R7386 vp_p.n13717 vp_p.n13714 14.806
R7387 vp_p.n13712 vp_p.n13709 14.806
R7388 vp_p.n12008 vp_p.n12005 14.806
R7389 vp_p.n10570 vp_p.n10567 14.806
R7390 vp_p.n9068 vp_p.n9065 14.806
R7391 vp_p.n329 vp_p.n326 14.806
R7392 vp_p.n1813 vp_p.n1810 14.806
R7393 vp_p.n3238 vp_p.n3235 14.806
R7394 vp_p.n4662 vp_p.n4659 14.806
R7395 vp_p.n6085 vp_p.n6082 14.806
R7396 vp_p.n7507 vp_p.n7504 14.806
R7397 vp_p.n14811 vp_p.n14808 14.806
R7398 vp_p.n16239 vp_p.n16236 14.806
R7399 vp_p.n17666 vp_p.n17663 14.806
R7400 vp_p.n19092 vp_p.n19089 14.806
R7401 vp_p.n20517 vp_p.n20514 14.806
R7402 vp_p.n21941 vp_p.n21938 14.806
R7403 vp_p.n23364 vp_p.n23361 14.806
R7404 vp_p.n24786 vp_p.n24783 14.806
R7405 vp_p.n26212 vp_p.n26209 14.806
R7406 vp_p.n13707 vp_p.n13704 14.806
R7407 vp_p.n13702 vp_p.n13699 14.806
R7408 vp_p.n12003 vp_p.n12000 14.806
R7409 vp_p.n10565 vp_p.n10562 14.806
R7410 vp_p.n9063 vp_p.n9060 14.806
R7411 vp_p.n324 vp_p.n321 14.806
R7412 vp_p.n1808 vp_p.n1805 14.806
R7413 vp_p.n3233 vp_p.n3230 14.806
R7414 vp_p.n4657 vp_p.n4654 14.806
R7415 vp_p.n6080 vp_p.n6077 14.806
R7416 vp_p.n7502 vp_p.n7499 14.806
R7417 vp_p.n14806 vp_p.n14803 14.806
R7418 vp_p.n16234 vp_p.n16231 14.806
R7419 vp_p.n17661 vp_p.n17658 14.806
R7420 vp_p.n19087 vp_p.n19084 14.806
R7421 vp_p.n20512 vp_p.n20509 14.806
R7422 vp_p.n21936 vp_p.n21933 14.806
R7423 vp_p.n23359 vp_p.n23356 14.806
R7424 vp_p.n24781 vp_p.n24778 14.806
R7425 vp_p.n26207 vp_p.n26204 14.806
R7426 vp_p.n13697 vp_p.n13694 14.806
R7427 vp_p.n13692 vp_p.n13689 14.806
R7428 vp_p.n11998 vp_p.n11995 14.806
R7429 vp_p.n10560 vp_p.n10557 14.806
R7430 vp_p.n9058 vp_p.n9055 14.806
R7431 vp_p.n319 vp_p.n316 14.806
R7432 vp_p.n1803 vp_p.n1800 14.806
R7433 vp_p.n3228 vp_p.n3225 14.806
R7434 vp_p.n4652 vp_p.n4649 14.806
R7435 vp_p.n6075 vp_p.n6072 14.806
R7436 vp_p.n7497 vp_p.n7494 14.806
R7437 vp_p.n14801 vp_p.n14798 14.806
R7438 vp_p.n16229 vp_p.n16226 14.806
R7439 vp_p.n17656 vp_p.n17653 14.806
R7440 vp_p.n19082 vp_p.n19079 14.806
R7441 vp_p.n20507 vp_p.n20504 14.806
R7442 vp_p.n21931 vp_p.n21928 14.806
R7443 vp_p.n23354 vp_p.n23351 14.806
R7444 vp_p.n24776 vp_p.n24773 14.806
R7445 vp_p.n26202 vp_p.n26199 14.806
R7446 vp_p.n13687 vp_p.n13684 14.806
R7447 vp_p.n13682 vp_p.n13679 14.806
R7448 vp_p.n11993 vp_p.n11990 14.806
R7449 vp_p.n10555 vp_p.n10552 14.806
R7450 vp_p.n9053 vp_p.n9050 14.806
R7451 vp_p.n314 vp_p.n311 14.806
R7452 vp_p.n1798 vp_p.n1795 14.806
R7453 vp_p.n3223 vp_p.n3220 14.806
R7454 vp_p.n4647 vp_p.n4644 14.806
R7455 vp_p.n6070 vp_p.n6067 14.806
R7456 vp_p.n7492 vp_p.n7489 14.806
R7457 vp_p.n14796 vp_p.n14793 14.806
R7458 vp_p.n16224 vp_p.n16221 14.806
R7459 vp_p.n17651 vp_p.n17648 14.806
R7460 vp_p.n19077 vp_p.n19074 14.806
R7461 vp_p.n20502 vp_p.n20499 14.806
R7462 vp_p.n21926 vp_p.n21923 14.806
R7463 vp_p.n23349 vp_p.n23346 14.806
R7464 vp_p.n24771 vp_p.n24768 14.806
R7465 vp_p.n26197 vp_p.n26194 14.806
R7466 vp_p.n13677 vp_p.n13674 14.806
R7467 vp_p.n13672 vp_p.n13669 14.806
R7468 vp_p.n11988 vp_p.n11985 14.806
R7469 vp_p.n10550 vp_p.n10547 14.806
R7470 vp_p.n9048 vp_p.n9045 14.806
R7471 vp_p.n309 vp_p.n306 14.806
R7472 vp_p.n1793 vp_p.n1790 14.806
R7473 vp_p.n3218 vp_p.n3215 14.806
R7474 vp_p.n4642 vp_p.n4639 14.806
R7475 vp_p.n6065 vp_p.n6062 14.806
R7476 vp_p.n7487 vp_p.n7484 14.806
R7477 vp_p.n14791 vp_p.n14788 14.806
R7478 vp_p.n16219 vp_p.n16216 14.806
R7479 vp_p.n17646 vp_p.n17643 14.806
R7480 vp_p.n19072 vp_p.n19069 14.806
R7481 vp_p.n20497 vp_p.n20494 14.806
R7482 vp_p.n21921 vp_p.n21918 14.806
R7483 vp_p.n23344 vp_p.n23341 14.806
R7484 vp_p.n24766 vp_p.n24763 14.806
R7485 vp_p.n26192 vp_p.n26189 14.806
R7486 vp_p.n13667 vp_p.n13664 14.806
R7487 vp_p.n13662 vp_p.n13659 14.806
R7488 vp_p.n11983 vp_p.n11980 14.806
R7489 vp_p.n10545 vp_p.n10542 14.806
R7490 vp_p.n9043 vp_p.n9040 14.806
R7491 vp_p.n304 vp_p.n301 14.806
R7492 vp_p.n1788 vp_p.n1785 14.806
R7493 vp_p.n3213 vp_p.n3210 14.806
R7494 vp_p.n4637 vp_p.n4634 14.806
R7495 vp_p.n6060 vp_p.n6057 14.806
R7496 vp_p.n7482 vp_p.n7479 14.806
R7497 vp_p.n14786 vp_p.n14783 14.806
R7498 vp_p.n16214 vp_p.n16211 14.806
R7499 vp_p.n17641 vp_p.n17638 14.806
R7500 vp_p.n19067 vp_p.n19064 14.806
R7501 vp_p.n20492 vp_p.n20489 14.806
R7502 vp_p.n21916 vp_p.n21913 14.806
R7503 vp_p.n23339 vp_p.n23336 14.806
R7504 vp_p.n24761 vp_p.n24758 14.806
R7505 vp_p.n26187 vp_p.n26184 14.806
R7506 vp_p.n13657 vp_p.n13654 14.806
R7507 vp_p.n13652 vp_p.n13649 14.806
R7508 vp_p.n11978 vp_p.n11975 14.806
R7509 vp_p.n10540 vp_p.n10537 14.806
R7510 vp_p.n9038 vp_p.n9035 14.806
R7511 vp_p.n299 vp_p.n296 14.806
R7512 vp_p.n1783 vp_p.n1780 14.806
R7513 vp_p.n3208 vp_p.n3205 14.806
R7514 vp_p.n4632 vp_p.n4629 14.806
R7515 vp_p.n6055 vp_p.n6052 14.806
R7516 vp_p.n7477 vp_p.n7474 14.806
R7517 vp_p.n14781 vp_p.n14778 14.806
R7518 vp_p.n16209 vp_p.n16206 14.806
R7519 vp_p.n17636 vp_p.n17633 14.806
R7520 vp_p.n19062 vp_p.n19059 14.806
R7521 vp_p.n20487 vp_p.n20484 14.806
R7522 vp_p.n21911 vp_p.n21908 14.806
R7523 vp_p.n23334 vp_p.n23331 14.806
R7524 vp_p.n24756 vp_p.n24753 14.806
R7525 vp_p.n26182 vp_p.n26179 14.806
R7526 vp_p.n13647 vp_p.n13644 14.806
R7527 vp_p.n13642 vp_p.n13639 14.806
R7528 vp_p.n11973 vp_p.n11970 14.806
R7529 vp_p.n10535 vp_p.n10532 14.806
R7530 vp_p.n9033 vp_p.n9030 14.806
R7531 vp_p.n294 vp_p.n291 14.806
R7532 vp_p.n1778 vp_p.n1775 14.806
R7533 vp_p.n3203 vp_p.n3200 14.806
R7534 vp_p.n4627 vp_p.n4624 14.806
R7535 vp_p.n6050 vp_p.n6047 14.806
R7536 vp_p.n7472 vp_p.n7469 14.806
R7537 vp_p.n14776 vp_p.n14773 14.806
R7538 vp_p.n16204 vp_p.n16201 14.806
R7539 vp_p.n17631 vp_p.n17628 14.806
R7540 vp_p.n19057 vp_p.n19054 14.806
R7541 vp_p.n20482 vp_p.n20479 14.806
R7542 vp_p.n21906 vp_p.n21903 14.806
R7543 vp_p.n23329 vp_p.n23326 14.806
R7544 vp_p.n24751 vp_p.n24748 14.806
R7545 vp_p.n26177 vp_p.n26174 14.806
R7546 vp_p.n13637 vp_p.n13634 14.806
R7547 vp_p.n13632 vp_p.n13629 14.806
R7548 vp_p.n11968 vp_p.n11965 14.806
R7549 vp_p.n10530 vp_p.n10527 14.806
R7550 vp_p.n9028 vp_p.n9025 14.806
R7551 vp_p.n289 vp_p.n286 14.806
R7552 vp_p.n1773 vp_p.n1770 14.806
R7553 vp_p.n3198 vp_p.n3195 14.806
R7554 vp_p.n4622 vp_p.n4619 14.806
R7555 vp_p.n6045 vp_p.n6042 14.806
R7556 vp_p.n7467 vp_p.n7464 14.806
R7557 vp_p.n14771 vp_p.n14768 14.806
R7558 vp_p.n16199 vp_p.n16196 14.806
R7559 vp_p.n17626 vp_p.n17623 14.806
R7560 vp_p.n19052 vp_p.n19049 14.806
R7561 vp_p.n20477 vp_p.n20474 14.806
R7562 vp_p.n21901 vp_p.n21898 14.806
R7563 vp_p.n23324 vp_p.n23321 14.806
R7564 vp_p.n24746 vp_p.n24743 14.806
R7565 vp_p.n26172 vp_p.n26169 14.806
R7566 vp_p.n13627 vp_p.n13624 14.806
R7567 vp_p.n13622 vp_p.n13619 14.806
R7568 vp_p.n11963 vp_p.n11960 14.806
R7569 vp_p.n10525 vp_p.n10522 14.806
R7570 vp_p.n9023 vp_p.n9020 14.806
R7571 vp_p.n284 vp_p.n281 14.806
R7572 vp_p.n1768 vp_p.n1765 14.806
R7573 vp_p.n3193 vp_p.n3190 14.806
R7574 vp_p.n4617 vp_p.n4614 14.806
R7575 vp_p.n6040 vp_p.n6037 14.806
R7576 vp_p.n7462 vp_p.n7459 14.806
R7577 vp_p.n14766 vp_p.n14763 14.806
R7578 vp_p.n16194 vp_p.n16191 14.806
R7579 vp_p.n17621 vp_p.n17618 14.806
R7580 vp_p.n19047 vp_p.n19044 14.806
R7581 vp_p.n20472 vp_p.n20469 14.806
R7582 vp_p.n21896 vp_p.n21893 14.806
R7583 vp_p.n23319 vp_p.n23316 14.806
R7584 vp_p.n24741 vp_p.n24738 14.806
R7585 vp_p.n26167 vp_p.n26164 14.806
R7586 vp_p.n13617 vp_p.n13614 14.806
R7587 vp_p.n13612 vp_p.n13609 14.806
R7588 vp_p.n11958 vp_p.n11955 14.806
R7589 vp_p.n10520 vp_p.n10517 14.806
R7590 vp_p.n9018 vp_p.n9015 14.806
R7591 vp_p.n279 vp_p.n276 14.806
R7592 vp_p.n1763 vp_p.n1760 14.806
R7593 vp_p.n3188 vp_p.n3185 14.806
R7594 vp_p.n4612 vp_p.n4609 14.806
R7595 vp_p.n6035 vp_p.n6032 14.806
R7596 vp_p.n7457 vp_p.n7454 14.806
R7597 vp_p.n14761 vp_p.n14758 14.806
R7598 vp_p.n16189 vp_p.n16186 14.806
R7599 vp_p.n17616 vp_p.n17613 14.806
R7600 vp_p.n19042 vp_p.n19039 14.806
R7601 vp_p.n20467 vp_p.n20464 14.806
R7602 vp_p.n21891 vp_p.n21888 14.806
R7603 vp_p.n23314 vp_p.n23311 14.806
R7604 vp_p.n24736 vp_p.n24733 14.806
R7605 vp_p.n26162 vp_p.n26159 14.806
R7606 vp_p.n13607 vp_p.n13604 14.806
R7607 vp_p.n13602 vp_p.n13599 14.806
R7608 vp_p.n11953 vp_p.n11950 14.806
R7609 vp_p.n10515 vp_p.n10512 14.806
R7610 vp_p.n9013 vp_p.n9010 14.806
R7611 vp_p.n274 vp_p.n271 14.806
R7612 vp_p.n1758 vp_p.n1755 14.806
R7613 vp_p.n3183 vp_p.n3180 14.806
R7614 vp_p.n4607 vp_p.n4604 14.806
R7615 vp_p.n6030 vp_p.n6027 14.806
R7616 vp_p.n7452 vp_p.n7449 14.806
R7617 vp_p.n14756 vp_p.n14753 14.806
R7618 vp_p.n16184 vp_p.n16181 14.806
R7619 vp_p.n17611 vp_p.n17608 14.806
R7620 vp_p.n19037 vp_p.n19034 14.806
R7621 vp_p.n20462 vp_p.n20459 14.806
R7622 vp_p.n21886 vp_p.n21883 14.806
R7623 vp_p.n23309 vp_p.n23306 14.806
R7624 vp_p.n24731 vp_p.n24728 14.806
R7625 vp_p.n26157 vp_p.n26154 14.806
R7626 vp_p.n13597 vp_p.n13594 14.806
R7627 vp_p.n13592 vp_p.n13589 14.806
R7628 vp_p.n11948 vp_p.n11945 14.806
R7629 vp_p.n10510 vp_p.n10507 14.806
R7630 vp_p.n9008 vp_p.n9005 14.806
R7631 vp_p.n269 vp_p.n266 14.806
R7632 vp_p.n1753 vp_p.n1750 14.806
R7633 vp_p.n3178 vp_p.n3175 14.806
R7634 vp_p.n4602 vp_p.n4599 14.806
R7635 vp_p.n6025 vp_p.n6022 14.806
R7636 vp_p.n7447 vp_p.n7444 14.806
R7637 vp_p.n14751 vp_p.n14748 14.806
R7638 vp_p.n16179 vp_p.n16176 14.806
R7639 vp_p.n17606 vp_p.n17603 14.806
R7640 vp_p.n19032 vp_p.n19029 14.806
R7641 vp_p.n20457 vp_p.n20454 14.806
R7642 vp_p.n21881 vp_p.n21878 14.806
R7643 vp_p.n23304 vp_p.n23301 14.806
R7644 vp_p.n24726 vp_p.n24723 14.806
R7645 vp_p.n26152 vp_p.n26149 14.806
R7646 vp_p.n13587 vp_p.n13584 14.806
R7647 vp_p.n13582 vp_p.n13579 14.806
R7648 vp_p.n11943 vp_p.n11940 14.806
R7649 vp_p.n10505 vp_p.n10502 14.806
R7650 vp_p.n9003 vp_p.n9000 14.806
R7651 vp_p.n264 vp_p.n261 14.806
R7652 vp_p.n1748 vp_p.n1745 14.806
R7653 vp_p.n3173 vp_p.n3170 14.806
R7654 vp_p.n4597 vp_p.n4594 14.806
R7655 vp_p.n6020 vp_p.n6017 14.806
R7656 vp_p.n7442 vp_p.n7439 14.806
R7657 vp_p.n14746 vp_p.n14743 14.806
R7658 vp_p.n16174 vp_p.n16171 14.806
R7659 vp_p.n17601 vp_p.n17598 14.806
R7660 vp_p.n19027 vp_p.n19024 14.806
R7661 vp_p.n20452 vp_p.n20449 14.806
R7662 vp_p.n21876 vp_p.n21873 14.806
R7663 vp_p.n23299 vp_p.n23296 14.806
R7664 vp_p.n24721 vp_p.n24718 14.806
R7665 vp_p.n26147 vp_p.n26144 14.806
R7666 vp_p.n13577 vp_p.n13574 14.806
R7667 vp_p.n13572 vp_p.n13569 14.806
R7668 vp_p.n11938 vp_p.n11935 14.806
R7669 vp_p.n10500 vp_p.n10497 14.806
R7670 vp_p.n8998 vp_p.n8995 14.806
R7671 vp_p.n259 vp_p.n256 14.806
R7672 vp_p.n1743 vp_p.n1740 14.806
R7673 vp_p.n3168 vp_p.n3165 14.806
R7674 vp_p.n4592 vp_p.n4589 14.806
R7675 vp_p.n6015 vp_p.n6012 14.806
R7676 vp_p.n7437 vp_p.n7434 14.806
R7677 vp_p.n14741 vp_p.n14738 14.806
R7678 vp_p.n16169 vp_p.n16166 14.806
R7679 vp_p.n17596 vp_p.n17593 14.806
R7680 vp_p.n19022 vp_p.n19019 14.806
R7681 vp_p.n20447 vp_p.n20444 14.806
R7682 vp_p.n21871 vp_p.n21868 14.806
R7683 vp_p.n23294 vp_p.n23291 14.806
R7684 vp_p.n24716 vp_p.n24713 14.806
R7685 vp_p.n26142 vp_p.n26139 14.806
R7686 vp_p.n13567 vp_p.n13564 14.806
R7687 vp_p.n13562 vp_p.n13559 14.806
R7688 vp_p.n11933 vp_p.n11930 14.806
R7689 vp_p.n10495 vp_p.n10492 14.806
R7690 vp_p.n8993 vp_p.n8990 14.806
R7691 vp_p.n254 vp_p.n251 14.806
R7692 vp_p.n1738 vp_p.n1735 14.806
R7693 vp_p.n3163 vp_p.n3160 14.806
R7694 vp_p.n4587 vp_p.n4584 14.806
R7695 vp_p.n6010 vp_p.n6007 14.806
R7696 vp_p.n7432 vp_p.n7429 14.806
R7697 vp_p.n14736 vp_p.n14733 14.806
R7698 vp_p.n16164 vp_p.n16161 14.806
R7699 vp_p.n17591 vp_p.n17588 14.806
R7700 vp_p.n19017 vp_p.n19014 14.806
R7701 vp_p.n20442 vp_p.n20439 14.806
R7702 vp_p.n21866 vp_p.n21863 14.806
R7703 vp_p.n23289 vp_p.n23286 14.806
R7704 vp_p.n24711 vp_p.n24708 14.806
R7705 vp_p.n26137 vp_p.n26134 14.806
R7706 vp_p.n13557 vp_p.n13554 14.806
R7707 vp_p.n13552 vp_p.n13549 14.806
R7708 vp_p.n11928 vp_p.n11925 14.806
R7709 vp_p.n10490 vp_p.n10487 14.806
R7710 vp_p.n8988 vp_p.n8985 14.806
R7711 vp_p.n249 vp_p.n246 14.806
R7712 vp_p.n1733 vp_p.n1730 14.806
R7713 vp_p.n3158 vp_p.n3155 14.806
R7714 vp_p.n4582 vp_p.n4579 14.806
R7715 vp_p.n6005 vp_p.n6002 14.806
R7716 vp_p.n7427 vp_p.n7424 14.806
R7717 vp_p.n14731 vp_p.n14728 14.806
R7718 vp_p.n16159 vp_p.n16156 14.806
R7719 vp_p.n17586 vp_p.n17583 14.806
R7720 vp_p.n19012 vp_p.n19009 14.806
R7721 vp_p.n20437 vp_p.n20434 14.806
R7722 vp_p.n21861 vp_p.n21858 14.806
R7723 vp_p.n23284 vp_p.n23281 14.806
R7724 vp_p.n24706 vp_p.n24703 14.806
R7725 vp_p.n26132 vp_p.n26129 14.806
R7726 vp_p.n13547 vp_p.n13544 14.806
R7727 vp_p.n13542 vp_p.n13539 14.806
R7728 vp_p.n11923 vp_p.n11920 14.806
R7729 vp_p.n10485 vp_p.n10482 14.806
R7730 vp_p.n8983 vp_p.n8980 14.806
R7731 vp_p.n244 vp_p.n241 14.806
R7732 vp_p.n1728 vp_p.n1725 14.806
R7733 vp_p.n3153 vp_p.n3150 14.806
R7734 vp_p.n4577 vp_p.n4574 14.806
R7735 vp_p.n6000 vp_p.n5997 14.806
R7736 vp_p.n7422 vp_p.n7419 14.806
R7737 vp_p.n14726 vp_p.n14723 14.806
R7738 vp_p.n16154 vp_p.n16151 14.806
R7739 vp_p.n17581 vp_p.n17578 14.806
R7740 vp_p.n19007 vp_p.n19004 14.806
R7741 vp_p.n20432 vp_p.n20429 14.806
R7742 vp_p.n21856 vp_p.n21853 14.806
R7743 vp_p.n23279 vp_p.n23276 14.806
R7744 vp_p.n24701 vp_p.n24698 14.806
R7745 vp_p.n26127 vp_p.n26124 14.806
R7746 vp_p.n13537 vp_p.n13534 14.806
R7747 vp_p.n13532 vp_p.n13529 14.806
R7748 vp_p.n11918 vp_p.n11915 14.806
R7749 vp_p.n10480 vp_p.n10477 14.806
R7750 vp_p.n8978 vp_p.n8975 14.806
R7751 vp_p.n239 vp_p.n236 14.806
R7752 vp_p.n1723 vp_p.n1720 14.806
R7753 vp_p.n3148 vp_p.n3145 14.806
R7754 vp_p.n4572 vp_p.n4569 14.806
R7755 vp_p.n5995 vp_p.n5992 14.806
R7756 vp_p.n7417 vp_p.n7414 14.806
R7757 vp_p.n14721 vp_p.n14718 14.806
R7758 vp_p.n16149 vp_p.n16146 14.806
R7759 vp_p.n17576 vp_p.n17573 14.806
R7760 vp_p.n19002 vp_p.n18999 14.806
R7761 vp_p.n20427 vp_p.n20424 14.806
R7762 vp_p.n21851 vp_p.n21848 14.806
R7763 vp_p.n23274 vp_p.n23271 14.806
R7764 vp_p.n24696 vp_p.n24693 14.806
R7765 vp_p.n26122 vp_p.n26119 14.806
R7766 vp_p.n13527 vp_p.n13524 14.806
R7767 vp_p.n13522 vp_p.n13519 14.806
R7768 vp_p.n11913 vp_p.n11910 14.806
R7769 vp_p.n10475 vp_p.n10472 14.806
R7770 vp_p.n8973 vp_p.n8970 14.806
R7771 vp_p.n234 vp_p.n231 14.806
R7772 vp_p.n1718 vp_p.n1715 14.806
R7773 vp_p.n3143 vp_p.n3140 14.806
R7774 vp_p.n4567 vp_p.n4564 14.806
R7775 vp_p.n5990 vp_p.n5987 14.806
R7776 vp_p.n7412 vp_p.n7409 14.806
R7777 vp_p.n14716 vp_p.n14713 14.806
R7778 vp_p.n16144 vp_p.n16141 14.806
R7779 vp_p.n17571 vp_p.n17568 14.806
R7780 vp_p.n18997 vp_p.n18994 14.806
R7781 vp_p.n20422 vp_p.n20419 14.806
R7782 vp_p.n21846 vp_p.n21843 14.806
R7783 vp_p.n23269 vp_p.n23266 14.806
R7784 vp_p.n24691 vp_p.n24688 14.806
R7785 vp_p.n26117 vp_p.n26114 14.806
R7786 vp_p.n13517 vp_p.n13514 14.806
R7787 vp_p.n13512 vp_p.n13509 14.806
R7788 vp_p.n11908 vp_p.n11905 14.806
R7789 vp_p.n10470 vp_p.n10467 14.806
R7790 vp_p.n8968 vp_p.n8965 14.806
R7791 vp_p.n229 vp_p.n226 14.806
R7792 vp_p.n1713 vp_p.n1710 14.806
R7793 vp_p.n3138 vp_p.n3135 14.806
R7794 vp_p.n4562 vp_p.n4559 14.806
R7795 vp_p.n5985 vp_p.n5982 14.806
R7796 vp_p.n7407 vp_p.n7404 14.806
R7797 vp_p.n14711 vp_p.n14708 14.806
R7798 vp_p.n16139 vp_p.n16136 14.806
R7799 vp_p.n17566 vp_p.n17563 14.806
R7800 vp_p.n18992 vp_p.n18989 14.806
R7801 vp_p.n20417 vp_p.n20414 14.806
R7802 vp_p.n21841 vp_p.n21838 14.806
R7803 vp_p.n23264 vp_p.n23261 14.806
R7804 vp_p.n24686 vp_p.n24683 14.806
R7805 vp_p.n26112 vp_p.n26109 14.806
R7806 vp_p.n13507 vp_p.n13504 14.806
R7807 vp_p.n13502 vp_p.n13499 14.806
R7808 vp_p.n11903 vp_p.n11900 14.806
R7809 vp_p.n10465 vp_p.n10462 14.806
R7810 vp_p.n8963 vp_p.n8960 14.806
R7811 vp_p.n224 vp_p.n221 14.806
R7812 vp_p.n1708 vp_p.n1705 14.806
R7813 vp_p.n3133 vp_p.n3130 14.806
R7814 vp_p.n4557 vp_p.n4554 14.806
R7815 vp_p.n5980 vp_p.n5977 14.806
R7816 vp_p.n7402 vp_p.n7399 14.806
R7817 vp_p.n14706 vp_p.n14703 14.806
R7818 vp_p.n16134 vp_p.n16131 14.806
R7819 vp_p.n17561 vp_p.n17558 14.806
R7820 vp_p.n18987 vp_p.n18984 14.806
R7821 vp_p.n20412 vp_p.n20409 14.806
R7822 vp_p.n21836 vp_p.n21833 14.806
R7823 vp_p.n23259 vp_p.n23256 14.806
R7824 vp_p.n24681 vp_p.n24678 14.806
R7825 vp_p.n26107 vp_p.n26104 14.806
R7826 vp_p.n13497 vp_p.n13494 14.806
R7827 vp_p.n13492 vp_p.n13489 14.806
R7828 vp_p.n11898 vp_p.n11895 14.806
R7829 vp_p.n10460 vp_p.n10457 14.806
R7830 vp_p.n8958 vp_p.n8955 14.806
R7831 vp_p.n219 vp_p.n216 14.806
R7832 vp_p.n1703 vp_p.n1700 14.806
R7833 vp_p.n3128 vp_p.n3125 14.806
R7834 vp_p.n4552 vp_p.n4549 14.806
R7835 vp_p.n5975 vp_p.n5972 14.806
R7836 vp_p.n7397 vp_p.n7394 14.806
R7837 vp_p.n14701 vp_p.n14698 14.806
R7838 vp_p.n16129 vp_p.n16126 14.806
R7839 vp_p.n17556 vp_p.n17553 14.806
R7840 vp_p.n18982 vp_p.n18979 14.806
R7841 vp_p.n20407 vp_p.n20404 14.806
R7842 vp_p.n21831 vp_p.n21828 14.806
R7843 vp_p.n23254 vp_p.n23251 14.806
R7844 vp_p.n24676 vp_p.n24673 14.806
R7845 vp_p.n26102 vp_p.n26099 14.806
R7846 vp_p.n13487 vp_p.n13484 14.806
R7847 vp_p.n13482 vp_p.n13479 14.806
R7848 vp_p.n11893 vp_p.n11890 14.806
R7849 vp_p.n10455 vp_p.n10452 14.806
R7850 vp_p.n8953 vp_p.n8950 14.806
R7851 vp_p.n214 vp_p.n211 14.806
R7852 vp_p.n1698 vp_p.n1695 14.806
R7853 vp_p.n3123 vp_p.n3120 14.806
R7854 vp_p.n4547 vp_p.n4544 14.806
R7855 vp_p.n5970 vp_p.n5967 14.806
R7856 vp_p.n7392 vp_p.n7389 14.806
R7857 vp_p.n14696 vp_p.n14693 14.806
R7858 vp_p.n16124 vp_p.n16121 14.806
R7859 vp_p.n17551 vp_p.n17548 14.806
R7860 vp_p.n18977 vp_p.n18974 14.806
R7861 vp_p.n20402 vp_p.n20399 14.806
R7862 vp_p.n21826 vp_p.n21823 14.806
R7863 vp_p.n23249 vp_p.n23246 14.806
R7864 vp_p.n24671 vp_p.n24668 14.806
R7865 vp_p.n26097 vp_p.n26094 14.806
R7866 vp_p.n13477 vp_p.n13474 14.806
R7867 vp_p.n13472 vp_p.n13469 14.806
R7868 vp_p.n11888 vp_p.n11885 14.806
R7869 vp_p.n10450 vp_p.n10447 14.806
R7870 vp_p.n8948 vp_p.n8945 14.806
R7871 vp_p.n209 vp_p.n206 14.806
R7872 vp_p.n1693 vp_p.n1690 14.806
R7873 vp_p.n3118 vp_p.n3115 14.806
R7874 vp_p.n4542 vp_p.n4539 14.806
R7875 vp_p.n5965 vp_p.n5962 14.806
R7876 vp_p.n7387 vp_p.n7384 14.806
R7877 vp_p.n14691 vp_p.n14688 14.806
R7878 vp_p.n16119 vp_p.n16116 14.806
R7879 vp_p.n17546 vp_p.n17543 14.806
R7880 vp_p.n18972 vp_p.n18969 14.806
R7881 vp_p.n20397 vp_p.n20394 14.806
R7882 vp_p.n21821 vp_p.n21818 14.806
R7883 vp_p.n23244 vp_p.n23241 14.806
R7884 vp_p.n24666 vp_p.n24663 14.806
R7885 vp_p.n26092 vp_p.n26089 14.806
R7886 vp_p.n13467 vp_p.n13464 14.806
R7887 vp_p.n13462 vp_p.n13459 14.806
R7888 vp_p.n11883 vp_p.n11880 14.806
R7889 vp_p.n10445 vp_p.n10442 14.806
R7890 vp_p.n8943 vp_p.n8940 14.806
R7891 vp_p.n204 vp_p.n201 14.806
R7892 vp_p.n1688 vp_p.n1685 14.806
R7893 vp_p.n3113 vp_p.n3110 14.806
R7894 vp_p.n4537 vp_p.n4534 14.806
R7895 vp_p.n5960 vp_p.n5957 14.806
R7896 vp_p.n7382 vp_p.n7379 14.806
R7897 vp_p.n14686 vp_p.n14683 14.806
R7898 vp_p.n16114 vp_p.n16111 14.806
R7899 vp_p.n17541 vp_p.n17538 14.806
R7900 vp_p.n18967 vp_p.n18964 14.806
R7901 vp_p.n20392 vp_p.n20389 14.806
R7902 vp_p.n21816 vp_p.n21813 14.806
R7903 vp_p.n23239 vp_p.n23236 14.806
R7904 vp_p.n24661 vp_p.n24658 14.806
R7905 vp_p.n26087 vp_p.n26084 14.806
R7906 vp_p.n13457 vp_p.n13454 14.806
R7907 vp_p.n13452 vp_p.n13449 14.806
R7908 vp_p.n11878 vp_p.n11875 14.806
R7909 vp_p.n10440 vp_p.n10437 14.806
R7910 vp_p.n8938 vp_p.n8935 14.806
R7911 vp_p.n199 vp_p.n196 14.806
R7912 vp_p.n1683 vp_p.n1680 14.806
R7913 vp_p.n3108 vp_p.n3105 14.806
R7914 vp_p.n4532 vp_p.n4529 14.806
R7915 vp_p.n5955 vp_p.n5952 14.806
R7916 vp_p.n7377 vp_p.n7374 14.806
R7917 vp_p.n14681 vp_p.n14678 14.806
R7918 vp_p.n16109 vp_p.n16106 14.806
R7919 vp_p.n17536 vp_p.n17533 14.806
R7920 vp_p.n18962 vp_p.n18959 14.806
R7921 vp_p.n20387 vp_p.n20384 14.806
R7922 vp_p.n21811 vp_p.n21808 14.806
R7923 vp_p.n23234 vp_p.n23231 14.806
R7924 vp_p.n24656 vp_p.n24653 14.806
R7925 vp_p.n26082 vp_p.n26079 14.806
R7926 vp_p.n13447 vp_p.n13444 14.806
R7927 vp_p.n13442 vp_p.n13439 14.806
R7928 vp_p.n11873 vp_p.n11870 14.806
R7929 vp_p.n10435 vp_p.n10432 14.806
R7930 vp_p.n8933 vp_p.n8930 14.806
R7931 vp_p.n194 vp_p.n191 14.806
R7932 vp_p.n1678 vp_p.n1675 14.806
R7933 vp_p.n3103 vp_p.n3100 14.806
R7934 vp_p.n4527 vp_p.n4524 14.806
R7935 vp_p.n5950 vp_p.n5947 14.806
R7936 vp_p.n7372 vp_p.n7369 14.806
R7937 vp_p.n14676 vp_p.n14673 14.806
R7938 vp_p.n16104 vp_p.n16101 14.806
R7939 vp_p.n17531 vp_p.n17528 14.806
R7940 vp_p.n18957 vp_p.n18954 14.806
R7941 vp_p.n20382 vp_p.n20379 14.806
R7942 vp_p.n21806 vp_p.n21803 14.806
R7943 vp_p.n23229 vp_p.n23226 14.806
R7944 vp_p.n24651 vp_p.n24648 14.806
R7945 vp_p.n26077 vp_p.n26074 14.806
R7946 vp_p.n13437 vp_p.n13434 14.806
R7947 vp_p.n13432 vp_p.n13429 14.806
R7948 vp_p.n11868 vp_p.n11865 14.806
R7949 vp_p.n10430 vp_p.n10427 14.806
R7950 vp_p.n8928 vp_p.n8925 14.806
R7951 vp_p.n189 vp_p.n186 14.806
R7952 vp_p.n1673 vp_p.n1670 14.806
R7953 vp_p.n3098 vp_p.n3095 14.806
R7954 vp_p.n4522 vp_p.n4519 14.806
R7955 vp_p.n5945 vp_p.n5942 14.806
R7956 vp_p.n7367 vp_p.n7364 14.806
R7957 vp_p.n14671 vp_p.n14668 14.806
R7958 vp_p.n16099 vp_p.n16096 14.806
R7959 vp_p.n17526 vp_p.n17523 14.806
R7960 vp_p.n18952 vp_p.n18949 14.806
R7961 vp_p.n20377 vp_p.n20374 14.806
R7962 vp_p.n21801 vp_p.n21798 14.806
R7963 vp_p.n23224 vp_p.n23221 14.806
R7964 vp_p.n24646 vp_p.n24643 14.806
R7965 vp_p.n26072 vp_p.n26069 14.806
R7966 vp_p.n13427 vp_p.n13424 14.806
R7967 vp_p.n13422 vp_p.n13419 14.806
R7968 vp_p.n11863 vp_p.n11860 14.806
R7969 vp_p.n10425 vp_p.n10422 14.806
R7970 vp_p.n8923 vp_p.n8920 14.806
R7971 vp_p.n184 vp_p.n181 14.806
R7972 vp_p.n1668 vp_p.n1665 14.806
R7973 vp_p.n3093 vp_p.n3090 14.806
R7974 vp_p.n4517 vp_p.n4514 14.806
R7975 vp_p.n5940 vp_p.n5937 14.806
R7976 vp_p.n7362 vp_p.n7359 14.806
R7977 vp_p.n14666 vp_p.n14663 14.806
R7978 vp_p.n16094 vp_p.n16091 14.806
R7979 vp_p.n17521 vp_p.n17518 14.806
R7980 vp_p.n18947 vp_p.n18944 14.806
R7981 vp_p.n20372 vp_p.n20369 14.806
R7982 vp_p.n21796 vp_p.n21793 14.806
R7983 vp_p.n23219 vp_p.n23216 14.806
R7984 vp_p.n24641 vp_p.n24638 14.806
R7985 vp_p.n26067 vp_p.n26064 14.806
R7986 vp_p.n13417 vp_p.n13414 14.806
R7987 vp_p.n13412 vp_p.n13409 14.806
R7988 vp_p.n11858 vp_p.n11855 14.806
R7989 vp_p.n10420 vp_p.n10417 14.806
R7990 vp_p.n8918 vp_p.n8915 14.806
R7991 vp_p.n179 vp_p.n176 14.806
R7992 vp_p.n1663 vp_p.n1660 14.806
R7993 vp_p.n3088 vp_p.n3085 14.806
R7994 vp_p.n4512 vp_p.n4509 14.806
R7995 vp_p.n5935 vp_p.n5932 14.806
R7996 vp_p.n7357 vp_p.n7354 14.806
R7997 vp_p.n14661 vp_p.n14658 14.806
R7998 vp_p.n16089 vp_p.n16086 14.806
R7999 vp_p.n17516 vp_p.n17513 14.806
R8000 vp_p.n18942 vp_p.n18939 14.806
R8001 vp_p.n20367 vp_p.n20364 14.806
R8002 vp_p.n21791 vp_p.n21788 14.806
R8003 vp_p.n23214 vp_p.n23211 14.806
R8004 vp_p.n24636 vp_p.n24633 14.806
R8005 vp_p.n26062 vp_p.n26059 14.806
R8006 vp_p.n13407 vp_p.n13404 14.806
R8007 vp_p.n13402 vp_p.n13399 14.806
R8008 vp_p.n11853 vp_p.n11850 14.806
R8009 vp_p.n10415 vp_p.n10412 14.806
R8010 vp_p.n8913 vp_p.n8910 14.806
R8011 vp_p.n174 vp_p.n171 14.806
R8012 vp_p.n1658 vp_p.n1655 14.806
R8013 vp_p.n3083 vp_p.n3080 14.806
R8014 vp_p.n4507 vp_p.n4504 14.806
R8015 vp_p.n5930 vp_p.n5927 14.806
R8016 vp_p.n7352 vp_p.n7349 14.806
R8017 vp_p.n14656 vp_p.n14653 14.806
R8018 vp_p.n16084 vp_p.n16081 14.806
R8019 vp_p.n17511 vp_p.n17508 14.806
R8020 vp_p.n18937 vp_p.n18934 14.806
R8021 vp_p.n20362 vp_p.n20359 14.806
R8022 vp_p.n21786 vp_p.n21783 14.806
R8023 vp_p.n23209 vp_p.n23206 14.806
R8024 vp_p.n24631 vp_p.n24628 14.806
R8025 vp_p.n26057 vp_p.n26054 14.806
R8026 vp_p.n13397 vp_p.n13394 14.806
R8027 vp_p.n13392 vp_p.n13389 14.806
R8028 vp_p.n11848 vp_p.n11845 14.806
R8029 vp_p.n10410 vp_p.n10407 14.806
R8030 vp_p.n8908 vp_p.n8905 14.806
R8031 vp_p.n169 vp_p.n166 14.806
R8032 vp_p.n1653 vp_p.n1650 14.806
R8033 vp_p.n3078 vp_p.n3075 14.806
R8034 vp_p.n4502 vp_p.n4499 14.806
R8035 vp_p.n5925 vp_p.n5922 14.806
R8036 vp_p.n7347 vp_p.n7344 14.806
R8037 vp_p.n14651 vp_p.n14648 14.806
R8038 vp_p.n16079 vp_p.n16076 14.806
R8039 vp_p.n17506 vp_p.n17503 14.806
R8040 vp_p.n18932 vp_p.n18929 14.806
R8041 vp_p.n20357 vp_p.n20354 14.806
R8042 vp_p.n21781 vp_p.n21778 14.806
R8043 vp_p.n23204 vp_p.n23201 14.806
R8044 vp_p.n24626 vp_p.n24623 14.806
R8045 vp_p.n26052 vp_p.n26049 14.806
R8046 vp_p.n13387 vp_p.n13384 14.806
R8047 vp_p.n13382 vp_p.n13379 14.806
R8048 vp_p.n11843 vp_p.n11840 14.806
R8049 vp_p.n10405 vp_p.n10402 14.806
R8050 vp_p.n8903 vp_p.n8900 14.806
R8051 vp_p.n164 vp_p.n161 14.806
R8052 vp_p.n1648 vp_p.n1645 14.806
R8053 vp_p.n3073 vp_p.n3070 14.806
R8054 vp_p.n4497 vp_p.n4494 14.806
R8055 vp_p.n5920 vp_p.n5917 14.806
R8056 vp_p.n7342 vp_p.n7339 14.806
R8057 vp_p.n14646 vp_p.n14643 14.806
R8058 vp_p.n16074 vp_p.n16071 14.806
R8059 vp_p.n17501 vp_p.n17498 14.806
R8060 vp_p.n18927 vp_p.n18924 14.806
R8061 vp_p.n20352 vp_p.n20349 14.806
R8062 vp_p.n21776 vp_p.n21773 14.806
R8063 vp_p.n23199 vp_p.n23196 14.806
R8064 vp_p.n24621 vp_p.n24618 14.806
R8065 vp_p.n26047 vp_p.n26044 14.806
R8066 vp_p.n13377 vp_p.n13374 14.806
R8067 vp_p.n13372 vp_p.n13369 14.806
R8068 vp_p.n11838 vp_p.n11835 14.806
R8069 vp_p.n10400 vp_p.n10397 14.806
R8070 vp_p.n8898 vp_p.n8895 14.806
R8071 vp_p.n159 vp_p.n156 14.806
R8072 vp_p.n1643 vp_p.n1640 14.806
R8073 vp_p.n3068 vp_p.n3065 14.806
R8074 vp_p.n4492 vp_p.n4489 14.806
R8075 vp_p.n5915 vp_p.n5912 14.806
R8076 vp_p.n7337 vp_p.n7334 14.806
R8077 vp_p.n14641 vp_p.n14638 14.806
R8078 vp_p.n16069 vp_p.n16066 14.806
R8079 vp_p.n17496 vp_p.n17493 14.806
R8080 vp_p.n18922 vp_p.n18919 14.806
R8081 vp_p.n20347 vp_p.n20344 14.806
R8082 vp_p.n21771 vp_p.n21768 14.806
R8083 vp_p.n23194 vp_p.n23191 14.806
R8084 vp_p.n24616 vp_p.n24613 14.806
R8085 vp_p.n26042 vp_p.n26039 14.806
R8086 vp_p.n13367 vp_p.n13364 14.806
R8087 vp_p.n13362 vp_p.n13359 14.806
R8088 vp_p.n11833 vp_p.n11830 14.806
R8089 vp_p.n10395 vp_p.n10392 14.806
R8090 vp_p.n8893 vp_p.n8890 14.806
R8091 vp_p.n154 vp_p.n151 14.806
R8092 vp_p.n1638 vp_p.n1635 14.806
R8093 vp_p.n3063 vp_p.n3060 14.806
R8094 vp_p.n4487 vp_p.n4484 14.806
R8095 vp_p.n5910 vp_p.n5907 14.806
R8096 vp_p.n7332 vp_p.n7329 14.806
R8097 vp_p.n14636 vp_p.n14633 14.806
R8098 vp_p.n16064 vp_p.n16061 14.806
R8099 vp_p.n17491 vp_p.n17488 14.806
R8100 vp_p.n18917 vp_p.n18914 14.806
R8101 vp_p.n20342 vp_p.n20339 14.806
R8102 vp_p.n21766 vp_p.n21763 14.806
R8103 vp_p.n23189 vp_p.n23186 14.806
R8104 vp_p.n24611 vp_p.n24608 14.806
R8105 vp_p.n26037 vp_p.n26034 14.806
R8106 vp_p.n13357 vp_p.n13354 14.806
R8107 vp_p.n13352 vp_p.n13349 14.806
R8108 vp_p.n11828 vp_p.n11825 14.806
R8109 vp_p.n10390 vp_p.n10387 14.806
R8110 vp_p.n8888 vp_p.n8885 14.806
R8111 vp_p.n149 vp_p.n146 14.806
R8112 vp_p.n1633 vp_p.n1630 14.806
R8113 vp_p.n3058 vp_p.n3055 14.806
R8114 vp_p.n4482 vp_p.n4479 14.806
R8115 vp_p.n5905 vp_p.n5902 14.806
R8116 vp_p.n7327 vp_p.n7324 14.806
R8117 vp_p.n14631 vp_p.n14628 14.806
R8118 vp_p.n16059 vp_p.n16056 14.806
R8119 vp_p.n17486 vp_p.n17483 14.806
R8120 vp_p.n18912 vp_p.n18909 14.806
R8121 vp_p.n20337 vp_p.n20334 14.806
R8122 vp_p.n21761 vp_p.n21758 14.806
R8123 vp_p.n23184 vp_p.n23181 14.806
R8124 vp_p.n24606 vp_p.n24603 14.806
R8125 vp_p.n26032 vp_p.n26029 14.806
R8126 vp_p.n13347 vp_p.n13344 14.806
R8127 vp_p.n13342 vp_p.n13339 14.806
R8128 vp_p.n11823 vp_p.n11820 14.806
R8129 vp_p.n10385 vp_p.n10382 14.806
R8130 vp_p.n8883 vp_p.n8880 14.806
R8131 vp_p.n144 vp_p.n141 14.806
R8132 vp_p.n1628 vp_p.n1625 14.806
R8133 vp_p.n3053 vp_p.n3050 14.806
R8134 vp_p.n4477 vp_p.n4474 14.806
R8135 vp_p.n5900 vp_p.n5897 14.806
R8136 vp_p.n7322 vp_p.n7319 14.806
R8137 vp_p.n14626 vp_p.n14623 14.806
R8138 vp_p.n16054 vp_p.n16051 14.806
R8139 vp_p.n17481 vp_p.n17478 14.806
R8140 vp_p.n18907 vp_p.n18904 14.806
R8141 vp_p.n20332 vp_p.n20329 14.806
R8142 vp_p.n21756 vp_p.n21753 14.806
R8143 vp_p.n23179 vp_p.n23176 14.806
R8144 vp_p.n24601 vp_p.n24598 14.806
R8145 vp_p.n26027 vp_p.n26024 14.806
R8146 vp_p.n13337 vp_p.n13334 14.806
R8147 vp_p.n13332 vp_p.n13329 14.806
R8148 vp_p.n11818 vp_p.n11815 14.806
R8149 vp_p.n10380 vp_p.n10377 14.806
R8150 vp_p.n8878 vp_p.n8875 14.806
R8151 vp_p.n139 vp_p.n136 14.806
R8152 vp_p.n1623 vp_p.n1620 14.806
R8153 vp_p.n3048 vp_p.n3045 14.806
R8154 vp_p.n4472 vp_p.n4469 14.806
R8155 vp_p.n5895 vp_p.n5892 14.806
R8156 vp_p.n7317 vp_p.n7314 14.806
R8157 vp_p.n14621 vp_p.n14618 14.806
R8158 vp_p.n16049 vp_p.n16046 14.806
R8159 vp_p.n17476 vp_p.n17473 14.806
R8160 vp_p.n18902 vp_p.n18899 14.806
R8161 vp_p.n20327 vp_p.n20324 14.806
R8162 vp_p.n21751 vp_p.n21748 14.806
R8163 vp_p.n23174 vp_p.n23171 14.806
R8164 vp_p.n24596 vp_p.n24593 14.806
R8165 vp_p.n26022 vp_p.n26019 14.806
R8166 vp_p.n13327 vp_p.n13324 14.806
R8167 vp_p.n13322 vp_p.n13319 14.806
R8168 vp_p.n11813 vp_p.n11810 14.806
R8169 vp_p.n10375 vp_p.n10372 14.806
R8170 vp_p.n8873 vp_p.n8870 14.806
R8171 vp_p.n134 vp_p.n131 14.806
R8172 vp_p.n1618 vp_p.n1615 14.806
R8173 vp_p.n3043 vp_p.n3040 14.806
R8174 vp_p.n4467 vp_p.n4464 14.806
R8175 vp_p.n5890 vp_p.n5887 14.806
R8176 vp_p.n7312 vp_p.n7309 14.806
R8177 vp_p.n14616 vp_p.n14613 14.806
R8178 vp_p.n16044 vp_p.n16041 14.806
R8179 vp_p.n17471 vp_p.n17468 14.806
R8180 vp_p.n18897 vp_p.n18894 14.806
R8181 vp_p.n20322 vp_p.n20319 14.806
R8182 vp_p.n21746 vp_p.n21743 14.806
R8183 vp_p.n23169 vp_p.n23166 14.806
R8184 vp_p.n24591 vp_p.n24588 14.806
R8185 vp_p.n26017 vp_p.n26014 14.806
R8186 vp_p.n13317 vp_p.n13314 14.806
R8187 vp_p.n13312 vp_p.n13309 14.806
R8188 vp_p.n11808 vp_p.n11805 14.806
R8189 vp_p.n10370 vp_p.n10367 14.806
R8190 vp_p.n8868 vp_p.n8865 14.806
R8191 vp_p.n129 vp_p.n126 14.806
R8192 vp_p.n1613 vp_p.n1610 14.806
R8193 vp_p.n3038 vp_p.n3035 14.806
R8194 vp_p.n4462 vp_p.n4459 14.806
R8195 vp_p.n5885 vp_p.n5882 14.806
R8196 vp_p.n7307 vp_p.n7304 14.806
R8197 vp_p.n14611 vp_p.n14608 14.806
R8198 vp_p.n16039 vp_p.n16036 14.806
R8199 vp_p.n17466 vp_p.n17463 14.806
R8200 vp_p.n18892 vp_p.n18889 14.806
R8201 vp_p.n20317 vp_p.n20314 14.806
R8202 vp_p.n21741 vp_p.n21738 14.806
R8203 vp_p.n23164 vp_p.n23161 14.806
R8204 vp_p.n24586 vp_p.n24583 14.806
R8205 vp_p.n26012 vp_p.n26009 14.806
R8206 vp_p.n13307 vp_p.n13304 14.806
R8207 vp_p.n13302 vp_p.n13299 14.806
R8208 vp_p.n11803 vp_p.n11800 14.806
R8209 vp_p.n10365 vp_p.n10362 14.806
R8210 vp_p.n8863 vp_p.n8860 14.806
R8211 vp_p.n124 vp_p.n121 14.806
R8212 vp_p.n1608 vp_p.n1605 14.806
R8213 vp_p.n3033 vp_p.n3030 14.806
R8214 vp_p.n4457 vp_p.n4454 14.806
R8215 vp_p.n5880 vp_p.n5877 14.806
R8216 vp_p.n7302 vp_p.n7299 14.806
R8217 vp_p.n14606 vp_p.n14603 14.806
R8218 vp_p.n16034 vp_p.n16031 14.806
R8219 vp_p.n17461 vp_p.n17458 14.806
R8220 vp_p.n18887 vp_p.n18884 14.806
R8221 vp_p.n20312 vp_p.n20309 14.806
R8222 vp_p.n21736 vp_p.n21733 14.806
R8223 vp_p.n23159 vp_p.n23156 14.806
R8224 vp_p.n24581 vp_p.n24578 14.806
R8225 vp_p.n26007 vp_p.n26004 14.806
R8226 vp_p.n13297 vp_p.n13294 14.806
R8227 vp_p.n13292 vp_p.n13289 14.806
R8228 vp_p.n11798 vp_p.n11795 14.806
R8229 vp_p.n10360 vp_p.n10357 14.806
R8230 vp_p.n8858 vp_p.n8855 14.806
R8231 vp_p.n119 vp_p.n116 14.806
R8232 vp_p.n1603 vp_p.n1600 14.806
R8233 vp_p.n3028 vp_p.n3025 14.806
R8234 vp_p.n4452 vp_p.n4449 14.806
R8235 vp_p.n5875 vp_p.n5872 14.806
R8236 vp_p.n7297 vp_p.n7294 14.806
R8237 vp_p.n14601 vp_p.n14598 14.806
R8238 vp_p.n16029 vp_p.n16026 14.806
R8239 vp_p.n17456 vp_p.n17453 14.806
R8240 vp_p.n18882 vp_p.n18879 14.806
R8241 vp_p.n20307 vp_p.n20304 14.806
R8242 vp_p.n21731 vp_p.n21728 14.806
R8243 vp_p.n23154 vp_p.n23151 14.806
R8244 vp_p.n24576 vp_p.n24573 14.806
R8245 vp_p.n26002 vp_p.n25999 14.806
R8246 vp_p.n13287 vp_p.n13284 14.806
R8247 vp_p.n13282 vp_p.n13279 14.806
R8248 vp_p.n11793 vp_p.n11790 14.806
R8249 vp_p.n10355 vp_p.n10352 14.806
R8250 vp_p.n8853 vp_p.n8850 14.806
R8251 vp_p.n114 vp_p.n111 14.806
R8252 vp_p.n1598 vp_p.n1595 14.806
R8253 vp_p.n3023 vp_p.n3020 14.806
R8254 vp_p.n4447 vp_p.n4444 14.806
R8255 vp_p.n5870 vp_p.n5867 14.806
R8256 vp_p.n7292 vp_p.n7289 14.806
R8257 vp_p.n14596 vp_p.n14593 14.806
R8258 vp_p.n16024 vp_p.n16021 14.806
R8259 vp_p.n17451 vp_p.n17448 14.806
R8260 vp_p.n18877 vp_p.n18874 14.806
R8261 vp_p.n20302 vp_p.n20299 14.806
R8262 vp_p.n21726 vp_p.n21723 14.806
R8263 vp_p.n23149 vp_p.n23146 14.806
R8264 vp_p.n24571 vp_p.n24568 14.806
R8265 vp_p.n25997 vp_p.n25994 14.806
R8266 vp_p.n13277 vp_p.n13274 14.806
R8267 vp_p.n13272 vp_p.n13269 14.806
R8268 vp_p.n11788 vp_p.n11785 14.806
R8269 vp_p.n10350 vp_p.n10347 14.806
R8270 vp_p.n8848 vp_p.n8845 14.806
R8271 vp_p.n109 vp_p.n106 14.806
R8272 vp_p.n1593 vp_p.n1590 14.806
R8273 vp_p.n3018 vp_p.n3015 14.806
R8274 vp_p.n4442 vp_p.n4439 14.806
R8275 vp_p.n5865 vp_p.n5862 14.806
R8276 vp_p.n7287 vp_p.n7284 14.806
R8277 vp_p.n14591 vp_p.n14588 14.806
R8278 vp_p.n16019 vp_p.n16016 14.806
R8279 vp_p.n17446 vp_p.n17443 14.806
R8280 vp_p.n18872 vp_p.n18869 14.806
R8281 vp_p.n20297 vp_p.n20294 14.806
R8282 vp_p.n21721 vp_p.n21718 14.806
R8283 vp_p.n23144 vp_p.n23141 14.806
R8284 vp_p.n24566 vp_p.n24563 14.806
R8285 vp_p.n25992 vp_p.n25989 14.806
R8286 vp_p.n13267 vp_p.n13264 14.806
R8287 vp_p.n13262 vp_p.n13259 14.806
R8288 vp_p.n11783 vp_p.n11780 14.806
R8289 vp_p.n10345 vp_p.n10342 14.806
R8290 vp_p.n8843 vp_p.n8840 14.806
R8291 vp_p.n104 vp_p.n101 14.806
R8292 vp_p.n1588 vp_p.n1585 14.806
R8293 vp_p.n3013 vp_p.n3010 14.806
R8294 vp_p.n4437 vp_p.n4434 14.806
R8295 vp_p.n5860 vp_p.n5857 14.806
R8296 vp_p.n7282 vp_p.n7279 14.806
R8297 vp_p.n14586 vp_p.n14583 14.806
R8298 vp_p.n16014 vp_p.n16011 14.806
R8299 vp_p.n17441 vp_p.n17438 14.806
R8300 vp_p.n18867 vp_p.n18864 14.806
R8301 vp_p.n20292 vp_p.n20289 14.806
R8302 vp_p.n21716 vp_p.n21713 14.806
R8303 vp_p.n23139 vp_p.n23136 14.806
R8304 vp_p.n24561 vp_p.n24558 14.806
R8305 vp_p.n25987 vp_p.n25984 14.806
R8306 vp_p.n13257 vp_p.n13254 14.806
R8307 vp_p.n13252 vp_p.n13249 14.806
R8308 vp_p.n11778 vp_p.n11775 14.806
R8309 vp_p.n10340 vp_p.n10337 14.806
R8310 vp_p.n8838 vp_p.n8835 14.806
R8311 vp_p.n99 vp_p.n96 14.806
R8312 vp_p.n1583 vp_p.n1580 14.806
R8313 vp_p.n3008 vp_p.n3005 14.806
R8314 vp_p.n4432 vp_p.n4429 14.806
R8315 vp_p.n5855 vp_p.n5852 14.806
R8316 vp_p.n7277 vp_p.n7274 14.806
R8317 vp_p.n14581 vp_p.n14578 14.806
R8318 vp_p.n16009 vp_p.n16006 14.806
R8319 vp_p.n17436 vp_p.n17433 14.806
R8320 vp_p.n18862 vp_p.n18859 14.806
R8321 vp_p.n20287 vp_p.n20284 14.806
R8322 vp_p.n21711 vp_p.n21708 14.806
R8323 vp_p.n23134 vp_p.n23131 14.806
R8324 vp_p.n24556 vp_p.n24553 14.806
R8325 vp_p.n25982 vp_p.n25979 14.806
R8326 vp_p.n13247 vp_p.n13244 14.806
R8327 vp_p.n13242 vp_p.n13239 14.806
R8328 vp_p.n11773 vp_p.n11770 14.806
R8329 vp_p.n10335 vp_p.n10332 14.806
R8330 vp_p.n8833 vp_p.n8830 14.806
R8331 vp_p.n94 vp_p.n91 14.806
R8332 vp_p.n1578 vp_p.n1575 14.806
R8333 vp_p.n3003 vp_p.n3000 14.806
R8334 vp_p.n4427 vp_p.n4424 14.806
R8335 vp_p.n5850 vp_p.n5847 14.806
R8336 vp_p.n7272 vp_p.n7269 14.806
R8337 vp_p.n14576 vp_p.n14573 14.806
R8338 vp_p.n16004 vp_p.n16001 14.806
R8339 vp_p.n17431 vp_p.n17428 14.806
R8340 vp_p.n18857 vp_p.n18854 14.806
R8341 vp_p.n20282 vp_p.n20279 14.806
R8342 vp_p.n21706 vp_p.n21703 14.806
R8343 vp_p.n23129 vp_p.n23126 14.806
R8344 vp_p.n24551 vp_p.n24548 14.806
R8345 vp_p.n25977 vp_p.n25974 14.806
R8346 vp_p.n13237 vp_p.n13234 14.806
R8347 vp_p.n13232 vp_p.n13229 14.806
R8348 vp_p.n11768 vp_p.n11765 14.806
R8349 vp_p.n10330 vp_p.n10327 14.806
R8350 vp_p.n8828 vp_p.n8825 14.806
R8351 vp_p.n89 vp_p.n86 14.806
R8352 vp_p.n1573 vp_p.n1570 14.806
R8353 vp_p.n2998 vp_p.n2995 14.806
R8354 vp_p.n4422 vp_p.n4419 14.806
R8355 vp_p.n5845 vp_p.n5842 14.806
R8356 vp_p.n7267 vp_p.n7264 14.806
R8357 vp_p.n14571 vp_p.n14568 14.806
R8358 vp_p.n15999 vp_p.n15996 14.806
R8359 vp_p.n17426 vp_p.n17423 14.806
R8360 vp_p.n18852 vp_p.n18849 14.806
R8361 vp_p.n20277 vp_p.n20274 14.806
R8362 vp_p.n21701 vp_p.n21698 14.806
R8363 vp_p.n23124 vp_p.n23121 14.806
R8364 vp_p.n24546 vp_p.n24543 14.806
R8365 vp_p.n25972 vp_p.n25969 14.806
R8366 vp_p.n13227 vp_p.n13224 14.806
R8367 vp_p.n13222 vp_p.n13219 14.806
R8368 vp_p.n11763 vp_p.n11760 14.806
R8369 vp_p.n10325 vp_p.n10322 14.806
R8370 vp_p.n8823 vp_p.n8820 14.806
R8371 vp_p.n84 vp_p.n81 14.806
R8372 vp_p.n1568 vp_p.n1565 14.806
R8373 vp_p.n2993 vp_p.n2990 14.806
R8374 vp_p.n4417 vp_p.n4414 14.806
R8375 vp_p.n5840 vp_p.n5837 14.806
R8376 vp_p.n7262 vp_p.n7259 14.806
R8377 vp_p.n14566 vp_p.n14563 14.806
R8378 vp_p.n15994 vp_p.n15991 14.806
R8379 vp_p.n17421 vp_p.n17418 14.806
R8380 vp_p.n18847 vp_p.n18844 14.806
R8381 vp_p.n20272 vp_p.n20269 14.806
R8382 vp_p.n21696 vp_p.n21693 14.806
R8383 vp_p.n23119 vp_p.n23116 14.806
R8384 vp_p.n24541 vp_p.n24538 14.806
R8385 vp_p.n25967 vp_p.n25964 14.806
R8386 vp_p.n13217 vp_p.n13214 14.806
R8387 vp_p.n13212 vp_p.n13209 14.806
R8388 vp_p.n11758 vp_p.n11755 14.806
R8389 vp_p.n10320 vp_p.n10317 14.806
R8390 vp_p.n8818 vp_p.n8815 14.806
R8391 vp_p.n79 vp_p.n76 14.806
R8392 vp_p.n1563 vp_p.n1560 14.806
R8393 vp_p.n2988 vp_p.n2985 14.806
R8394 vp_p.n4412 vp_p.n4409 14.806
R8395 vp_p.n5835 vp_p.n5832 14.806
R8396 vp_p.n7257 vp_p.n7254 14.806
R8397 vp_p.n14561 vp_p.n14558 14.806
R8398 vp_p.n15989 vp_p.n15986 14.806
R8399 vp_p.n17416 vp_p.n17413 14.806
R8400 vp_p.n18842 vp_p.n18839 14.806
R8401 vp_p.n20267 vp_p.n20264 14.806
R8402 vp_p.n21691 vp_p.n21688 14.806
R8403 vp_p.n23114 vp_p.n23111 14.806
R8404 vp_p.n24536 vp_p.n24533 14.806
R8405 vp_p.n25962 vp_p.n25959 14.806
R8406 vp_p.n13207 vp_p.n13204 14.806
R8407 vp_p.n13202 vp_p.n13199 14.806
R8408 vp_p.n11753 vp_p.n11750 14.806
R8409 vp_p.n10315 vp_p.n10312 14.806
R8410 vp_p.n8813 vp_p.n8810 14.806
R8411 vp_p.n74 vp_p.n71 14.806
R8412 vp_p.n1558 vp_p.n1555 14.806
R8413 vp_p.n2983 vp_p.n2980 14.806
R8414 vp_p.n4407 vp_p.n4404 14.806
R8415 vp_p.n5830 vp_p.n5827 14.806
R8416 vp_p.n7252 vp_p.n7249 14.806
R8417 vp_p.n14556 vp_p.n14553 14.806
R8418 vp_p.n15984 vp_p.n15981 14.806
R8419 vp_p.n17411 vp_p.n17408 14.806
R8420 vp_p.n18837 vp_p.n18834 14.806
R8421 vp_p.n20262 vp_p.n20259 14.806
R8422 vp_p.n21686 vp_p.n21683 14.806
R8423 vp_p.n23109 vp_p.n23106 14.806
R8424 vp_p.n24531 vp_p.n24528 14.806
R8425 vp_p.n25957 vp_p.n25954 14.806
R8426 vp_p.n13197 vp_p.n13194 14.806
R8427 vp_p.n13192 vp_p.n13189 14.806
R8428 vp_p.n11748 vp_p.n11745 14.806
R8429 vp_p.n10310 vp_p.n10307 14.806
R8430 vp_p.n8808 vp_p.n8805 14.806
R8431 vp_p.n69 vp_p.n66 14.806
R8432 vp_p.n1553 vp_p.n1550 14.806
R8433 vp_p.n2978 vp_p.n2975 14.806
R8434 vp_p.n4402 vp_p.n4399 14.806
R8435 vp_p.n5825 vp_p.n5822 14.806
R8436 vp_p.n7247 vp_p.n7244 14.806
R8437 vp_p.n14551 vp_p.n14548 14.806
R8438 vp_p.n15979 vp_p.n15976 14.806
R8439 vp_p.n17406 vp_p.n17403 14.806
R8440 vp_p.n18832 vp_p.n18829 14.806
R8441 vp_p.n20257 vp_p.n20254 14.806
R8442 vp_p.n21681 vp_p.n21678 14.806
R8443 vp_p.n23104 vp_p.n23101 14.806
R8444 vp_p.n24526 vp_p.n24523 14.806
R8445 vp_p.n25952 vp_p.n25949 14.806
R8446 vp_p.n13187 vp_p.n13184 14.806
R8447 vp_p.n13182 vp_p.n13179 14.806
R8448 vp_p.n14546 vp_p.n14543 14.806
R8449 vp_p.n15974 vp_p.n15971 14.806
R8450 vp_p.n17401 vp_p.n17398 14.806
R8451 vp_p.n18827 vp_p.n18824 14.806
R8452 vp_p.n20252 vp_p.n20249 14.806
R8453 vp_p.n21676 vp_p.n21673 14.806
R8454 vp_p.n23099 vp_p.n23096 14.806
R8455 vp_p.n24521 vp_p.n24518 14.806
R8456 vp_p.n25947 vp_p.n25944 14.806
R8457 vp_p.n11743 vp_p.n11740 14.806
R8458 vp_p.n14541 vp_p.n14538 14.806
R8459 vp_p.n15969 vp_p.n15966 14.806
R8460 vp_p.n17396 vp_p.n17393 14.806
R8461 vp_p.n18822 vp_p.n18819 14.806
R8462 vp_p.n20247 vp_p.n20244 14.806
R8463 vp_p.n21671 vp_p.n21668 14.806
R8464 vp_p.n23094 vp_p.n23091 14.806
R8465 vp_p.n24516 vp_p.n24513 14.806
R8466 vp_p.n25942 vp_p.n25939 14.806
R8467 vp_p.n10300 vp_p.n10297 14.806
R8468 vp_p.n15964 vp_p.n15961 14.806
R8469 vp_p.n17391 vp_p.n17388 14.806
R8470 vp_p.n18817 vp_p.n18814 14.806
R8471 vp_p.n20242 vp_p.n20239 14.806
R8472 vp_p.n21666 vp_p.n21663 14.806
R8473 vp_p.n23089 vp_p.n23086 14.806
R8474 vp_p.n24511 vp_p.n24508 14.806
R8475 vp_p.n25937 vp_p.n25934 14.806
R8476 vp_p.n8793 vp_p.n8790 14.806
R8477 vp_p.n17386 vp_p.n17383 14.806
R8478 vp_p.n18812 vp_p.n18809 14.806
R8479 vp_p.n20237 vp_p.n20234 14.806
R8480 vp_p.n21661 vp_p.n21658 14.806
R8481 vp_p.n23084 vp_p.n23081 14.806
R8482 vp_p.n24506 vp_p.n24503 14.806
R8483 vp_p.n25932 vp_p.n25929 14.806
R8484 vp_p.n49 vp_p.n46 14.806
R8485 vp_p.n18807 vp_p.n18804 14.806
R8486 vp_p.n20232 vp_p.n20229 14.806
R8487 vp_p.n21656 vp_p.n21653 14.806
R8488 vp_p.n23079 vp_p.n23076 14.806
R8489 vp_p.n24501 vp_p.n24498 14.806
R8490 vp_p.n25927 vp_p.n25924 14.806
R8491 vp_p.n1528 vp_p.n1525 14.806
R8492 vp_p.n20227 vp_p.n20224 14.806
R8493 vp_p.n21651 vp_p.n21648 14.806
R8494 vp_p.n23074 vp_p.n23071 14.806
R8495 vp_p.n24496 vp_p.n24493 14.806
R8496 vp_p.n25922 vp_p.n25919 14.806
R8497 vp_p.n2948 vp_p.n2945 14.806
R8498 vp_p.n21646 vp_p.n21643 14.806
R8499 vp_p.n23069 vp_p.n23066 14.806
R8500 vp_p.n24491 vp_p.n24488 14.806
R8501 vp_p.n25917 vp_p.n25914 14.806
R8502 vp_p.n4367 vp_p.n4364 14.806
R8503 vp_p.n23064 vp_p.n23061 14.806
R8504 vp_p.n24486 vp_p.n24483 14.806
R8505 vp_p.n25912 vp_p.n25909 14.806
R8506 vp_p.n5785 vp_p.n5782 14.806
R8507 vp_p.n24481 vp_p.n24478 14.806
R8508 vp_p.n25907 vp_p.n25904 14.806
R8509 vp_p.n26277 vp_p.n26274 14.806
R8510 vp_p.n7572 vp_p.n7569 14.806
R8511 vp_p.n24856 vp_p.n24853 14.806
R8512 vp_p.n24851 vp_p.n24848 14.806
R8513 vp_p.n6155 vp_p.n6152 14.806
R8514 vp_p.n6150 vp_p.n6147 14.806
R8515 vp_p.n23434 vp_p.n23431 14.806
R8516 vp_p.n23429 vp_p.n23426 14.806
R8517 vp_p.n4732 vp_p.n4729 14.806
R8518 vp_p.n4727 vp_p.n4724 14.806
R8519 vp_p.n22011 vp_p.n22008 14.806
R8520 vp_p.n22006 vp_p.n22003 14.806
R8521 vp_p.n3308 vp_p.n3305 14.806
R8522 vp_p.n3303 vp_p.n3300 14.806
R8523 vp_p.n20587 vp_p.n20584 14.806
R8524 vp_p.n20582 vp_p.n20579 14.806
R8525 vp_p.n1883 vp_p.n1880 14.806
R8526 vp_p.n1878 vp_p.n1875 14.806
R8527 vp_p.n19162 vp_p.n19159 14.806
R8528 vp_p.n19157 vp_p.n19154 14.806
R8529 vp_p.n399 vp_p.n396 14.806
R8530 vp_p.n394 vp_p.n391 14.806
R8531 vp_p.n17736 vp_p.n17733 14.806
R8532 vp_p.n17731 vp_p.n17728 14.806
R8533 vp_p.n9138 vp_p.n9135 14.806
R8534 vp_p.n9133 vp_p.n9130 14.806
R8535 vp_p.n16309 vp_p.n16306 14.806
R8536 vp_p.n16304 vp_p.n16301 14.806
R8537 vp_p.n10640 vp_p.n10637 14.806
R8538 vp_p.n10635 vp_p.n10632 14.806
R8539 vp_p.n14881 vp_p.n14878 14.806
R8540 vp_p.n14876 vp_p.n14873 14.806
R8541 vp_p.n12078 vp_p.n12075 14.806
R8542 vp_p.n12073 vp_p.n12070 14.806
R8543 vp_p.n13842 vp_p.n13839 14.806
R8544 vp_p.n13837 vp_p.n13834 14.806
R8545 vp_p.n13177 vp_p.n13174 14.806
R8546 vp_p.n13172 vp_p.n13169 14.806
R8547 vp_p.n13167 vp_p.n13164 14.806
R8548 vp_p.n13162 vp_p.n13159 14.806
R8549 vp_p.n13157 vp_p.n13154 14.806
R8550 vp_p.n13152 vp_p.n13149 14.806
R8551 vp_p.n13147 vp_p.n13144 14.806
R8552 vp_p.n13142 vp_p.n13139 14.806
R8553 vp_p.n13137 vp_p.n13134 14.806
R8554 vp_p.n13132 vp_p.n13129 14.806
R8555 vp_p.n13127 vp_p.n13124 14.806
R8556 vp_p.n13122 vp_p.n13119 14.806
R8557 vp_p.n13117 vp_p.n13114 14.806
R8558 vp_p.n13112 vp_p.n13109 14.806
R8559 vp_p.n13107 vp_p.n13104 14.806
R8560 vp_p.n13102 vp_p.n13099 14.806
R8561 vp_p.n11738 vp_p.n11735 14.806
R8562 vp_p.n11733 vp_p.n11730 14.806
R8563 vp_p.n11728 vp_p.n11725 14.806
R8564 vp_p.n11723 vp_p.n11720 14.806
R8565 vp_p.n11718 vp_p.n11715 14.806
R8566 vp_p.n11713 vp_p.n11710 14.806
R8567 vp_p.n11708 vp_p.n11705 14.806
R8568 vp_p.n11703 vp_p.n11700 14.806
R8569 vp_p.n11698 vp_p.n11695 14.806
R8570 vp_p.n11693 vp_p.n11690 14.806
R8571 vp_p.n11688 vp_p.n11685 14.806
R8572 vp_p.n11683 vp_p.n11680 14.806
R8573 vp_p.n11678 vp_p.n11675 14.806
R8574 vp_p.n11673 vp_p.n11670 14.806
R8575 vp_p.n11668 vp_p.n11665 14.806
R8576 vp_p.n14536 vp_p.n14533 14.806
R8577 vp_p.n14531 vp_p.n14528 14.806
R8578 vp_p.n14526 vp_p.n14523 14.806
R8579 vp_p.n14521 vp_p.n14518 14.806
R8580 vp_p.n14516 vp_p.n14513 14.806
R8581 vp_p.n14511 vp_p.n14508 14.806
R8582 vp_p.n14506 vp_p.n14503 14.806
R8583 vp_p.n14501 vp_p.n14498 14.806
R8584 vp_p.n14496 vp_p.n14493 14.806
R8585 vp_p.n14491 vp_p.n14488 14.806
R8586 vp_p.n14486 vp_p.n14483 14.806
R8587 vp_p.n14481 vp_p.n14478 14.806
R8588 vp_p.n14476 vp_p.n14473 14.806
R8589 vp_p.n14471 vp_p.n14468 14.806
R8590 vp_p.n10295 vp_p.n10292 14.806
R8591 vp_p.n10290 vp_p.n10287 14.806
R8592 vp_p.n10285 vp_p.n10282 14.806
R8593 vp_p.n10280 vp_p.n10277 14.806
R8594 vp_p.n10275 vp_p.n10272 14.806
R8595 vp_p.n10270 vp_p.n10267 14.806
R8596 vp_p.n10265 vp_p.n10262 14.806
R8597 vp_p.n10260 vp_p.n10257 14.806
R8598 vp_p.n10255 vp_p.n10252 14.806
R8599 vp_p.n10250 vp_p.n10247 14.806
R8600 vp_p.n10245 vp_p.n10242 14.806
R8601 vp_p.n10240 vp_p.n10237 14.806
R8602 vp_p.n10235 vp_p.n10232 14.806
R8603 vp_p.n15959 vp_p.n15956 14.806
R8604 vp_p.n15954 vp_p.n15951 14.806
R8605 vp_p.n15949 vp_p.n15946 14.806
R8606 vp_p.n15944 vp_p.n15941 14.806
R8607 vp_p.n15939 vp_p.n15936 14.806
R8608 vp_p.n15934 vp_p.n15931 14.806
R8609 vp_p.n15929 vp_p.n15926 14.806
R8610 vp_p.n15924 vp_p.n15921 14.806
R8611 vp_p.n15919 vp_p.n15916 14.806
R8612 vp_p.n15914 vp_p.n15911 14.806
R8613 vp_p.n15909 vp_p.n15906 14.806
R8614 vp_p.n15904 vp_p.n15901 14.806
R8615 vp_p.n8788 vp_p.n8785 14.806
R8616 vp_p.n8783 vp_p.n8780 14.806
R8617 vp_p.n8778 vp_p.n8775 14.806
R8618 vp_p.n8773 vp_p.n8770 14.806
R8619 vp_p.n8768 vp_p.n8765 14.806
R8620 vp_p.n8763 vp_p.n8760 14.806
R8621 vp_p.n8758 vp_p.n8755 14.806
R8622 vp_p.n8753 vp_p.n8750 14.806
R8623 vp_p.n8748 vp_p.n8745 14.806
R8624 vp_p.n8743 vp_p.n8740 14.806
R8625 vp_p.n8738 vp_p.n8735 14.806
R8626 vp_p.n17381 vp_p.n17378 14.806
R8627 vp_p.n17376 vp_p.n17373 14.806
R8628 vp_p.n17371 vp_p.n17368 14.806
R8629 vp_p.n17366 vp_p.n17363 14.806
R8630 vp_p.n17361 vp_p.n17358 14.806
R8631 vp_p.n17356 vp_p.n17353 14.806
R8632 vp_p.n17351 vp_p.n17348 14.806
R8633 vp_p.n17346 vp_p.n17343 14.806
R8634 vp_p.n17341 vp_p.n17338 14.806
R8635 vp_p.n17336 vp_p.n17333 14.806
R8636 vp_p.n44 vp_p.n41 14.806
R8637 vp_p.n39 vp_p.n36 14.806
R8638 vp_p.n34 vp_p.n31 14.806
R8639 vp_p.n29 vp_p.n26 14.806
R8640 vp_p.n24 vp_p.n21 14.806
R8641 vp_p.n19 vp_p.n16 14.806
R8642 vp_p.n14 vp_p.n11 14.806
R8643 vp_p.n9 vp_p.n6 14.806
R8644 vp_p.n4 vp_p.n1 14.806
R8645 vp_p.n18802 vp_p.n18799 14.806
R8646 vp_p.n18797 vp_p.n18794 14.806
R8647 vp_p.n18792 vp_p.n18789 14.806
R8648 vp_p.n18787 vp_p.n18784 14.806
R8649 vp_p.n18782 vp_p.n18779 14.806
R8650 vp_p.n18777 vp_p.n18774 14.806
R8651 vp_p.n18772 vp_p.n18769 14.806
R8652 vp_p.n18767 vp_p.n18764 14.806
R8653 vp_p.n1523 vp_p.n1520 14.806
R8654 vp_p.n1518 vp_p.n1515 14.806
R8655 vp_p.n1513 vp_p.n1510 14.806
R8656 vp_p.n1508 vp_p.n1505 14.806
R8657 vp_p.n1503 vp_p.n1500 14.806
R8658 vp_p.n1498 vp_p.n1495 14.806
R8659 vp_p.n1493 vp_p.n1490 14.806
R8660 vp_p.n20222 vp_p.n20219 14.806
R8661 vp_p.n20217 vp_p.n20214 14.806
R8662 vp_p.n20212 vp_p.n20209 14.806
R8663 vp_p.n20207 vp_p.n20204 14.806
R8664 vp_p.n20202 vp_p.n20199 14.806
R8665 vp_p.n20197 vp_p.n20194 14.806
R8666 vp_p.n2943 vp_p.n2940 14.806
R8667 vp_p.n2938 vp_p.n2935 14.806
R8668 vp_p.n2933 vp_p.n2930 14.806
R8669 vp_p.n2928 vp_p.n2925 14.806
R8670 vp_p.n2923 vp_p.n2920 14.806
R8671 vp_p.n21641 vp_p.n21638 14.806
R8672 vp_p.n21636 vp_p.n21633 14.806
R8673 vp_p.n21631 vp_p.n21628 14.806
R8674 vp_p.n21626 vp_p.n21623 14.806
R8675 vp_p.n4362 vp_p.n4359 14.806
R8676 vp_p.n4357 vp_p.n4354 14.806
R8677 vp_p.n4352 vp_p.n4349 14.806
R8678 vp_p.n23059 vp_p.n23056 14.806
R8679 vp_p.n23054 vp_p.n23051 14.806
R8680 vp_p.n5780 vp_p.n5777 14.806
R8681 vp_p.n8626 vp_p.n8623 14.806
R8682 vp_p.n14383 vp_p.n14382 14.805
R8683 vp_p.n15826 vp_p.n15825 14.805
R8684 vp_p.n17268 vp_p.n17267 14.805
R8685 vp_p.n18709 vp_p.n18708 14.805
R8686 vp_p.n20149 vp_p.n20148 14.805
R8687 vp_p.n21588 vp_p.n21587 14.805
R8688 vp_p.n23026 vp_p.n23025 14.805
R8689 vp_p.n24463 vp_p.n24462 14.805
R8690 vp_p.n25899 vp_p.n25898 14.805
R8691 vp_p.n7584 vp_p.n7583 14.805
R8692 vp_p.n13019 vp_p.n13018 14.805
R8693 vp_p.n11595 vp_p.n11594 14.805
R8694 vp_p.n10172 vp_p.n10171 14.805
R8695 vp_p.n1440 vp_p.n1439 14.805
R8696 vp_p.n2880 vp_p.n2879 14.805
R8697 vp_p.n4319 vp_p.n4318 14.805
R8698 vp_p.n5757 vp_p.n5756 14.805
R8699 vp_p.n7194 vp_p.n7193 14.805
R8700 vp_p.n7204 vp_p.n7203 13.653
R8701 vp_p.n7209 vp_p.n7208 13.653
R8702 vp_p.n5787 vp_p.n5786 13.653
R8703 vp_p.n7214 vp_p.n7213 13.653
R8704 vp_p.n5792 vp_p.n5791 13.653
R8705 vp_p.n4369 vp_p.n4368 13.653
R8706 vp_p.n7219 vp_p.n7218 13.653
R8707 vp_p.n5797 vp_p.n5796 13.653
R8708 vp_p.n4374 vp_p.n4373 13.653
R8709 vp_p.n2950 vp_p.n2949 13.653
R8710 vp_p.n7224 vp_p.n7223 13.653
R8711 vp_p.n5802 vp_p.n5801 13.653
R8712 vp_p.n4379 vp_p.n4378 13.653
R8713 vp_p.n2955 vp_p.n2954 13.653
R8714 vp_p.n1530 vp_p.n1529 13.653
R8715 vp_p.n7229 vp_p.n7228 13.653
R8716 vp_p.n5807 vp_p.n5806 13.653
R8717 vp_p.n4384 vp_p.n4383 13.653
R8718 vp_p.n2960 vp_p.n2959 13.653
R8719 vp_p.n1535 vp_p.n1534 13.653
R8720 vp_p.n51 vp_p.n50 13.653
R8721 vp_p.n7234 vp_p.n7233 13.653
R8722 vp_p.n5812 vp_p.n5811 13.653
R8723 vp_p.n4389 vp_p.n4388 13.653
R8724 vp_p.n2965 vp_p.n2964 13.653
R8725 vp_p.n1540 vp_p.n1539 13.653
R8726 vp_p.n56 vp_p.n55 13.653
R8727 vp_p.n8795 vp_p.n8794 13.653
R8728 vp_p.n7239 vp_p.n7238 13.653
R8729 vp_p.n5817 vp_p.n5816 13.653
R8730 vp_p.n4394 vp_p.n4393 13.653
R8731 vp_p.n2970 vp_p.n2969 13.653
R8732 vp_p.n1545 vp_p.n1544 13.653
R8733 vp_p.n61 vp_p.n60 13.653
R8734 vp_p.n8800 vp_p.n8799 13.653
R8735 vp_p.n10302 vp_p.n10301 13.653
R8736 vp_p.n7593 vp_p.n7592 13.653
R8737 vp_p.n6171 vp_p.n6170 13.653
R8738 vp_p.n4748 vp_p.n4747 13.653
R8739 vp_p.n3324 vp_p.n3323 13.653
R8740 vp_p.n1899 vp_p.n1898 13.653
R8741 vp_p.n473 vp_p.n472 13.653
R8742 vp_p.n9219 vp_p.n9218 13.653
R8743 vp_p.n10656 vp_p.n10655 13.653
R8744 vp_p.n12094 vp_p.n12093 13.653
R8745 vp_p.n26297 vp_p.n26296 13.653
R8746 vp_p.n24872 vp_p.n24871 13.653
R8747 vp_p.n23450 vp_p.n23449 13.653
R8748 vp_p.n22027 vp_p.n22026 13.653
R8749 vp_p.n20603 vp_p.n20602 13.653
R8750 vp_p.n19178 vp_p.n19177 13.653
R8751 vp_p.n17752 vp_p.n17751 13.653
R8752 vp_p.n16325 vp_p.n16324 13.653
R8753 vp_p.n14897 vp_p.n14896 13.653
R8754 vp_p.n13831 vp_p.n13830 13.653
R8755 vp_p.n13829 vp_p.n13828 13.653
R8756 vp_p.n7564 vp_p.n7563 13.653
R8757 vp_p.n6142 vp_p.n6141 13.653
R8758 vp_p.n4719 vp_p.n4718 13.653
R8759 vp_p.n3295 vp_p.n3294 13.653
R8760 vp_p.n1870 vp_p.n1869 13.653
R8761 vp_p.n386 vp_p.n385 13.653
R8762 vp_p.n9125 vp_p.n9124 13.653
R8763 vp_p.n10627 vp_p.n10626 13.653
R8764 vp_p.n12065 vp_p.n12064 13.653
R8765 vp_p.n26269 vp_p.n26268 13.653
R8766 vp_p.n24843 vp_p.n24842 13.653
R8767 vp_p.n23421 vp_p.n23420 13.653
R8768 vp_p.n21998 vp_p.n21997 13.653
R8769 vp_p.n20574 vp_p.n20573 13.653
R8770 vp_p.n19149 vp_p.n19148 13.653
R8771 vp_p.n17723 vp_p.n17722 13.653
R8772 vp_p.n16296 vp_p.n16295 13.653
R8773 vp_p.n14868 vp_p.n14867 13.653
R8774 vp_p.n13824 vp_p.n13823 13.653
R8775 vp_p.n7607 vp_p.n7606 13.653
R8776 vp_p.n6185 vp_p.n6184 13.653
R8777 vp_p.n4762 vp_p.n4761 13.653
R8778 vp_p.n3338 vp_p.n3337 13.653
R8779 vp_p.n1913 vp_p.n1912 13.653
R8780 vp_p.n487 vp_p.n486 13.653
R8781 vp_p.n9233 vp_p.n9232 13.653
R8782 vp_p.n10670 vp_p.n10669 13.653
R8783 vp_p.n12108 vp_p.n12107 13.653
R8784 vp_p.n26311 vp_p.n26310 13.653
R8785 vp_p.n24886 vp_p.n24885 13.653
R8786 vp_p.n23464 vp_p.n23463 13.653
R8787 vp_p.n22041 vp_p.n22040 13.653
R8788 vp_p.n20617 vp_p.n20616 13.653
R8789 vp_p.n19192 vp_p.n19191 13.653
R8790 vp_p.n17766 vp_p.n17765 13.653
R8791 vp_p.n16339 vp_p.n16338 13.653
R8792 vp_p.n14911 vp_p.n14910 13.653
R8793 vp_p.n13821 vp_p.n13820 13.653
R8794 vp_p.n13819 vp_p.n13818 13.653
R8795 vp_p.n7559 vp_p.n7558 13.653
R8796 vp_p.n6137 vp_p.n6136 13.653
R8797 vp_p.n4714 vp_p.n4713 13.653
R8798 vp_p.n3290 vp_p.n3289 13.653
R8799 vp_p.n1865 vp_p.n1864 13.653
R8800 vp_p.n381 vp_p.n380 13.653
R8801 vp_p.n9120 vp_p.n9119 13.653
R8802 vp_p.n10622 vp_p.n10621 13.653
R8803 vp_p.n12060 vp_p.n12059 13.653
R8804 vp_p.n26264 vp_p.n26263 13.653
R8805 vp_p.n24838 vp_p.n24837 13.653
R8806 vp_p.n23416 vp_p.n23415 13.653
R8807 vp_p.n21993 vp_p.n21992 13.653
R8808 vp_p.n20569 vp_p.n20568 13.653
R8809 vp_p.n19144 vp_p.n19143 13.653
R8810 vp_p.n17718 vp_p.n17717 13.653
R8811 vp_p.n16291 vp_p.n16290 13.653
R8812 vp_p.n14863 vp_p.n14862 13.653
R8813 vp_p.n13814 vp_p.n13813 13.653
R8814 vp_p.n7621 vp_p.n7620 13.653
R8815 vp_p.n6199 vp_p.n6198 13.653
R8816 vp_p.n4776 vp_p.n4775 13.653
R8817 vp_p.n3352 vp_p.n3351 13.653
R8818 vp_p.n1927 vp_p.n1926 13.653
R8819 vp_p.n501 vp_p.n500 13.653
R8820 vp_p.n9247 vp_p.n9246 13.653
R8821 vp_p.n10684 vp_p.n10683 13.653
R8822 vp_p.n12122 vp_p.n12121 13.653
R8823 vp_p.n26325 vp_p.n26324 13.653
R8824 vp_p.n24900 vp_p.n24899 13.653
R8825 vp_p.n23478 vp_p.n23477 13.653
R8826 vp_p.n22055 vp_p.n22054 13.653
R8827 vp_p.n20631 vp_p.n20630 13.653
R8828 vp_p.n19206 vp_p.n19205 13.653
R8829 vp_p.n17780 vp_p.n17779 13.653
R8830 vp_p.n16353 vp_p.n16352 13.653
R8831 vp_p.n14925 vp_p.n14924 13.653
R8832 vp_p.n13811 vp_p.n13810 13.653
R8833 vp_p.n13809 vp_p.n13808 13.653
R8834 vp_p.n7554 vp_p.n7553 13.653
R8835 vp_p.n6132 vp_p.n6131 13.653
R8836 vp_p.n4709 vp_p.n4708 13.653
R8837 vp_p.n3285 vp_p.n3284 13.653
R8838 vp_p.n1860 vp_p.n1859 13.653
R8839 vp_p.n376 vp_p.n375 13.653
R8840 vp_p.n9115 vp_p.n9114 13.653
R8841 vp_p.n10617 vp_p.n10616 13.653
R8842 vp_p.n12055 vp_p.n12054 13.653
R8843 vp_p.n26259 vp_p.n26258 13.653
R8844 vp_p.n24833 vp_p.n24832 13.653
R8845 vp_p.n23411 vp_p.n23410 13.653
R8846 vp_p.n21988 vp_p.n21987 13.653
R8847 vp_p.n20564 vp_p.n20563 13.653
R8848 vp_p.n19139 vp_p.n19138 13.653
R8849 vp_p.n17713 vp_p.n17712 13.653
R8850 vp_p.n16286 vp_p.n16285 13.653
R8851 vp_p.n14858 vp_p.n14857 13.653
R8852 vp_p.n13804 vp_p.n13803 13.653
R8853 vp_p.n7635 vp_p.n7634 13.653
R8854 vp_p.n6213 vp_p.n6212 13.653
R8855 vp_p.n4790 vp_p.n4789 13.653
R8856 vp_p.n3366 vp_p.n3365 13.653
R8857 vp_p.n1941 vp_p.n1940 13.653
R8858 vp_p.n515 vp_p.n514 13.653
R8859 vp_p.n9261 vp_p.n9260 13.653
R8860 vp_p.n10698 vp_p.n10697 13.653
R8861 vp_p.n12136 vp_p.n12135 13.653
R8862 vp_p.n26339 vp_p.n26338 13.653
R8863 vp_p.n24914 vp_p.n24913 13.653
R8864 vp_p.n23492 vp_p.n23491 13.653
R8865 vp_p.n22069 vp_p.n22068 13.653
R8866 vp_p.n20645 vp_p.n20644 13.653
R8867 vp_p.n19220 vp_p.n19219 13.653
R8868 vp_p.n17794 vp_p.n17793 13.653
R8869 vp_p.n16367 vp_p.n16366 13.653
R8870 vp_p.n14939 vp_p.n14938 13.653
R8871 vp_p.n13801 vp_p.n13800 13.653
R8872 vp_p.n13799 vp_p.n13798 13.653
R8873 vp_p.n7549 vp_p.n7548 13.653
R8874 vp_p.n6127 vp_p.n6126 13.653
R8875 vp_p.n4704 vp_p.n4703 13.653
R8876 vp_p.n3280 vp_p.n3279 13.653
R8877 vp_p.n1855 vp_p.n1854 13.653
R8878 vp_p.n371 vp_p.n370 13.653
R8879 vp_p.n9110 vp_p.n9109 13.653
R8880 vp_p.n10612 vp_p.n10611 13.653
R8881 vp_p.n12050 vp_p.n12049 13.653
R8882 vp_p.n26254 vp_p.n26253 13.653
R8883 vp_p.n24828 vp_p.n24827 13.653
R8884 vp_p.n23406 vp_p.n23405 13.653
R8885 vp_p.n21983 vp_p.n21982 13.653
R8886 vp_p.n20559 vp_p.n20558 13.653
R8887 vp_p.n19134 vp_p.n19133 13.653
R8888 vp_p.n17708 vp_p.n17707 13.653
R8889 vp_p.n16281 vp_p.n16280 13.653
R8890 vp_p.n14853 vp_p.n14852 13.653
R8891 vp_p.n13794 vp_p.n13793 13.653
R8892 vp_p.n7649 vp_p.n7648 13.653
R8893 vp_p.n6227 vp_p.n6226 13.653
R8894 vp_p.n4804 vp_p.n4803 13.653
R8895 vp_p.n3380 vp_p.n3379 13.653
R8896 vp_p.n1955 vp_p.n1954 13.653
R8897 vp_p.n529 vp_p.n528 13.653
R8898 vp_p.n9275 vp_p.n9274 13.653
R8899 vp_p.n10712 vp_p.n10711 13.653
R8900 vp_p.n12150 vp_p.n12149 13.653
R8901 vp_p.n26353 vp_p.n26352 13.653
R8902 vp_p.n24928 vp_p.n24927 13.653
R8903 vp_p.n23506 vp_p.n23505 13.653
R8904 vp_p.n22083 vp_p.n22082 13.653
R8905 vp_p.n20659 vp_p.n20658 13.653
R8906 vp_p.n19234 vp_p.n19233 13.653
R8907 vp_p.n17808 vp_p.n17807 13.653
R8908 vp_p.n16381 vp_p.n16380 13.653
R8909 vp_p.n14953 vp_p.n14952 13.653
R8910 vp_p.n13791 vp_p.n13790 13.653
R8911 vp_p.n13789 vp_p.n13788 13.653
R8912 vp_p.n7544 vp_p.n7543 13.653
R8913 vp_p.n6122 vp_p.n6121 13.653
R8914 vp_p.n4699 vp_p.n4698 13.653
R8915 vp_p.n3275 vp_p.n3274 13.653
R8916 vp_p.n1850 vp_p.n1849 13.653
R8917 vp_p.n366 vp_p.n365 13.653
R8918 vp_p.n9105 vp_p.n9104 13.653
R8919 vp_p.n10607 vp_p.n10606 13.653
R8920 vp_p.n12045 vp_p.n12044 13.653
R8921 vp_p.n26249 vp_p.n26248 13.653
R8922 vp_p.n24823 vp_p.n24822 13.653
R8923 vp_p.n23401 vp_p.n23400 13.653
R8924 vp_p.n21978 vp_p.n21977 13.653
R8925 vp_p.n20554 vp_p.n20553 13.653
R8926 vp_p.n19129 vp_p.n19128 13.653
R8927 vp_p.n17703 vp_p.n17702 13.653
R8928 vp_p.n16276 vp_p.n16275 13.653
R8929 vp_p.n14848 vp_p.n14847 13.653
R8930 vp_p.n13784 vp_p.n13783 13.653
R8931 vp_p.n7663 vp_p.n7662 13.653
R8932 vp_p.n6241 vp_p.n6240 13.653
R8933 vp_p.n4818 vp_p.n4817 13.653
R8934 vp_p.n3394 vp_p.n3393 13.653
R8935 vp_p.n1969 vp_p.n1968 13.653
R8936 vp_p.n543 vp_p.n542 13.653
R8937 vp_p.n9289 vp_p.n9288 13.653
R8938 vp_p.n10726 vp_p.n10725 13.653
R8939 vp_p.n12164 vp_p.n12163 13.653
R8940 vp_p.n26367 vp_p.n26366 13.653
R8941 vp_p.n24942 vp_p.n24941 13.653
R8942 vp_p.n23520 vp_p.n23519 13.653
R8943 vp_p.n22097 vp_p.n22096 13.653
R8944 vp_p.n20673 vp_p.n20672 13.653
R8945 vp_p.n19248 vp_p.n19247 13.653
R8946 vp_p.n17822 vp_p.n17821 13.653
R8947 vp_p.n16395 vp_p.n16394 13.653
R8948 vp_p.n14967 vp_p.n14966 13.653
R8949 vp_p.n13781 vp_p.n13780 13.653
R8950 vp_p.n13779 vp_p.n13778 13.653
R8951 vp_p.n7539 vp_p.n7538 13.653
R8952 vp_p.n6117 vp_p.n6116 13.653
R8953 vp_p.n4694 vp_p.n4693 13.653
R8954 vp_p.n3270 vp_p.n3269 13.653
R8955 vp_p.n1845 vp_p.n1844 13.653
R8956 vp_p.n361 vp_p.n360 13.653
R8957 vp_p.n9100 vp_p.n9099 13.653
R8958 vp_p.n10602 vp_p.n10601 13.653
R8959 vp_p.n12040 vp_p.n12039 13.653
R8960 vp_p.n26244 vp_p.n26243 13.653
R8961 vp_p.n24818 vp_p.n24817 13.653
R8962 vp_p.n23396 vp_p.n23395 13.653
R8963 vp_p.n21973 vp_p.n21972 13.653
R8964 vp_p.n20549 vp_p.n20548 13.653
R8965 vp_p.n19124 vp_p.n19123 13.653
R8966 vp_p.n17698 vp_p.n17697 13.653
R8967 vp_p.n16271 vp_p.n16270 13.653
R8968 vp_p.n14843 vp_p.n14842 13.653
R8969 vp_p.n13774 vp_p.n13773 13.653
R8970 vp_p.n7677 vp_p.n7676 13.653
R8971 vp_p.n6255 vp_p.n6254 13.653
R8972 vp_p.n4832 vp_p.n4831 13.653
R8973 vp_p.n3408 vp_p.n3407 13.653
R8974 vp_p.n1983 vp_p.n1982 13.653
R8975 vp_p.n557 vp_p.n556 13.653
R8976 vp_p.n9303 vp_p.n9302 13.653
R8977 vp_p.n10740 vp_p.n10739 13.653
R8978 vp_p.n12178 vp_p.n12177 13.653
R8979 vp_p.n26381 vp_p.n26380 13.653
R8980 vp_p.n24956 vp_p.n24955 13.653
R8981 vp_p.n23534 vp_p.n23533 13.653
R8982 vp_p.n22111 vp_p.n22110 13.653
R8983 vp_p.n20687 vp_p.n20686 13.653
R8984 vp_p.n19262 vp_p.n19261 13.653
R8985 vp_p.n17836 vp_p.n17835 13.653
R8986 vp_p.n16409 vp_p.n16408 13.653
R8987 vp_p.n14981 vp_p.n14980 13.653
R8988 vp_p.n13771 vp_p.n13770 13.653
R8989 vp_p.n13769 vp_p.n13768 13.653
R8990 vp_p.n7534 vp_p.n7533 13.653
R8991 vp_p.n6112 vp_p.n6111 13.653
R8992 vp_p.n4689 vp_p.n4688 13.653
R8993 vp_p.n3265 vp_p.n3264 13.653
R8994 vp_p.n1840 vp_p.n1839 13.653
R8995 vp_p.n356 vp_p.n355 13.653
R8996 vp_p.n9095 vp_p.n9094 13.653
R8997 vp_p.n10597 vp_p.n10596 13.653
R8998 vp_p.n12035 vp_p.n12034 13.653
R8999 vp_p.n26239 vp_p.n26238 13.653
R9000 vp_p.n24813 vp_p.n24812 13.653
R9001 vp_p.n23391 vp_p.n23390 13.653
R9002 vp_p.n21968 vp_p.n21967 13.653
R9003 vp_p.n20544 vp_p.n20543 13.653
R9004 vp_p.n19119 vp_p.n19118 13.653
R9005 vp_p.n17693 vp_p.n17692 13.653
R9006 vp_p.n16266 vp_p.n16265 13.653
R9007 vp_p.n14838 vp_p.n14837 13.653
R9008 vp_p.n13764 vp_p.n13763 13.653
R9009 vp_p.n7691 vp_p.n7690 13.653
R9010 vp_p.n6269 vp_p.n6268 13.653
R9011 vp_p.n4846 vp_p.n4845 13.653
R9012 vp_p.n3422 vp_p.n3421 13.653
R9013 vp_p.n1997 vp_p.n1996 13.653
R9014 vp_p.n571 vp_p.n570 13.653
R9015 vp_p.n9317 vp_p.n9316 13.653
R9016 vp_p.n10754 vp_p.n10753 13.653
R9017 vp_p.n12192 vp_p.n12191 13.653
R9018 vp_p.n26395 vp_p.n26394 13.653
R9019 vp_p.n24970 vp_p.n24969 13.653
R9020 vp_p.n23548 vp_p.n23547 13.653
R9021 vp_p.n22125 vp_p.n22124 13.653
R9022 vp_p.n20701 vp_p.n20700 13.653
R9023 vp_p.n19276 vp_p.n19275 13.653
R9024 vp_p.n17850 vp_p.n17849 13.653
R9025 vp_p.n16423 vp_p.n16422 13.653
R9026 vp_p.n14995 vp_p.n14994 13.653
R9027 vp_p.n13761 vp_p.n13760 13.653
R9028 vp_p.n13759 vp_p.n13758 13.653
R9029 vp_p.n7529 vp_p.n7528 13.653
R9030 vp_p.n6107 vp_p.n6106 13.653
R9031 vp_p.n4684 vp_p.n4683 13.653
R9032 vp_p.n3260 vp_p.n3259 13.653
R9033 vp_p.n1835 vp_p.n1834 13.653
R9034 vp_p.n351 vp_p.n350 13.653
R9035 vp_p.n9090 vp_p.n9089 13.653
R9036 vp_p.n10592 vp_p.n10591 13.653
R9037 vp_p.n12030 vp_p.n12029 13.653
R9038 vp_p.n26234 vp_p.n26233 13.653
R9039 vp_p.n24808 vp_p.n24807 13.653
R9040 vp_p.n23386 vp_p.n23385 13.653
R9041 vp_p.n21963 vp_p.n21962 13.653
R9042 vp_p.n20539 vp_p.n20538 13.653
R9043 vp_p.n19114 vp_p.n19113 13.653
R9044 vp_p.n17688 vp_p.n17687 13.653
R9045 vp_p.n16261 vp_p.n16260 13.653
R9046 vp_p.n14833 vp_p.n14832 13.653
R9047 vp_p.n13754 vp_p.n13753 13.653
R9048 vp_p.n7705 vp_p.n7704 13.653
R9049 vp_p.n6283 vp_p.n6282 13.653
R9050 vp_p.n4860 vp_p.n4859 13.653
R9051 vp_p.n3436 vp_p.n3435 13.653
R9052 vp_p.n2011 vp_p.n2010 13.653
R9053 vp_p.n585 vp_p.n584 13.653
R9054 vp_p.n9331 vp_p.n9330 13.653
R9055 vp_p.n10768 vp_p.n10767 13.653
R9056 vp_p.n12206 vp_p.n12205 13.653
R9057 vp_p.n26409 vp_p.n26408 13.653
R9058 vp_p.n24984 vp_p.n24983 13.653
R9059 vp_p.n23562 vp_p.n23561 13.653
R9060 vp_p.n22139 vp_p.n22138 13.653
R9061 vp_p.n20715 vp_p.n20714 13.653
R9062 vp_p.n19290 vp_p.n19289 13.653
R9063 vp_p.n17864 vp_p.n17863 13.653
R9064 vp_p.n16437 vp_p.n16436 13.653
R9065 vp_p.n15009 vp_p.n15008 13.653
R9066 vp_p.n13751 vp_p.n13750 13.653
R9067 vp_p.n13749 vp_p.n13748 13.653
R9068 vp_p.n7524 vp_p.n7523 13.653
R9069 vp_p.n6102 vp_p.n6101 13.653
R9070 vp_p.n4679 vp_p.n4678 13.653
R9071 vp_p.n3255 vp_p.n3254 13.653
R9072 vp_p.n1830 vp_p.n1829 13.653
R9073 vp_p.n346 vp_p.n345 13.653
R9074 vp_p.n9085 vp_p.n9084 13.653
R9075 vp_p.n10587 vp_p.n10586 13.653
R9076 vp_p.n12025 vp_p.n12024 13.653
R9077 vp_p.n26229 vp_p.n26228 13.653
R9078 vp_p.n24803 vp_p.n24802 13.653
R9079 vp_p.n23381 vp_p.n23380 13.653
R9080 vp_p.n21958 vp_p.n21957 13.653
R9081 vp_p.n20534 vp_p.n20533 13.653
R9082 vp_p.n19109 vp_p.n19108 13.653
R9083 vp_p.n17683 vp_p.n17682 13.653
R9084 vp_p.n16256 vp_p.n16255 13.653
R9085 vp_p.n14828 vp_p.n14827 13.653
R9086 vp_p.n13744 vp_p.n13743 13.653
R9087 vp_p.n7719 vp_p.n7718 13.653
R9088 vp_p.n6297 vp_p.n6296 13.653
R9089 vp_p.n4874 vp_p.n4873 13.653
R9090 vp_p.n3450 vp_p.n3449 13.653
R9091 vp_p.n2025 vp_p.n2024 13.653
R9092 vp_p.n599 vp_p.n598 13.653
R9093 vp_p.n9345 vp_p.n9344 13.653
R9094 vp_p.n10782 vp_p.n10781 13.653
R9095 vp_p.n12220 vp_p.n12219 13.653
R9096 vp_p.n26423 vp_p.n26422 13.653
R9097 vp_p.n24998 vp_p.n24997 13.653
R9098 vp_p.n23576 vp_p.n23575 13.653
R9099 vp_p.n22153 vp_p.n22152 13.653
R9100 vp_p.n20729 vp_p.n20728 13.653
R9101 vp_p.n19304 vp_p.n19303 13.653
R9102 vp_p.n17878 vp_p.n17877 13.653
R9103 vp_p.n16451 vp_p.n16450 13.653
R9104 vp_p.n15023 vp_p.n15022 13.653
R9105 vp_p.n13741 vp_p.n13740 13.653
R9106 vp_p.n13739 vp_p.n13738 13.653
R9107 vp_p.n7519 vp_p.n7518 13.653
R9108 vp_p.n6097 vp_p.n6096 13.653
R9109 vp_p.n4674 vp_p.n4673 13.653
R9110 vp_p.n3250 vp_p.n3249 13.653
R9111 vp_p.n1825 vp_p.n1824 13.653
R9112 vp_p.n341 vp_p.n340 13.653
R9113 vp_p.n9080 vp_p.n9079 13.653
R9114 vp_p.n10582 vp_p.n10581 13.653
R9115 vp_p.n12020 vp_p.n12019 13.653
R9116 vp_p.n26224 vp_p.n26223 13.653
R9117 vp_p.n24798 vp_p.n24797 13.653
R9118 vp_p.n23376 vp_p.n23375 13.653
R9119 vp_p.n21953 vp_p.n21952 13.653
R9120 vp_p.n20529 vp_p.n20528 13.653
R9121 vp_p.n19104 vp_p.n19103 13.653
R9122 vp_p.n17678 vp_p.n17677 13.653
R9123 vp_p.n16251 vp_p.n16250 13.653
R9124 vp_p.n14823 vp_p.n14822 13.653
R9125 vp_p.n13734 vp_p.n13733 13.653
R9126 vp_p.n7733 vp_p.n7732 13.653
R9127 vp_p.n6311 vp_p.n6310 13.653
R9128 vp_p.n4888 vp_p.n4887 13.653
R9129 vp_p.n3464 vp_p.n3463 13.653
R9130 vp_p.n2039 vp_p.n2038 13.653
R9131 vp_p.n613 vp_p.n612 13.653
R9132 vp_p.n9359 vp_p.n9358 13.653
R9133 vp_p.n10796 vp_p.n10795 13.653
R9134 vp_p.n12234 vp_p.n12233 13.653
R9135 vp_p.n26437 vp_p.n26436 13.653
R9136 vp_p.n25012 vp_p.n25011 13.653
R9137 vp_p.n23590 vp_p.n23589 13.653
R9138 vp_p.n22167 vp_p.n22166 13.653
R9139 vp_p.n20743 vp_p.n20742 13.653
R9140 vp_p.n19318 vp_p.n19317 13.653
R9141 vp_p.n17892 vp_p.n17891 13.653
R9142 vp_p.n16465 vp_p.n16464 13.653
R9143 vp_p.n15037 vp_p.n15036 13.653
R9144 vp_p.n13731 vp_p.n13730 13.653
R9145 vp_p.n13729 vp_p.n13728 13.653
R9146 vp_p.n7514 vp_p.n7513 13.653
R9147 vp_p.n6092 vp_p.n6091 13.653
R9148 vp_p.n4669 vp_p.n4668 13.653
R9149 vp_p.n3245 vp_p.n3244 13.653
R9150 vp_p.n1820 vp_p.n1819 13.653
R9151 vp_p.n336 vp_p.n335 13.653
R9152 vp_p.n9075 vp_p.n9074 13.653
R9153 vp_p.n10577 vp_p.n10576 13.653
R9154 vp_p.n12015 vp_p.n12014 13.653
R9155 vp_p.n26219 vp_p.n26218 13.653
R9156 vp_p.n24793 vp_p.n24792 13.653
R9157 vp_p.n23371 vp_p.n23370 13.653
R9158 vp_p.n21948 vp_p.n21947 13.653
R9159 vp_p.n20524 vp_p.n20523 13.653
R9160 vp_p.n19099 vp_p.n19098 13.653
R9161 vp_p.n17673 vp_p.n17672 13.653
R9162 vp_p.n16246 vp_p.n16245 13.653
R9163 vp_p.n14818 vp_p.n14817 13.653
R9164 vp_p.n13724 vp_p.n13723 13.653
R9165 vp_p.n7747 vp_p.n7746 13.653
R9166 vp_p.n6325 vp_p.n6324 13.653
R9167 vp_p.n4902 vp_p.n4901 13.653
R9168 vp_p.n3478 vp_p.n3477 13.653
R9169 vp_p.n2053 vp_p.n2052 13.653
R9170 vp_p.n627 vp_p.n626 13.653
R9171 vp_p.n9373 vp_p.n9372 13.653
R9172 vp_p.n10810 vp_p.n10809 13.653
R9173 vp_p.n12248 vp_p.n12247 13.653
R9174 vp_p.n26451 vp_p.n26450 13.653
R9175 vp_p.n25026 vp_p.n25025 13.653
R9176 vp_p.n23604 vp_p.n23603 13.653
R9177 vp_p.n22181 vp_p.n22180 13.653
R9178 vp_p.n20757 vp_p.n20756 13.653
R9179 vp_p.n19332 vp_p.n19331 13.653
R9180 vp_p.n17906 vp_p.n17905 13.653
R9181 vp_p.n16479 vp_p.n16478 13.653
R9182 vp_p.n15051 vp_p.n15050 13.653
R9183 vp_p.n13721 vp_p.n13720 13.653
R9184 vp_p.n13719 vp_p.n13718 13.653
R9185 vp_p.n7509 vp_p.n7508 13.653
R9186 vp_p.n6087 vp_p.n6086 13.653
R9187 vp_p.n4664 vp_p.n4663 13.653
R9188 vp_p.n3240 vp_p.n3239 13.653
R9189 vp_p.n1815 vp_p.n1814 13.653
R9190 vp_p.n331 vp_p.n330 13.653
R9191 vp_p.n9070 vp_p.n9069 13.653
R9192 vp_p.n10572 vp_p.n10571 13.653
R9193 vp_p.n12010 vp_p.n12009 13.653
R9194 vp_p.n26214 vp_p.n26213 13.653
R9195 vp_p.n24788 vp_p.n24787 13.653
R9196 vp_p.n23366 vp_p.n23365 13.653
R9197 vp_p.n21943 vp_p.n21942 13.653
R9198 vp_p.n20519 vp_p.n20518 13.653
R9199 vp_p.n19094 vp_p.n19093 13.653
R9200 vp_p.n17668 vp_p.n17667 13.653
R9201 vp_p.n16241 vp_p.n16240 13.653
R9202 vp_p.n14813 vp_p.n14812 13.653
R9203 vp_p.n13714 vp_p.n13713 13.653
R9204 vp_p.n7761 vp_p.n7760 13.653
R9205 vp_p.n6339 vp_p.n6338 13.653
R9206 vp_p.n4916 vp_p.n4915 13.653
R9207 vp_p.n3492 vp_p.n3491 13.653
R9208 vp_p.n2067 vp_p.n2066 13.653
R9209 vp_p.n641 vp_p.n640 13.653
R9210 vp_p.n9387 vp_p.n9386 13.653
R9211 vp_p.n10824 vp_p.n10823 13.653
R9212 vp_p.n12262 vp_p.n12261 13.653
R9213 vp_p.n26465 vp_p.n26464 13.653
R9214 vp_p.n25040 vp_p.n25039 13.653
R9215 vp_p.n23618 vp_p.n23617 13.653
R9216 vp_p.n22195 vp_p.n22194 13.653
R9217 vp_p.n20771 vp_p.n20770 13.653
R9218 vp_p.n19346 vp_p.n19345 13.653
R9219 vp_p.n17920 vp_p.n17919 13.653
R9220 vp_p.n16493 vp_p.n16492 13.653
R9221 vp_p.n15065 vp_p.n15064 13.653
R9222 vp_p.n13711 vp_p.n13710 13.653
R9223 vp_p.n13709 vp_p.n13708 13.653
R9224 vp_p.n7504 vp_p.n7503 13.653
R9225 vp_p.n6082 vp_p.n6081 13.653
R9226 vp_p.n4659 vp_p.n4658 13.653
R9227 vp_p.n3235 vp_p.n3234 13.653
R9228 vp_p.n1810 vp_p.n1809 13.653
R9229 vp_p.n326 vp_p.n325 13.653
R9230 vp_p.n9065 vp_p.n9064 13.653
R9231 vp_p.n10567 vp_p.n10566 13.653
R9232 vp_p.n12005 vp_p.n12004 13.653
R9233 vp_p.n26209 vp_p.n26208 13.653
R9234 vp_p.n24783 vp_p.n24782 13.653
R9235 vp_p.n23361 vp_p.n23360 13.653
R9236 vp_p.n21938 vp_p.n21937 13.653
R9237 vp_p.n20514 vp_p.n20513 13.653
R9238 vp_p.n19089 vp_p.n19088 13.653
R9239 vp_p.n17663 vp_p.n17662 13.653
R9240 vp_p.n16236 vp_p.n16235 13.653
R9241 vp_p.n14808 vp_p.n14807 13.653
R9242 vp_p.n13704 vp_p.n13703 13.653
R9243 vp_p.n7775 vp_p.n7774 13.653
R9244 vp_p.n6353 vp_p.n6352 13.653
R9245 vp_p.n4930 vp_p.n4929 13.653
R9246 vp_p.n3506 vp_p.n3505 13.653
R9247 vp_p.n2081 vp_p.n2080 13.653
R9248 vp_p.n655 vp_p.n654 13.653
R9249 vp_p.n9401 vp_p.n9400 13.653
R9250 vp_p.n10838 vp_p.n10837 13.653
R9251 vp_p.n12276 vp_p.n12275 13.653
R9252 vp_p.n26479 vp_p.n26478 13.653
R9253 vp_p.n25054 vp_p.n25053 13.653
R9254 vp_p.n23632 vp_p.n23631 13.653
R9255 vp_p.n22209 vp_p.n22208 13.653
R9256 vp_p.n20785 vp_p.n20784 13.653
R9257 vp_p.n19360 vp_p.n19359 13.653
R9258 vp_p.n17934 vp_p.n17933 13.653
R9259 vp_p.n16507 vp_p.n16506 13.653
R9260 vp_p.n15079 vp_p.n15078 13.653
R9261 vp_p.n13701 vp_p.n13700 13.653
R9262 vp_p.n13699 vp_p.n13698 13.653
R9263 vp_p.n7499 vp_p.n7498 13.653
R9264 vp_p.n6077 vp_p.n6076 13.653
R9265 vp_p.n4654 vp_p.n4653 13.653
R9266 vp_p.n3230 vp_p.n3229 13.653
R9267 vp_p.n1805 vp_p.n1804 13.653
R9268 vp_p.n321 vp_p.n320 13.653
R9269 vp_p.n9060 vp_p.n9059 13.653
R9270 vp_p.n10562 vp_p.n10561 13.653
R9271 vp_p.n12000 vp_p.n11999 13.653
R9272 vp_p.n26204 vp_p.n26203 13.653
R9273 vp_p.n24778 vp_p.n24777 13.653
R9274 vp_p.n23356 vp_p.n23355 13.653
R9275 vp_p.n21933 vp_p.n21932 13.653
R9276 vp_p.n20509 vp_p.n20508 13.653
R9277 vp_p.n19084 vp_p.n19083 13.653
R9278 vp_p.n17658 vp_p.n17657 13.653
R9279 vp_p.n16231 vp_p.n16230 13.653
R9280 vp_p.n14803 vp_p.n14802 13.653
R9281 vp_p.n13694 vp_p.n13693 13.653
R9282 vp_p.n7789 vp_p.n7788 13.653
R9283 vp_p.n6367 vp_p.n6366 13.653
R9284 vp_p.n4944 vp_p.n4943 13.653
R9285 vp_p.n3520 vp_p.n3519 13.653
R9286 vp_p.n2095 vp_p.n2094 13.653
R9287 vp_p.n669 vp_p.n668 13.653
R9288 vp_p.n9415 vp_p.n9414 13.653
R9289 vp_p.n10852 vp_p.n10851 13.653
R9290 vp_p.n12290 vp_p.n12289 13.653
R9291 vp_p.n26493 vp_p.n26492 13.653
R9292 vp_p.n25068 vp_p.n25067 13.653
R9293 vp_p.n23646 vp_p.n23645 13.653
R9294 vp_p.n22223 vp_p.n22222 13.653
R9295 vp_p.n20799 vp_p.n20798 13.653
R9296 vp_p.n19374 vp_p.n19373 13.653
R9297 vp_p.n17948 vp_p.n17947 13.653
R9298 vp_p.n16521 vp_p.n16520 13.653
R9299 vp_p.n15093 vp_p.n15092 13.653
R9300 vp_p.n13691 vp_p.n13690 13.653
R9301 vp_p.n13689 vp_p.n13688 13.653
R9302 vp_p.n7494 vp_p.n7493 13.653
R9303 vp_p.n6072 vp_p.n6071 13.653
R9304 vp_p.n4649 vp_p.n4648 13.653
R9305 vp_p.n3225 vp_p.n3224 13.653
R9306 vp_p.n1800 vp_p.n1799 13.653
R9307 vp_p.n316 vp_p.n315 13.653
R9308 vp_p.n9055 vp_p.n9054 13.653
R9309 vp_p.n10557 vp_p.n10556 13.653
R9310 vp_p.n11995 vp_p.n11994 13.653
R9311 vp_p.n26199 vp_p.n26198 13.653
R9312 vp_p.n24773 vp_p.n24772 13.653
R9313 vp_p.n23351 vp_p.n23350 13.653
R9314 vp_p.n21928 vp_p.n21927 13.653
R9315 vp_p.n20504 vp_p.n20503 13.653
R9316 vp_p.n19079 vp_p.n19078 13.653
R9317 vp_p.n17653 vp_p.n17652 13.653
R9318 vp_p.n16226 vp_p.n16225 13.653
R9319 vp_p.n14798 vp_p.n14797 13.653
R9320 vp_p.n13684 vp_p.n13683 13.653
R9321 vp_p.n7803 vp_p.n7802 13.653
R9322 vp_p.n6381 vp_p.n6380 13.653
R9323 vp_p.n4958 vp_p.n4957 13.653
R9324 vp_p.n3534 vp_p.n3533 13.653
R9325 vp_p.n2109 vp_p.n2108 13.653
R9326 vp_p.n683 vp_p.n682 13.653
R9327 vp_p.n9429 vp_p.n9428 13.653
R9328 vp_p.n10866 vp_p.n10865 13.653
R9329 vp_p.n12304 vp_p.n12303 13.653
R9330 vp_p.n26507 vp_p.n26506 13.653
R9331 vp_p.n25082 vp_p.n25081 13.653
R9332 vp_p.n23660 vp_p.n23659 13.653
R9333 vp_p.n22237 vp_p.n22236 13.653
R9334 vp_p.n20813 vp_p.n20812 13.653
R9335 vp_p.n19388 vp_p.n19387 13.653
R9336 vp_p.n17962 vp_p.n17961 13.653
R9337 vp_p.n16535 vp_p.n16534 13.653
R9338 vp_p.n15107 vp_p.n15106 13.653
R9339 vp_p.n13681 vp_p.n13680 13.653
R9340 vp_p.n13679 vp_p.n13678 13.653
R9341 vp_p.n7489 vp_p.n7488 13.653
R9342 vp_p.n6067 vp_p.n6066 13.653
R9343 vp_p.n4644 vp_p.n4643 13.653
R9344 vp_p.n3220 vp_p.n3219 13.653
R9345 vp_p.n1795 vp_p.n1794 13.653
R9346 vp_p.n311 vp_p.n310 13.653
R9347 vp_p.n9050 vp_p.n9049 13.653
R9348 vp_p.n10552 vp_p.n10551 13.653
R9349 vp_p.n11990 vp_p.n11989 13.653
R9350 vp_p.n26194 vp_p.n26193 13.653
R9351 vp_p.n24768 vp_p.n24767 13.653
R9352 vp_p.n23346 vp_p.n23345 13.653
R9353 vp_p.n21923 vp_p.n21922 13.653
R9354 vp_p.n20499 vp_p.n20498 13.653
R9355 vp_p.n19074 vp_p.n19073 13.653
R9356 vp_p.n17648 vp_p.n17647 13.653
R9357 vp_p.n16221 vp_p.n16220 13.653
R9358 vp_p.n14793 vp_p.n14792 13.653
R9359 vp_p.n13674 vp_p.n13673 13.653
R9360 vp_p.n7817 vp_p.n7816 13.653
R9361 vp_p.n6395 vp_p.n6394 13.653
R9362 vp_p.n4972 vp_p.n4971 13.653
R9363 vp_p.n3548 vp_p.n3547 13.653
R9364 vp_p.n2123 vp_p.n2122 13.653
R9365 vp_p.n697 vp_p.n696 13.653
R9366 vp_p.n9443 vp_p.n9442 13.653
R9367 vp_p.n10880 vp_p.n10879 13.653
R9368 vp_p.n12318 vp_p.n12317 13.653
R9369 vp_p.n26521 vp_p.n26520 13.653
R9370 vp_p.n25096 vp_p.n25095 13.653
R9371 vp_p.n23674 vp_p.n23673 13.653
R9372 vp_p.n22251 vp_p.n22250 13.653
R9373 vp_p.n20827 vp_p.n20826 13.653
R9374 vp_p.n19402 vp_p.n19401 13.653
R9375 vp_p.n17976 vp_p.n17975 13.653
R9376 vp_p.n16549 vp_p.n16548 13.653
R9377 vp_p.n15121 vp_p.n15120 13.653
R9378 vp_p.n13671 vp_p.n13670 13.653
R9379 vp_p.n13669 vp_p.n13668 13.653
R9380 vp_p.n7484 vp_p.n7483 13.653
R9381 vp_p.n6062 vp_p.n6061 13.653
R9382 vp_p.n4639 vp_p.n4638 13.653
R9383 vp_p.n3215 vp_p.n3214 13.653
R9384 vp_p.n1790 vp_p.n1789 13.653
R9385 vp_p.n306 vp_p.n305 13.653
R9386 vp_p.n9045 vp_p.n9044 13.653
R9387 vp_p.n10547 vp_p.n10546 13.653
R9388 vp_p.n11985 vp_p.n11984 13.653
R9389 vp_p.n26189 vp_p.n26188 13.653
R9390 vp_p.n24763 vp_p.n24762 13.653
R9391 vp_p.n23341 vp_p.n23340 13.653
R9392 vp_p.n21918 vp_p.n21917 13.653
R9393 vp_p.n20494 vp_p.n20493 13.653
R9394 vp_p.n19069 vp_p.n19068 13.653
R9395 vp_p.n17643 vp_p.n17642 13.653
R9396 vp_p.n16216 vp_p.n16215 13.653
R9397 vp_p.n14788 vp_p.n14787 13.653
R9398 vp_p.n13664 vp_p.n13663 13.653
R9399 vp_p.n7831 vp_p.n7830 13.653
R9400 vp_p.n6409 vp_p.n6408 13.653
R9401 vp_p.n4986 vp_p.n4985 13.653
R9402 vp_p.n3562 vp_p.n3561 13.653
R9403 vp_p.n2137 vp_p.n2136 13.653
R9404 vp_p.n711 vp_p.n710 13.653
R9405 vp_p.n9457 vp_p.n9456 13.653
R9406 vp_p.n10894 vp_p.n10893 13.653
R9407 vp_p.n12332 vp_p.n12331 13.653
R9408 vp_p.n26535 vp_p.n26534 13.653
R9409 vp_p.n25110 vp_p.n25109 13.653
R9410 vp_p.n23688 vp_p.n23687 13.653
R9411 vp_p.n22265 vp_p.n22264 13.653
R9412 vp_p.n20841 vp_p.n20840 13.653
R9413 vp_p.n19416 vp_p.n19415 13.653
R9414 vp_p.n17990 vp_p.n17989 13.653
R9415 vp_p.n16563 vp_p.n16562 13.653
R9416 vp_p.n15135 vp_p.n15134 13.653
R9417 vp_p.n13661 vp_p.n13660 13.653
R9418 vp_p.n13659 vp_p.n13658 13.653
R9419 vp_p.n7479 vp_p.n7478 13.653
R9420 vp_p.n6057 vp_p.n6056 13.653
R9421 vp_p.n4634 vp_p.n4633 13.653
R9422 vp_p.n3210 vp_p.n3209 13.653
R9423 vp_p.n1785 vp_p.n1784 13.653
R9424 vp_p.n301 vp_p.n300 13.653
R9425 vp_p.n9040 vp_p.n9039 13.653
R9426 vp_p.n10542 vp_p.n10541 13.653
R9427 vp_p.n11980 vp_p.n11979 13.653
R9428 vp_p.n26184 vp_p.n26183 13.653
R9429 vp_p.n24758 vp_p.n24757 13.653
R9430 vp_p.n23336 vp_p.n23335 13.653
R9431 vp_p.n21913 vp_p.n21912 13.653
R9432 vp_p.n20489 vp_p.n20488 13.653
R9433 vp_p.n19064 vp_p.n19063 13.653
R9434 vp_p.n17638 vp_p.n17637 13.653
R9435 vp_p.n16211 vp_p.n16210 13.653
R9436 vp_p.n14783 vp_p.n14782 13.653
R9437 vp_p.n13654 vp_p.n13653 13.653
R9438 vp_p.n7845 vp_p.n7844 13.653
R9439 vp_p.n6423 vp_p.n6422 13.653
R9440 vp_p.n5000 vp_p.n4999 13.653
R9441 vp_p.n3576 vp_p.n3575 13.653
R9442 vp_p.n2151 vp_p.n2150 13.653
R9443 vp_p.n725 vp_p.n724 13.653
R9444 vp_p.n9471 vp_p.n9470 13.653
R9445 vp_p.n10908 vp_p.n10907 13.653
R9446 vp_p.n12346 vp_p.n12345 13.653
R9447 vp_p.n26549 vp_p.n26548 13.653
R9448 vp_p.n25124 vp_p.n25123 13.653
R9449 vp_p.n23702 vp_p.n23701 13.653
R9450 vp_p.n22279 vp_p.n22278 13.653
R9451 vp_p.n20855 vp_p.n20854 13.653
R9452 vp_p.n19430 vp_p.n19429 13.653
R9453 vp_p.n18004 vp_p.n18003 13.653
R9454 vp_p.n16577 vp_p.n16576 13.653
R9455 vp_p.n15149 vp_p.n15148 13.653
R9456 vp_p.n13651 vp_p.n13650 13.653
R9457 vp_p.n13649 vp_p.n13648 13.653
R9458 vp_p.n7474 vp_p.n7473 13.653
R9459 vp_p.n6052 vp_p.n6051 13.653
R9460 vp_p.n4629 vp_p.n4628 13.653
R9461 vp_p.n3205 vp_p.n3204 13.653
R9462 vp_p.n1780 vp_p.n1779 13.653
R9463 vp_p.n296 vp_p.n295 13.653
R9464 vp_p.n9035 vp_p.n9034 13.653
R9465 vp_p.n10537 vp_p.n10536 13.653
R9466 vp_p.n11975 vp_p.n11974 13.653
R9467 vp_p.n26179 vp_p.n26178 13.653
R9468 vp_p.n24753 vp_p.n24752 13.653
R9469 vp_p.n23331 vp_p.n23330 13.653
R9470 vp_p.n21908 vp_p.n21907 13.653
R9471 vp_p.n20484 vp_p.n20483 13.653
R9472 vp_p.n19059 vp_p.n19058 13.653
R9473 vp_p.n17633 vp_p.n17632 13.653
R9474 vp_p.n16206 vp_p.n16205 13.653
R9475 vp_p.n14778 vp_p.n14777 13.653
R9476 vp_p.n13644 vp_p.n13643 13.653
R9477 vp_p.n7859 vp_p.n7858 13.653
R9478 vp_p.n6437 vp_p.n6436 13.653
R9479 vp_p.n5014 vp_p.n5013 13.653
R9480 vp_p.n3590 vp_p.n3589 13.653
R9481 vp_p.n2165 vp_p.n2164 13.653
R9482 vp_p.n739 vp_p.n738 13.653
R9483 vp_p.n9485 vp_p.n9484 13.653
R9484 vp_p.n10922 vp_p.n10921 13.653
R9485 vp_p.n12360 vp_p.n12359 13.653
R9486 vp_p.n26563 vp_p.n26562 13.653
R9487 vp_p.n25138 vp_p.n25137 13.653
R9488 vp_p.n23716 vp_p.n23715 13.653
R9489 vp_p.n22293 vp_p.n22292 13.653
R9490 vp_p.n20869 vp_p.n20868 13.653
R9491 vp_p.n19444 vp_p.n19443 13.653
R9492 vp_p.n18018 vp_p.n18017 13.653
R9493 vp_p.n16591 vp_p.n16590 13.653
R9494 vp_p.n15163 vp_p.n15162 13.653
R9495 vp_p.n13641 vp_p.n13640 13.653
R9496 vp_p.n13639 vp_p.n13638 13.653
R9497 vp_p.n7469 vp_p.n7468 13.653
R9498 vp_p.n6047 vp_p.n6046 13.653
R9499 vp_p.n4624 vp_p.n4623 13.653
R9500 vp_p.n3200 vp_p.n3199 13.653
R9501 vp_p.n1775 vp_p.n1774 13.653
R9502 vp_p.n291 vp_p.n290 13.653
R9503 vp_p.n9030 vp_p.n9029 13.653
R9504 vp_p.n10532 vp_p.n10531 13.653
R9505 vp_p.n11970 vp_p.n11969 13.653
R9506 vp_p.n26174 vp_p.n26173 13.653
R9507 vp_p.n24748 vp_p.n24747 13.653
R9508 vp_p.n23326 vp_p.n23325 13.653
R9509 vp_p.n21903 vp_p.n21902 13.653
R9510 vp_p.n20479 vp_p.n20478 13.653
R9511 vp_p.n19054 vp_p.n19053 13.653
R9512 vp_p.n17628 vp_p.n17627 13.653
R9513 vp_p.n16201 vp_p.n16200 13.653
R9514 vp_p.n14773 vp_p.n14772 13.653
R9515 vp_p.n13634 vp_p.n13633 13.653
R9516 vp_p.n7873 vp_p.n7872 13.653
R9517 vp_p.n6451 vp_p.n6450 13.653
R9518 vp_p.n5028 vp_p.n5027 13.653
R9519 vp_p.n3604 vp_p.n3603 13.653
R9520 vp_p.n2179 vp_p.n2178 13.653
R9521 vp_p.n753 vp_p.n752 13.653
R9522 vp_p.n9499 vp_p.n9498 13.653
R9523 vp_p.n10936 vp_p.n10935 13.653
R9524 vp_p.n12374 vp_p.n12373 13.653
R9525 vp_p.n26577 vp_p.n26576 13.653
R9526 vp_p.n25152 vp_p.n25151 13.653
R9527 vp_p.n23730 vp_p.n23729 13.653
R9528 vp_p.n22307 vp_p.n22306 13.653
R9529 vp_p.n20883 vp_p.n20882 13.653
R9530 vp_p.n19458 vp_p.n19457 13.653
R9531 vp_p.n18032 vp_p.n18031 13.653
R9532 vp_p.n16605 vp_p.n16604 13.653
R9533 vp_p.n15177 vp_p.n15176 13.653
R9534 vp_p.n13631 vp_p.n13630 13.653
R9535 vp_p.n13629 vp_p.n13628 13.653
R9536 vp_p.n7464 vp_p.n7463 13.653
R9537 vp_p.n6042 vp_p.n6041 13.653
R9538 vp_p.n4619 vp_p.n4618 13.653
R9539 vp_p.n3195 vp_p.n3194 13.653
R9540 vp_p.n1770 vp_p.n1769 13.653
R9541 vp_p.n286 vp_p.n285 13.653
R9542 vp_p.n9025 vp_p.n9024 13.653
R9543 vp_p.n10527 vp_p.n10526 13.653
R9544 vp_p.n11965 vp_p.n11964 13.653
R9545 vp_p.n26169 vp_p.n26168 13.653
R9546 vp_p.n24743 vp_p.n24742 13.653
R9547 vp_p.n23321 vp_p.n23320 13.653
R9548 vp_p.n21898 vp_p.n21897 13.653
R9549 vp_p.n20474 vp_p.n20473 13.653
R9550 vp_p.n19049 vp_p.n19048 13.653
R9551 vp_p.n17623 vp_p.n17622 13.653
R9552 vp_p.n16196 vp_p.n16195 13.653
R9553 vp_p.n14768 vp_p.n14767 13.653
R9554 vp_p.n13624 vp_p.n13623 13.653
R9555 vp_p.n7887 vp_p.n7886 13.653
R9556 vp_p.n6465 vp_p.n6464 13.653
R9557 vp_p.n5042 vp_p.n5041 13.653
R9558 vp_p.n3618 vp_p.n3617 13.653
R9559 vp_p.n2193 vp_p.n2192 13.653
R9560 vp_p.n767 vp_p.n766 13.653
R9561 vp_p.n9513 vp_p.n9512 13.653
R9562 vp_p.n10950 vp_p.n10949 13.653
R9563 vp_p.n12388 vp_p.n12387 13.653
R9564 vp_p.n26591 vp_p.n26590 13.653
R9565 vp_p.n25166 vp_p.n25165 13.653
R9566 vp_p.n23744 vp_p.n23743 13.653
R9567 vp_p.n22321 vp_p.n22320 13.653
R9568 vp_p.n20897 vp_p.n20896 13.653
R9569 vp_p.n19472 vp_p.n19471 13.653
R9570 vp_p.n18046 vp_p.n18045 13.653
R9571 vp_p.n16619 vp_p.n16618 13.653
R9572 vp_p.n15191 vp_p.n15190 13.653
R9573 vp_p.n13621 vp_p.n13620 13.653
R9574 vp_p.n13619 vp_p.n13618 13.653
R9575 vp_p.n7459 vp_p.n7458 13.653
R9576 vp_p.n6037 vp_p.n6036 13.653
R9577 vp_p.n4614 vp_p.n4613 13.653
R9578 vp_p.n3190 vp_p.n3189 13.653
R9579 vp_p.n1765 vp_p.n1764 13.653
R9580 vp_p.n281 vp_p.n280 13.653
R9581 vp_p.n9020 vp_p.n9019 13.653
R9582 vp_p.n10522 vp_p.n10521 13.653
R9583 vp_p.n11960 vp_p.n11959 13.653
R9584 vp_p.n26164 vp_p.n26163 13.653
R9585 vp_p.n24738 vp_p.n24737 13.653
R9586 vp_p.n23316 vp_p.n23315 13.653
R9587 vp_p.n21893 vp_p.n21892 13.653
R9588 vp_p.n20469 vp_p.n20468 13.653
R9589 vp_p.n19044 vp_p.n19043 13.653
R9590 vp_p.n17618 vp_p.n17617 13.653
R9591 vp_p.n16191 vp_p.n16190 13.653
R9592 vp_p.n14763 vp_p.n14762 13.653
R9593 vp_p.n13614 vp_p.n13613 13.653
R9594 vp_p.n7901 vp_p.n7900 13.653
R9595 vp_p.n6479 vp_p.n6478 13.653
R9596 vp_p.n5056 vp_p.n5055 13.653
R9597 vp_p.n3632 vp_p.n3631 13.653
R9598 vp_p.n2207 vp_p.n2206 13.653
R9599 vp_p.n781 vp_p.n780 13.653
R9600 vp_p.n9527 vp_p.n9526 13.653
R9601 vp_p.n10964 vp_p.n10963 13.653
R9602 vp_p.n12402 vp_p.n12401 13.653
R9603 vp_p.n26605 vp_p.n26604 13.653
R9604 vp_p.n25180 vp_p.n25179 13.653
R9605 vp_p.n23758 vp_p.n23757 13.653
R9606 vp_p.n22335 vp_p.n22334 13.653
R9607 vp_p.n20911 vp_p.n20910 13.653
R9608 vp_p.n19486 vp_p.n19485 13.653
R9609 vp_p.n18060 vp_p.n18059 13.653
R9610 vp_p.n16633 vp_p.n16632 13.653
R9611 vp_p.n15205 vp_p.n15204 13.653
R9612 vp_p.n13611 vp_p.n13610 13.653
R9613 vp_p.n13609 vp_p.n13608 13.653
R9614 vp_p.n7454 vp_p.n7453 13.653
R9615 vp_p.n6032 vp_p.n6031 13.653
R9616 vp_p.n4609 vp_p.n4608 13.653
R9617 vp_p.n3185 vp_p.n3184 13.653
R9618 vp_p.n1760 vp_p.n1759 13.653
R9619 vp_p.n276 vp_p.n275 13.653
R9620 vp_p.n9015 vp_p.n9014 13.653
R9621 vp_p.n10517 vp_p.n10516 13.653
R9622 vp_p.n11955 vp_p.n11954 13.653
R9623 vp_p.n26159 vp_p.n26158 13.653
R9624 vp_p.n24733 vp_p.n24732 13.653
R9625 vp_p.n23311 vp_p.n23310 13.653
R9626 vp_p.n21888 vp_p.n21887 13.653
R9627 vp_p.n20464 vp_p.n20463 13.653
R9628 vp_p.n19039 vp_p.n19038 13.653
R9629 vp_p.n17613 vp_p.n17612 13.653
R9630 vp_p.n16186 vp_p.n16185 13.653
R9631 vp_p.n14758 vp_p.n14757 13.653
R9632 vp_p.n13604 vp_p.n13603 13.653
R9633 vp_p.n7915 vp_p.n7914 13.653
R9634 vp_p.n6493 vp_p.n6492 13.653
R9635 vp_p.n5070 vp_p.n5069 13.653
R9636 vp_p.n3646 vp_p.n3645 13.653
R9637 vp_p.n2221 vp_p.n2220 13.653
R9638 vp_p.n795 vp_p.n794 13.653
R9639 vp_p.n9541 vp_p.n9540 13.653
R9640 vp_p.n10978 vp_p.n10977 13.653
R9641 vp_p.n12416 vp_p.n12415 13.653
R9642 vp_p.n26619 vp_p.n26618 13.653
R9643 vp_p.n25194 vp_p.n25193 13.653
R9644 vp_p.n23772 vp_p.n23771 13.653
R9645 vp_p.n22349 vp_p.n22348 13.653
R9646 vp_p.n20925 vp_p.n20924 13.653
R9647 vp_p.n19500 vp_p.n19499 13.653
R9648 vp_p.n18074 vp_p.n18073 13.653
R9649 vp_p.n16647 vp_p.n16646 13.653
R9650 vp_p.n15219 vp_p.n15218 13.653
R9651 vp_p.n13601 vp_p.n13600 13.653
R9652 vp_p.n13599 vp_p.n13598 13.653
R9653 vp_p.n7449 vp_p.n7448 13.653
R9654 vp_p.n6027 vp_p.n6026 13.653
R9655 vp_p.n4604 vp_p.n4603 13.653
R9656 vp_p.n3180 vp_p.n3179 13.653
R9657 vp_p.n1755 vp_p.n1754 13.653
R9658 vp_p.n271 vp_p.n270 13.653
R9659 vp_p.n9010 vp_p.n9009 13.653
R9660 vp_p.n10512 vp_p.n10511 13.653
R9661 vp_p.n11950 vp_p.n11949 13.653
R9662 vp_p.n26154 vp_p.n26153 13.653
R9663 vp_p.n24728 vp_p.n24727 13.653
R9664 vp_p.n23306 vp_p.n23305 13.653
R9665 vp_p.n21883 vp_p.n21882 13.653
R9666 vp_p.n20459 vp_p.n20458 13.653
R9667 vp_p.n19034 vp_p.n19033 13.653
R9668 vp_p.n17608 vp_p.n17607 13.653
R9669 vp_p.n16181 vp_p.n16180 13.653
R9670 vp_p.n14753 vp_p.n14752 13.653
R9671 vp_p.n13594 vp_p.n13593 13.653
R9672 vp_p.n7929 vp_p.n7928 13.653
R9673 vp_p.n6507 vp_p.n6506 13.653
R9674 vp_p.n5084 vp_p.n5083 13.653
R9675 vp_p.n3660 vp_p.n3659 13.653
R9676 vp_p.n2235 vp_p.n2234 13.653
R9677 vp_p.n809 vp_p.n808 13.653
R9678 vp_p.n9555 vp_p.n9554 13.653
R9679 vp_p.n10992 vp_p.n10991 13.653
R9680 vp_p.n12430 vp_p.n12429 13.653
R9681 vp_p.n26633 vp_p.n26632 13.653
R9682 vp_p.n25208 vp_p.n25207 13.653
R9683 vp_p.n23786 vp_p.n23785 13.653
R9684 vp_p.n22363 vp_p.n22362 13.653
R9685 vp_p.n20939 vp_p.n20938 13.653
R9686 vp_p.n19514 vp_p.n19513 13.653
R9687 vp_p.n18088 vp_p.n18087 13.653
R9688 vp_p.n16661 vp_p.n16660 13.653
R9689 vp_p.n15233 vp_p.n15232 13.653
R9690 vp_p.n13591 vp_p.n13590 13.653
R9691 vp_p.n13589 vp_p.n13588 13.653
R9692 vp_p.n7444 vp_p.n7443 13.653
R9693 vp_p.n6022 vp_p.n6021 13.653
R9694 vp_p.n4599 vp_p.n4598 13.653
R9695 vp_p.n3175 vp_p.n3174 13.653
R9696 vp_p.n1750 vp_p.n1749 13.653
R9697 vp_p.n266 vp_p.n265 13.653
R9698 vp_p.n9005 vp_p.n9004 13.653
R9699 vp_p.n10507 vp_p.n10506 13.653
R9700 vp_p.n11945 vp_p.n11944 13.653
R9701 vp_p.n26149 vp_p.n26148 13.653
R9702 vp_p.n24723 vp_p.n24722 13.653
R9703 vp_p.n23301 vp_p.n23300 13.653
R9704 vp_p.n21878 vp_p.n21877 13.653
R9705 vp_p.n20454 vp_p.n20453 13.653
R9706 vp_p.n19029 vp_p.n19028 13.653
R9707 vp_p.n17603 vp_p.n17602 13.653
R9708 vp_p.n16176 vp_p.n16175 13.653
R9709 vp_p.n14748 vp_p.n14747 13.653
R9710 vp_p.n13584 vp_p.n13583 13.653
R9711 vp_p.n7943 vp_p.n7942 13.653
R9712 vp_p.n6521 vp_p.n6520 13.653
R9713 vp_p.n5098 vp_p.n5097 13.653
R9714 vp_p.n3674 vp_p.n3673 13.653
R9715 vp_p.n2249 vp_p.n2248 13.653
R9716 vp_p.n823 vp_p.n822 13.653
R9717 vp_p.n9569 vp_p.n9568 13.653
R9718 vp_p.n11006 vp_p.n11005 13.653
R9719 vp_p.n12444 vp_p.n12443 13.653
R9720 vp_p.n26647 vp_p.n26646 13.653
R9721 vp_p.n25222 vp_p.n25221 13.653
R9722 vp_p.n23800 vp_p.n23799 13.653
R9723 vp_p.n22377 vp_p.n22376 13.653
R9724 vp_p.n20953 vp_p.n20952 13.653
R9725 vp_p.n19528 vp_p.n19527 13.653
R9726 vp_p.n18102 vp_p.n18101 13.653
R9727 vp_p.n16675 vp_p.n16674 13.653
R9728 vp_p.n15247 vp_p.n15246 13.653
R9729 vp_p.n13581 vp_p.n13580 13.653
R9730 vp_p.n13579 vp_p.n13578 13.653
R9731 vp_p.n7439 vp_p.n7438 13.653
R9732 vp_p.n6017 vp_p.n6016 13.653
R9733 vp_p.n4594 vp_p.n4593 13.653
R9734 vp_p.n3170 vp_p.n3169 13.653
R9735 vp_p.n1745 vp_p.n1744 13.653
R9736 vp_p.n261 vp_p.n260 13.653
R9737 vp_p.n9000 vp_p.n8999 13.653
R9738 vp_p.n10502 vp_p.n10501 13.653
R9739 vp_p.n11940 vp_p.n11939 13.653
R9740 vp_p.n26144 vp_p.n26143 13.653
R9741 vp_p.n24718 vp_p.n24717 13.653
R9742 vp_p.n23296 vp_p.n23295 13.653
R9743 vp_p.n21873 vp_p.n21872 13.653
R9744 vp_p.n20449 vp_p.n20448 13.653
R9745 vp_p.n19024 vp_p.n19023 13.653
R9746 vp_p.n17598 vp_p.n17597 13.653
R9747 vp_p.n16171 vp_p.n16170 13.653
R9748 vp_p.n14743 vp_p.n14742 13.653
R9749 vp_p.n13574 vp_p.n13573 13.653
R9750 vp_p.n7957 vp_p.n7956 13.653
R9751 vp_p.n6535 vp_p.n6534 13.653
R9752 vp_p.n5112 vp_p.n5111 13.653
R9753 vp_p.n3688 vp_p.n3687 13.653
R9754 vp_p.n2263 vp_p.n2262 13.653
R9755 vp_p.n837 vp_p.n836 13.653
R9756 vp_p.n9583 vp_p.n9582 13.653
R9757 vp_p.n11020 vp_p.n11019 13.653
R9758 vp_p.n12458 vp_p.n12457 13.653
R9759 vp_p.n26661 vp_p.n26660 13.653
R9760 vp_p.n25236 vp_p.n25235 13.653
R9761 vp_p.n23814 vp_p.n23813 13.653
R9762 vp_p.n22391 vp_p.n22390 13.653
R9763 vp_p.n20967 vp_p.n20966 13.653
R9764 vp_p.n19542 vp_p.n19541 13.653
R9765 vp_p.n18116 vp_p.n18115 13.653
R9766 vp_p.n16689 vp_p.n16688 13.653
R9767 vp_p.n15261 vp_p.n15260 13.653
R9768 vp_p.n13571 vp_p.n13570 13.653
R9769 vp_p.n13569 vp_p.n13568 13.653
R9770 vp_p.n7434 vp_p.n7433 13.653
R9771 vp_p.n6012 vp_p.n6011 13.653
R9772 vp_p.n4589 vp_p.n4588 13.653
R9773 vp_p.n3165 vp_p.n3164 13.653
R9774 vp_p.n1740 vp_p.n1739 13.653
R9775 vp_p.n256 vp_p.n255 13.653
R9776 vp_p.n8995 vp_p.n8994 13.653
R9777 vp_p.n10497 vp_p.n10496 13.653
R9778 vp_p.n11935 vp_p.n11934 13.653
R9779 vp_p.n26139 vp_p.n26138 13.653
R9780 vp_p.n24713 vp_p.n24712 13.653
R9781 vp_p.n23291 vp_p.n23290 13.653
R9782 vp_p.n21868 vp_p.n21867 13.653
R9783 vp_p.n20444 vp_p.n20443 13.653
R9784 vp_p.n19019 vp_p.n19018 13.653
R9785 vp_p.n17593 vp_p.n17592 13.653
R9786 vp_p.n16166 vp_p.n16165 13.653
R9787 vp_p.n14738 vp_p.n14737 13.653
R9788 vp_p.n13564 vp_p.n13563 13.653
R9789 vp_p.n7971 vp_p.n7970 13.653
R9790 vp_p.n6549 vp_p.n6548 13.653
R9791 vp_p.n5126 vp_p.n5125 13.653
R9792 vp_p.n3702 vp_p.n3701 13.653
R9793 vp_p.n2277 vp_p.n2276 13.653
R9794 vp_p.n851 vp_p.n850 13.653
R9795 vp_p.n9597 vp_p.n9596 13.653
R9796 vp_p.n11034 vp_p.n11033 13.653
R9797 vp_p.n12472 vp_p.n12471 13.653
R9798 vp_p.n26675 vp_p.n26674 13.653
R9799 vp_p.n25250 vp_p.n25249 13.653
R9800 vp_p.n23828 vp_p.n23827 13.653
R9801 vp_p.n22405 vp_p.n22404 13.653
R9802 vp_p.n20981 vp_p.n20980 13.653
R9803 vp_p.n19556 vp_p.n19555 13.653
R9804 vp_p.n18130 vp_p.n18129 13.653
R9805 vp_p.n16703 vp_p.n16702 13.653
R9806 vp_p.n15275 vp_p.n15274 13.653
R9807 vp_p.n13561 vp_p.n13560 13.653
R9808 vp_p.n13559 vp_p.n13558 13.653
R9809 vp_p.n7429 vp_p.n7428 13.653
R9810 vp_p.n6007 vp_p.n6006 13.653
R9811 vp_p.n4584 vp_p.n4583 13.653
R9812 vp_p.n3160 vp_p.n3159 13.653
R9813 vp_p.n1735 vp_p.n1734 13.653
R9814 vp_p.n251 vp_p.n250 13.653
R9815 vp_p.n8990 vp_p.n8989 13.653
R9816 vp_p.n10492 vp_p.n10491 13.653
R9817 vp_p.n11930 vp_p.n11929 13.653
R9818 vp_p.n26134 vp_p.n26133 13.653
R9819 vp_p.n24708 vp_p.n24707 13.653
R9820 vp_p.n23286 vp_p.n23285 13.653
R9821 vp_p.n21863 vp_p.n21862 13.653
R9822 vp_p.n20439 vp_p.n20438 13.653
R9823 vp_p.n19014 vp_p.n19013 13.653
R9824 vp_p.n17588 vp_p.n17587 13.653
R9825 vp_p.n16161 vp_p.n16160 13.653
R9826 vp_p.n14733 vp_p.n14732 13.653
R9827 vp_p.n13554 vp_p.n13553 13.653
R9828 vp_p.n7985 vp_p.n7984 13.653
R9829 vp_p.n6563 vp_p.n6562 13.653
R9830 vp_p.n5140 vp_p.n5139 13.653
R9831 vp_p.n3716 vp_p.n3715 13.653
R9832 vp_p.n2291 vp_p.n2290 13.653
R9833 vp_p.n865 vp_p.n864 13.653
R9834 vp_p.n9611 vp_p.n9610 13.653
R9835 vp_p.n11048 vp_p.n11047 13.653
R9836 vp_p.n12486 vp_p.n12485 13.653
R9837 vp_p.n26689 vp_p.n26688 13.653
R9838 vp_p.n25264 vp_p.n25263 13.653
R9839 vp_p.n23842 vp_p.n23841 13.653
R9840 vp_p.n22419 vp_p.n22418 13.653
R9841 vp_p.n20995 vp_p.n20994 13.653
R9842 vp_p.n19570 vp_p.n19569 13.653
R9843 vp_p.n18144 vp_p.n18143 13.653
R9844 vp_p.n16717 vp_p.n16716 13.653
R9845 vp_p.n15289 vp_p.n15288 13.653
R9846 vp_p.n13551 vp_p.n13550 13.653
R9847 vp_p.n13549 vp_p.n13548 13.653
R9848 vp_p.n7424 vp_p.n7423 13.653
R9849 vp_p.n6002 vp_p.n6001 13.653
R9850 vp_p.n4579 vp_p.n4578 13.653
R9851 vp_p.n3155 vp_p.n3154 13.653
R9852 vp_p.n1730 vp_p.n1729 13.653
R9853 vp_p.n246 vp_p.n245 13.653
R9854 vp_p.n8985 vp_p.n8984 13.653
R9855 vp_p.n10487 vp_p.n10486 13.653
R9856 vp_p.n11925 vp_p.n11924 13.653
R9857 vp_p.n26129 vp_p.n26128 13.653
R9858 vp_p.n24703 vp_p.n24702 13.653
R9859 vp_p.n23281 vp_p.n23280 13.653
R9860 vp_p.n21858 vp_p.n21857 13.653
R9861 vp_p.n20434 vp_p.n20433 13.653
R9862 vp_p.n19009 vp_p.n19008 13.653
R9863 vp_p.n17583 vp_p.n17582 13.653
R9864 vp_p.n16156 vp_p.n16155 13.653
R9865 vp_p.n14728 vp_p.n14727 13.653
R9866 vp_p.n13544 vp_p.n13543 13.653
R9867 vp_p.n7999 vp_p.n7998 13.653
R9868 vp_p.n6577 vp_p.n6576 13.653
R9869 vp_p.n5154 vp_p.n5153 13.653
R9870 vp_p.n3730 vp_p.n3729 13.653
R9871 vp_p.n2305 vp_p.n2304 13.653
R9872 vp_p.n879 vp_p.n878 13.653
R9873 vp_p.n9625 vp_p.n9624 13.653
R9874 vp_p.n11062 vp_p.n11061 13.653
R9875 vp_p.n12500 vp_p.n12499 13.653
R9876 vp_p.n26703 vp_p.n26702 13.653
R9877 vp_p.n25278 vp_p.n25277 13.653
R9878 vp_p.n23856 vp_p.n23855 13.653
R9879 vp_p.n22433 vp_p.n22432 13.653
R9880 vp_p.n21009 vp_p.n21008 13.653
R9881 vp_p.n19584 vp_p.n19583 13.653
R9882 vp_p.n18158 vp_p.n18157 13.653
R9883 vp_p.n16731 vp_p.n16730 13.653
R9884 vp_p.n15303 vp_p.n15302 13.653
R9885 vp_p.n13541 vp_p.n13540 13.653
R9886 vp_p.n13539 vp_p.n13538 13.653
R9887 vp_p.n7419 vp_p.n7418 13.653
R9888 vp_p.n5997 vp_p.n5996 13.653
R9889 vp_p.n4574 vp_p.n4573 13.653
R9890 vp_p.n3150 vp_p.n3149 13.653
R9891 vp_p.n1725 vp_p.n1724 13.653
R9892 vp_p.n241 vp_p.n240 13.653
R9893 vp_p.n8980 vp_p.n8979 13.653
R9894 vp_p.n10482 vp_p.n10481 13.653
R9895 vp_p.n11920 vp_p.n11919 13.653
R9896 vp_p.n26124 vp_p.n26123 13.653
R9897 vp_p.n24698 vp_p.n24697 13.653
R9898 vp_p.n23276 vp_p.n23275 13.653
R9899 vp_p.n21853 vp_p.n21852 13.653
R9900 vp_p.n20429 vp_p.n20428 13.653
R9901 vp_p.n19004 vp_p.n19003 13.653
R9902 vp_p.n17578 vp_p.n17577 13.653
R9903 vp_p.n16151 vp_p.n16150 13.653
R9904 vp_p.n14723 vp_p.n14722 13.653
R9905 vp_p.n13534 vp_p.n13533 13.653
R9906 vp_p.n8013 vp_p.n8012 13.653
R9907 vp_p.n6591 vp_p.n6590 13.653
R9908 vp_p.n5168 vp_p.n5167 13.653
R9909 vp_p.n3744 vp_p.n3743 13.653
R9910 vp_p.n2319 vp_p.n2318 13.653
R9911 vp_p.n893 vp_p.n892 13.653
R9912 vp_p.n9639 vp_p.n9638 13.653
R9913 vp_p.n11076 vp_p.n11075 13.653
R9914 vp_p.n12514 vp_p.n12513 13.653
R9915 vp_p.n26717 vp_p.n26716 13.653
R9916 vp_p.n25292 vp_p.n25291 13.653
R9917 vp_p.n23870 vp_p.n23869 13.653
R9918 vp_p.n22447 vp_p.n22446 13.653
R9919 vp_p.n21023 vp_p.n21022 13.653
R9920 vp_p.n19598 vp_p.n19597 13.653
R9921 vp_p.n18172 vp_p.n18171 13.653
R9922 vp_p.n16745 vp_p.n16744 13.653
R9923 vp_p.n15317 vp_p.n15316 13.653
R9924 vp_p.n13531 vp_p.n13530 13.653
R9925 vp_p.n13529 vp_p.n13528 13.653
R9926 vp_p.n7414 vp_p.n7413 13.653
R9927 vp_p.n5992 vp_p.n5991 13.653
R9928 vp_p.n4569 vp_p.n4568 13.653
R9929 vp_p.n3145 vp_p.n3144 13.653
R9930 vp_p.n1720 vp_p.n1719 13.653
R9931 vp_p.n236 vp_p.n235 13.653
R9932 vp_p.n8975 vp_p.n8974 13.653
R9933 vp_p.n10477 vp_p.n10476 13.653
R9934 vp_p.n11915 vp_p.n11914 13.653
R9935 vp_p.n26119 vp_p.n26118 13.653
R9936 vp_p.n24693 vp_p.n24692 13.653
R9937 vp_p.n23271 vp_p.n23270 13.653
R9938 vp_p.n21848 vp_p.n21847 13.653
R9939 vp_p.n20424 vp_p.n20423 13.653
R9940 vp_p.n18999 vp_p.n18998 13.653
R9941 vp_p.n17573 vp_p.n17572 13.653
R9942 vp_p.n16146 vp_p.n16145 13.653
R9943 vp_p.n14718 vp_p.n14717 13.653
R9944 vp_p.n13524 vp_p.n13523 13.653
R9945 vp_p.n8027 vp_p.n8026 13.653
R9946 vp_p.n6605 vp_p.n6604 13.653
R9947 vp_p.n5182 vp_p.n5181 13.653
R9948 vp_p.n3758 vp_p.n3757 13.653
R9949 vp_p.n2333 vp_p.n2332 13.653
R9950 vp_p.n907 vp_p.n906 13.653
R9951 vp_p.n9653 vp_p.n9652 13.653
R9952 vp_p.n11090 vp_p.n11089 13.653
R9953 vp_p.n12528 vp_p.n12527 13.653
R9954 vp_p.n26731 vp_p.n26730 13.653
R9955 vp_p.n25306 vp_p.n25305 13.653
R9956 vp_p.n23884 vp_p.n23883 13.653
R9957 vp_p.n22461 vp_p.n22460 13.653
R9958 vp_p.n21037 vp_p.n21036 13.653
R9959 vp_p.n19612 vp_p.n19611 13.653
R9960 vp_p.n18186 vp_p.n18185 13.653
R9961 vp_p.n16759 vp_p.n16758 13.653
R9962 vp_p.n15331 vp_p.n15330 13.653
R9963 vp_p.n13521 vp_p.n13520 13.653
R9964 vp_p.n13519 vp_p.n13518 13.653
R9965 vp_p.n7409 vp_p.n7408 13.653
R9966 vp_p.n5987 vp_p.n5986 13.653
R9967 vp_p.n4564 vp_p.n4563 13.653
R9968 vp_p.n3140 vp_p.n3139 13.653
R9969 vp_p.n1715 vp_p.n1714 13.653
R9970 vp_p.n231 vp_p.n230 13.653
R9971 vp_p.n8970 vp_p.n8969 13.653
R9972 vp_p.n10472 vp_p.n10471 13.653
R9973 vp_p.n11910 vp_p.n11909 13.653
R9974 vp_p.n26114 vp_p.n26113 13.653
R9975 vp_p.n24688 vp_p.n24687 13.653
R9976 vp_p.n23266 vp_p.n23265 13.653
R9977 vp_p.n21843 vp_p.n21842 13.653
R9978 vp_p.n20419 vp_p.n20418 13.653
R9979 vp_p.n18994 vp_p.n18993 13.653
R9980 vp_p.n17568 vp_p.n17567 13.653
R9981 vp_p.n16141 vp_p.n16140 13.653
R9982 vp_p.n14713 vp_p.n14712 13.653
R9983 vp_p.n13514 vp_p.n13513 13.653
R9984 vp_p.n8041 vp_p.n8040 13.653
R9985 vp_p.n6619 vp_p.n6618 13.653
R9986 vp_p.n5196 vp_p.n5195 13.653
R9987 vp_p.n3772 vp_p.n3771 13.653
R9988 vp_p.n2347 vp_p.n2346 13.653
R9989 vp_p.n921 vp_p.n920 13.653
R9990 vp_p.n9667 vp_p.n9666 13.653
R9991 vp_p.n11104 vp_p.n11103 13.653
R9992 vp_p.n12542 vp_p.n12541 13.653
R9993 vp_p.n26745 vp_p.n26744 13.653
R9994 vp_p.n25320 vp_p.n25319 13.653
R9995 vp_p.n23898 vp_p.n23897 13.653
R9996 vp_p.n22475 vp_p.n22474 13.653
R9997 vp_p.n21051 vp_p.n21050 13.653
R9998 vp_p.n19626 vp_p.n19625 13.653
R9999 vp_p.n18200 vp_p.n18199 13.653
R10000 vp_p.n16773 vp_p.n16772 13.653
R10001 vp_p.n15345 vp_p.n15344 13.653
R10002 vp_p.n13511 vp_p.n13510 13.653
R10003 vp_p.n13509 vp_p.n13508 13.653
R10004 vp_p.n7404 vp_p.n7403 13.653
R10005 vp_p.n5982 vp_p.n5981 13.653
R10006 vp_p.n4559 vp_p.n4558 13.653
R10007 vp_p.n3135 vp_p.n3134 13.653
R10008 vp_p.n1710 vp_p.n1709 13.653
R10009 vp_p.n226 vp_p.n225 13.653
R10010 vp_p.n8965 vp_p.n8964 13.653
R10011 vp_p.n10467 vp_p.n10466 13.653
R10012 vp_p.n11905 vp_p.n11904 13.653
R10013 vp_p.n26109 vp_p.n26108 13.653
R10014 vp_p.n24683 vp_p.n24682 13.653
R10015 vp_p.n23261 vp_p.n23260 13.653
R10016 vp_p.n21838 vp_p.n21837 13.653
R10017 vp_p.n20414 vp_p.n20413 13.653
R10018 vp_p.n18989 vp_p.n18988 13.653
R10019 vp_p.n17563 vp_p.n17562 13.653
R10020 vp_p.n16136 vp_p.n16135 13.653
R10021 vp_p.n14708 vp_p.n14707 13.653
R10022 vp_p.n13504 vp_p.n13503 13.653
R10023 vp_p.n8055 vp_p.n8054 13.653
R10024 vp_p.n6633 vp_p.n6632 13.653
R10025 vp_p.n5210 vp_p.n5209 13.653
R10026 vp_p.n3786 vp_p.n3785 13.653
R10027 vp_p.n2361 vp_p.n2360 13.653
R10028 vp_p.n935 vp_p.n934 13.653
R10029 vp_p.n9681 vp_p.n9680 13.653
R10030 vp_p.n11118 vp_p.n11117 13.653
R10031 vp_p.n12556 vp_p.n12555 13.653
R10032 vp_p.n26759 vp_p.n26758 13.653
R10033 vp_p.n25334 vp_p.n25333 13.653
R10034 vp_p.n23912 vp_p.n23911 13.653
R10035 vp_p.n22489 vp_p.n22488 13.653
R10036 vp_p.n21065 vp_p.n21064 13.653
R10037 vp_p.n19640 vp_p.n19639 13.653
R10038 vp_p.n18214 vp_p.n18213 13.653
R10039 vp_p.n16787 vp_p.n16786 13.653
R10040 vp_p.n15359 vp_p.n15358 13.653
R10041 vp_p.n13501 vp_p.n13500 13.653
R10042 vp_p.n13499 vp_p.n13498 13.653
R10043 vp_p.n7399 vp_p.n7398 13.653
R10044 vp_p.n5977 vp_p.n5976 13.653
R10045 vp_p.n4554 vp_p.n4553 13.653
R10046 vp_p.n3130 vp_p.n3129 13.653
R10047 vp_p.n1705 vp_p.n1704 13.653
R10048 vp_p.n221 vp_p.n220 13.653
R10049 vp_p.n8960 vp_p.n8959 13.653
R10050 vp_p.n10462 vp_p.n10461 13.653
R10051 vp_p.n11900 vp_p.n11899 13.653
R10052 vp_p.n26104 vp_p.n26103 13.653
R10053 vp_p.n24678 vp_p.n24677 13.653
R10054 vp_p.n23256 vp_p.n23255 13.653
R10055 vp_p.n21833 vp_p.n21832 13.653
R10056 vp_p.n20409 vp_p.n20408 13.653
R10057 vp_p.n18984 vp_p.n18983 13.653
R10058 vp_p.n17558 vp_p.n17557 13.653
R10059 vp_p.n16131 vp_p.n16130 13.653
R10060 vp_p.n14703 vp_p.n14702 13.653
R10061 vp_p.n13494 vp_p.n13493 13.653
R10062 vp_p.n8069 vp_p.n8068 13.653
R10063 vp_p.n6647 vp_p.n6646 13.653
R10064 vp_p.n5224 vp_p.n5223 13.653
R10065 vp_p.n3800 vp_p.n3799 13.653
R10066 vp_p.n2375 vp_p.n2374 13.653
R10067 vp_p.n949 vp_p.n948 13.653
R10068 vp_p.n9695 vp_p.n9694 13.653
R10069 vp_p.n11132 vp_p.n11131 13.653
R10070 vp_p.n12570 vp_p.n12569 13.653
R10071 vp_p.n26773 vp_p.n26772 13.653
R10072 vp_p.n25348 vp_p.n25347 13.653
R10073 vp_p.n23926 vp_p.n23925 13.653
R10074 vp_p.n22503 vp_p.n22502 13.653
R10075 vp_p.n21079 vp_p.n21078 13.653
R10076 vp_p.n19654 vp_p.n19653 13.653
R10077 vp_p.n18228 vp_p.n18227 13.653
R10078 vp_p.n16801 vp_p.n16800 13.653
R10079 vp_p.n15373 vp_p.n15372 13.653
R10080 vp_p.n13491 vp_p.n13490 13.653
R10081 vp_p.n13489 vp_p.n13488 13.653
R10082 vp_p.n7394 vp_p.n7393 13.653
R10083 vp_p.n5972 vp_p.n5971 13.653
R10084 vp_p.n4549 vp_p.n4548 13.653
R10085 vp_p.n3125 vp_p.n3124 13.653
R10086 vp_p.n1700 vp_p.n1699 13.653
R10087 vp_p.n216 vp_p.n215 13.653
R10088 vp_p.n8955 vp_p.n8954 13.653
R10089 vp_p.n10457 vp_p.n10456 13.653
R10090 vp_p.n11895 vp_p.n11894 13.653
R10091 vp_p.n26099 vp_p.n26098 13.653
R10092 vp_p.n24673 vp_p.n24672 13.653
R10093 vp_p.n23251 vp_p.n23250 13.653
R10094 vp_p.n21828 vp_p.n21827 13.653
R10095 vp_p.n20404 vp_p.n20403 13.653
R10096 vp_p.n18979 vp_p.n18978 13.653
R10097 vp_p.n17553 vp_p.n17552 13.653
R10098 vp_p.n16126 vp_p.n16125 13.653
R10099 vp_p.n14698 vp_p.n14697 13.653
R10100 vp_p.n13484 vp_p.n13483 13.653
R10101 vp_p.n8083 vp_p.n8082 13.653
R10102 vp_p.n6661 vp_p.n6660 13.653
R10103 vp_p.n5238 vp_p.n5237 13.653
R10104 vp_p.n3814 vp_p.n3813 13.653
R10105 vp_p.n2389 vp_p.n2388 13.653
R10106 vp_p.n963 vp_p.n962 13.653
R10107 vp_p.n9709 vp_p.n9708 13.653
R10108 vp_p.n11146 vp_p.n11145 13.653
R10109 vp_p.n12584 vp_p.n12583 13.653
R10110 vp_p.n26787 vp_p.n26786 13.653
R10111 vp_p.n25362 vp_p.n25361 13.653
R10112 vp_p.n23940 vp_p.n23939 13.653
R10113 vp_p.n22517 vp_p.n22516 13.653
R10114 vp_p.n21093 vp_p.n21092 13.653
R10115 vp_p.n19668 vp_p.n19667 13.653
R10116 vp_p.n18242 vp_p.n18241 13.653
R10117 vp_p.n16815 vp_p.n16814 13.653
R10118 vp_p.n15387 vp_p.n15386 13.653
R10119 vp_p.n13481 vp_p.n13480 13.653
R10120 vp_p.n13479 vp_p.n13478 13.653
R10121 vp_p.n7389 vp_p.n7388 13.653
R10122 vp_p.n5967 vp_p.n5966 13.653
R10123 vp_p.n4544 vp_p.n4543 13.653
R10124 vp_p.n3120 vp_p.n3119 13.653
R10125 vp_p.n1695 vp_p.n1694 13.653
R10126 vp_p.n211 vp_p.n210 13.653
R10127 vp_p.n8950 vp_p.n8949 13.653
R10128 vp_p.n10452 vp_p.n10451 13.653
R10129 vp_p.n11890 vp_p.n11889 13.653
R10130 vp_p.n26094 vp_p.n26093 13.653
R10131 vp_p.n24668 vp_p.n24667 13.653
R10132 vp_p.n23246 vp_p.n23245 13.653
R10133 vp_p.n21823 vp_p.n21822 13.653
R10134 vp_p.n20399 vp_p.n20398 13.653
R10135 vp_p.n18974 vp_p.n18973 13.653
R10136 vp_p.n17548 vp_p.n17547 13.653
R10137 vp_p.n16121 vp_p.n16120 13.653
R10138 vp_p.n14693 vp_p.n14692 13.653
R10139 vp_p.n13474 vp_p.n13473 13.653
R10140 vp_p.n8097 vp_p.n8096 13.653
R10141 vp_p.n6675 vp_p.n6674 13.653
R10142 vp_p.n5252 vp_p.n5251 13.653
R10143 vp_p.n3828 vp_p.n3827 13.653
R10144 vp_p.n2403 vp_p.n2402 13.653
R10145 vp_p.n977 vp_p.n976 13.653
R10146 vp_p.n9723 vp_p.n9722 13.653
R10147 vp_p.n11160 vp_p.n11159 13.653
R10148 vp_p.n12598 vp_p.n12597 13.653
R10149 vp_p.n26801 vp_p.n26800 13.653
R10150 vp_p.n25376 vp_p.n25375 13.653
R10151 vp_p.n23954 vp_p.n23953 13.653
R10152 vp_p.n22531 vp_p.n22530 13.653
R10153 vp_p.n21107 vp_p.n21106 13.653
R10154 vp_p.n19682 vp_p.n19681 13.653
R10155 vp_p.n18256 vp_p.n18255 13.653
R10156 vp_p.n16829 vp_p.n16828 13.653
R10157 vp_p.n15401 vp_p.n15400 13.653
R10158 vp_p.n13471 vp_p.n13470 13.653
R10159 vp_p.n13469 vp_p.n13468 13.653
R10160 vp_p.n7384 vp_p.n7383 13.653
R10161 vp_p.n5962 vp_p.n5961 13.653
R10162 vp_p.n4539 vp_p.n4538 13.653
R10163 vp_p.n3115 vp_p.n3114 13.653
R10164 vp_p.n1690 vp_p.n1689 13.653
R10165 vp_p.n206 vp_p.n205 13.653
R10166 vp_p.n8945 vp_p.n8944 13.653
R10167 vp_p.n10447 vp_p.n10446 13.653
R10168 vp_p.n11885 vp_p.n11884 13.653
R10169 vp_p.n26089 vp_p.n26088 13.653
R10170 vp_p.n24663 vp_p.n24662 13.653
R10171 vp_p.n23241 vp_p.n23240 13.653
R10172 vp_p.n21818 vp_p.n21817 13.653
R10173 vp_p.n20394 vp_p.n20393 13.653
R10174 vp_p.n18969 vp_p.n18968 13.653
R10175 vp_p.n17543 vp_p.n17542 13.653
R10176 vp_p.n16116 vp_p.n16115 13.653
R10177 vp_p.n14688 vp_p.n14687 13.653
R10178 vp_p.n13464 vp_p.n13463 13.653
R10179 vp_p.n8111 vp_p.n8110 13.653
R10180 vp_p.n6689 vp_p.n6688 13.653
R10181 vp_p.n5266 vp_p.n5265 13.653
R10182 vp_p.n3842 vp_p.n3841 13.653
R10183 vp_p.n2417 vp_p.n2416 13.653
R10184 vp_p.n991 vp_p.n990 13.653
R10185 vp_p.n9737 vp_p.n9736 13.653
R10186 vp_p.n11174 vp_p.n11173 13.653
R10187 vp_p.n12612 vp_p.n12611 13.653
R10188 vp_p.n26815 vp_p.n26814 13.653
R10189 vp_p.n25390 vp_p.n25389 13.653
R10190 vp_p.n23968 vp_p.n23967 13.653
R10191 vp_p.n22545 vp_p.n22544 13.653
R10192 vp_p.n21121 vp_p.n21120 13.653
R10193 vp_p.n19696 vp_p.n19695 13.653
R10194 vp_p.n18270 vp_p.n18269 13.653
R10195 vp_p.n16843 vp_p.n16842 13.653
R10196 vp_p.n15415 vp_p.n15414 13.653
R10197 vp_p.n13461 vp_p.n13460 13.653
R10198 vp_p.n13459 vp_p.n13458 13.653
R10199 vp_p.n7379 vp_p.n7378 13.653
R10200 vp_p.n5957 vp_p.n5956 13.653
R10201 vp_p.n4534 vp_p.n4533 13.653
R10202 vp_p.n3110 vp_p.n3109 13.653
R10203 vp_p.n1685 vp_p.n1684 13.653
R10204 vp_p.n201 vp_p.n200 13.653
R10205 vp_p.n8940 vp_p.n8939 13.653
R10206 vp_p.n10442 vp_p.n10441 13.653
R10207 vp_p.n11880 vp_p.n11879 13.653
R10208 vp_p.n26084 vp_p.n26083 13.653
R10209 vp_p.n24658 vp_p.n24657 13.653
R10210 vp_p.n23236 vp_p.n23235 13.653
R10211 vp_p.n21813 vp_p.n21812 13.653
R10212 vp_p.n20389 vp_p.n20388 13.653
R10213 vp_p.n18964 vp_p.n18963 13.653
R10214 vp_p.n17538 vp_p.n17537 13.653
R10215 vp_p.n16111 vp_p.n16110 13.653
R10216 vp_p.n14683 vp_p.n14682 13.653
R10217 vp_p.n13454 vp_p.n13453 13.653
R10218 vp_p.n8125 vp_p.n8124 13.653
R10219 vp_p.n6703 vp_p.n6702 13.653
R10220 vp_p.n5280 vp_p.n5279 13.653
R10221 vp_p.n3856 vp_p.n3855 13.653
R10222 vp_p.n2431 vp_p.n2430 13.653
R10223 vp_p.n1005 vp_p.n1004 13.653
R10224 vp_p.n9751 vp_p.n9750 13.653
R10225 vp_p.n11188 vp_p.n11187 13.653
R10226 vp_p.n12626 vp_p.n12625 13.653
R10227 vp_p.n26829 vp_p.n26828 13.653
R10228 vp_p.n25404 vp_p.n25403 13.653
R10229 vp_p.n23982 vp_p.n23981 13.653
R10230 vp_p.n22559 vp_p.n22558 13.653
R10231 vp_p.n21135 vp_p.n21134 13.653
R10232 vp_p.n19710 vp_p.n19709 13.653
R10233 vp_p.n18284 vp_p.n18283 13.653
R10234 vp_p.n16857 vp_p.n16856 13.653
R10235 vp_p.n15429 vp_p.n15428 13.653
R10236 vp_p.n13451 vp_p.n13450 13.653
R10237 vp_p.n13449 vp_p.n13448 13.653
R10238 vp_p.n7374 vp_p.n7373 13.653
R10239 vp_p.n5952 vp_p.n5951 13.653
R10240 vp_p.n4529 vp_p.n4528 13.653
R10241 vp_p.n3105 vp_p.n3104 13.653
R10242 vp_p.n1680 vp_p.n1679 13.653
R10243 vp_p.n196 vp_p.n195 13.653
R10244 vp_p.n8935 vp_p.n8934 13.653
R10245 vp_p.n10437 vp_p.n10436 13.653
R10246 vp_p.n11875 vp_p.n11874 13.653
R10247 vp_p.n26079 vp_p.n26078 13.653
R10248 vp_p.n24653 vp_p.n24652 13.653
R10249 vp_p.n23231 vp_p.n23230 13.653
R10250 vp_p.n21808 vp_p.n21807 13.653
R10251 vp_p.n20384 vp_p.n20383 13.653
R10252 vp_p.n18959 vp_p.n18958 13.653
R10253 vp_p.n17533 vp_p.n17532 13.653
R10254 vp_p.n16106 vp_p.n16105 13.653
R10255 vp_p.n14678 vp_p.n14677 13.653
R10256 vp_p.n13444 vp_p.n13443 13.653
R10257 vp_p.n8139 vp_p.n8138 13.653
R10258 vp_p.n6717 vp_p.n6716 13.653
R10259 vp_p.n5294 vp_p.n5293 13.653
R10260 vp_p.n3870 vp_p.n3869 13.653
R10261 vp_p.n2445 vp_p.n2444 13.653
R10262 vp_p.n1019 vp_p.n1018 13.653
R10263 vp_p.n9765 vp_p.n9764 13.653
R10264 vp_p.n11202 vp_p.n11201 13.653
R10265 vp_p.n12640 vp_p.n12639 13.653
R10266 vp_p.n26843 vp_p.n26842 13.653
R10267 vp_p.n25418 vp_p.n25417 13.653
R10268 vp_p.n23996 vp_p.n23995 13.653
R10269 vp_p.n22573 vp_p.n22572 13.653
R10270 vp_p.n21149 vp_p.n21148 13.653
R10271 vp_p.n19724 vp_p.n19723 13.653
R10272 vp_p.n18298 vp_p.n18297 13.653
R10273 vp_p.n16871 vp_p.n16870 13.653
R10274 vp_p.n15443 vp_p.n15442 13.653
R10275 vp_p.n13441 vp_p.n13440 13.653
R10276 vp_p.n13439 vp_p.n13438 13.653
R10277 vp_p.n7369 vp_p.n7368 13.653
R10278 vp_p.n5947 vp_p.n5946 13.653
R10279 vp_p.n4524 vp_p.n4523 13.653
R10280 vp_p.n3100 vp_p.n3099 13.653
R10281 vp_p.n1675 vp_p.n1674 13.653
R10282 vp_p.n191 vp_p.n190 13.653
R10283 vp_p.n8930 vp_p.n8929 13.653
R10284 vp_p.n10432 vp_p.n10431 13.653
R10285 vp_p.n11870 vp_p.n11869 13.653
R10286 vp_p.n26074 vp_p.n26073 13.653
R10287 vp_p.n24648 vp_p.n24647 13.653
R10288 vp_p.n23226 vp_p.n23225 13.653
R10289 vp_p.n21803 vp_p.n21802 13.653
R10290 vp_p.n20379 vp_p.n20378 13.653
R10291 vp_p.n18954 vp_p.n18953 13.653
R10292 vp_p.n17528 vp_p.n17527 13.653
R10293 vp_p.n16101 vp_p.n16100 13.653
R10294 vp_p.n14673 vp_p.n14672 13.653
R10295 vp_p.n13434 vp_p.n13433 13.653
R10296 vp_p.n8153 vp_p.n8152 13.653
R10297 vp_p.n6731 vp_p.n6730 13.653
R10298 vp_p.n5308 vp_p.n5307 13.653
R10299 vp_p.n3884 vp_p.n3883 13.653
R10300 vp_p.n2459 vp_p.n2458 13.653
R10301 vp_p.n1033 vp_p.n1032 13.653
R10302 vp_p.n9779 vp_p.n9778 13.653
R10303 vp_p.n11216 vp_p.n11215 13.653
R10304 vp_p.n12654 vp_p.n12653 13.653
R10305 vp_p.n26857 vp_p.n26856 13.653
R10306 vp_p.n25432 vp_p.n25431 13.653
R10307 vp_p.n24010 vp_p.n24009 13.653
R10308 vp_p.n22587 vp_p.n22586 13.653
R10309 vp_p.n21163 vp_p.n21162 13.653
R10310 vp_p.n19738 vp_p.n19737 13.653
R10311 vp_p.n18312 vp_p.n18311 13.653
R10312 vp_p.n16885 vp_p.n16884 13.653
R10313 vp_p.n15457 vp_p.n15456 13.653
R10314 vp_p.n13431 vp_p.n13430 13.653
R10315 vp_p.n13429 vp_p.n13428 13.653
R10316 vp_p.n7364 vp_p.n7363 13.653
R10317 vp_p.n5942 vp_p.n5941 13.653
R10318 vp_p.n4519 vp_p.n4518 13.653
R10319 vp_p.n3095 vp_p.n3094 13.653
R10320 vp_p.n1670 vp_p.n1669 13.653
R10321 vp_p.n186 vp_p.n185 13.653
R10322 vp_p.n8925 vp_p.n8924 13.653
R10323 vp_p.n10427 vp_p.n10426 13.653
R10324 vp_p.n11865 vp_p.n11864 13.653
R10325 vp_p.n26069 vp_p.n26068 13.653
R10326 vp_p.n24643 vp_p.n24642 13.653
R10327 vp_p.n23221 vp_p.n23220 13.653
R10328 vp_p.n21798 vp_p.n21797 13.653
R10329 vp_p.n20374 vp_p.n20373 13.653
R10330 vp_p.n18949 vp_p.n18948 13.653
R10331 vp_p.n17523 vp_p.n17522 13.653
R10332 vp_p.n16096 vp_p.n16095 13.653
R10333 vp_p.n14668 vp_p.n14667 13.653
R10334 vp_p.n13424 vp_p.n13423 13.653
R10335 vp_p.n8167 vp_p.n8166 13.653
R10336 vp_p.n6745 vp_p.n6744 13.653
R10337 vp_p.n5322 vp_p.n5321 13.653
R10338 vp_p.n3898 vp_p.n3897 13.653
R10339 vp_p.n2473 vp_p.n2472 13.653
R10340 vp_p.n1047 vp_p.n1046 13.653
R10341 vp_p.n9793 vp_p.n9792 13.653
R10342 vp_p.n11230 vp_p.n11229 13.653
R10343 vp_p.n12668 vp_p.n12667 13.653
R10344 vp_p.n26871 vp_p.n26870 13.653
R10345 vp_p.n25446 vp_p.n25445 13.653
R10346 vp_p.n24024 vp_p.n24023 13.653
R10347 vp_p.n22601 vp_p.n22600 13.653
R10348 vp_p.n21177 vp_p.n21176 13.653
R10349 vp_p.n19752 vp_p.n19751 13.653
R10350 vp_p.n18326 vp_p.n18325 13.653
R10351 vp_p.n16899 vp_p.n16898 13.653
R10352 vp_p.n15471 vp_p.n15470 13.653
R10353 vp_p.n13421 vp_p.n13420 13.653
R10354 vp_p.n13419 vp_p.n13418 13.653
R10355 vp_p.n7359 vp_p.n7358 13.653
R10356 vp_p.n5937 vp_p.n5936 13.653
R10357 vp_p.n4514 vp_p.n4513 13.653
R10358 vp_p.n3090 vp_p.n3089 13.653
R10359 vp_p.n1665 vp_p.n1664 13.653
R10360 vp_p.n181 vp_p.n180 13.653
R10361 vp_p.n8920 vp_p.n8919 13.653
R10362 vp_p.n10422 vp_p.n10421 13.653
R10363 vp_p.n11860 vp_p.n11859 13.653
R10364 vp_p.n26064 vp_p.n26063 13.653
R10365 vp_p.n24638 vp_p.n24637 13.653
R10366 vp_p.n23216 vp_p.n23215 13.653
R10367 vp_p.n21793 vp_p.n21792 13.653
R10368 vp_p.n20369 vp_p.n20368 13.653
R10369 vp_p.n18944 vp_p.n18943 13.653
R10370 vp_p.n17518 vp_p.n17517 13.653
R10371 vp_p.n16091 vp_p.n16090 13.653
R10372 vp_p.n14663 vp_p.n14662 13.653
R10373 vp_p.n13414 vp_p.n13413 13.653
R10374 vp_p.n8181 vp_p.n8180 13.653
R10375 vp_p.n6759 vp_p.n6758 13.653
R10376 vp_p.n5336 vp_p.n5335 13.653
R10377 vp_p.n3912 vp_p.n3911 13.653
R10378 vp_p.n2487 vp_p.n2486 13.653
R10379 vp_p.n1061 vp_p.n1060 13.653
R10380 vp_p.n9807 vp_p.n9806 13.653
R10381 vp_p.n11244 vp_p.n11243 13.653
R10382 vp_p.n12682 vp_p.n12681 13.653
R10383 vp_p.n26885 vp_p.n26884 13.653
R10384 vp_p.n25460 vp_p.n25459 13.653
R10385 vp_p.n24038 vp_p.n24037 13.653
R10386 vp_p.n22615 vp_p.n22614 13.653
R10387 vp_p.n21191 vp_p.n21190 13.653
R10388 vp_p.n19766 vp_p.n19765 13.653
R10389 vp_p.n18340 vp_p.n18339 13.653
R10390 vp_p.n16913 vp_p.n16912 13.653
R10391 vp_p.n15485 vp_p.n15484 13.653
R10392 vp_p.n13411 vp_p.n13410 13.653
R10393 vp_p.n13409 vp_p.n13408 13.653
R10394 vp_p.n7354 vp_p.n7353 13.653
R10395 vp_p.n5932 vp_p.n5931 13.653
R10396 vp_p.n4509 vp_p.n4508 13.653
R10397 vp_p.n3085 vp_p.n3084 13.653
R10398 vp_p.n1660 vp_p.n1659 13.653
R10399 vp_p.n176 vp_p.n175 13.653
R10400 vp_p.n8915 vp_p.n8914 13.653
R10401 vp_p.n10417 vp_p.n10416 13.653
R10402 vp_p.n11855 vp_p.n11854 13.653
R10403 vp_p.n26059 vp_p.n26058 13.653
R10404 vp_p.n24633 vp_p.n24632 13.653
R10405 vp_p.n23211 vp_p.n23210 13.653
R10406 vp_p.n21788 vp_p.n21787 13.653
R10407 vp_p.n20364 vp_p.n20363 13.653
R10408 vp_p.n18939 vp_p.n18938 13.653
R10409 vp_p.n17513 vp_p.n17512 13.653
R10410 vp_p.n16086 vp_p.n16085 13.653
R10411 vp_p.n14658 vp_p.n14657 13.653
R10412 vp_p.n13404 vp_p.n13403 13.653
R10413 vp_p.n8195 vp_p.n8194 13.653
R10414 vp_p.n6773 vp_p.n6772 13.653
R10415 vp_p.n5350 vp_p.n5349 13.653
R10416 vp_p.n3926 vp_p.n3925 13.653
R10417 vp_p.n2501 vp_p.n2500 13.653
R10418 vp_p.n1075 vp_p.n1074 13.653
R10419 vp_p.n9821 vp_p.n9820 13.653
R10420 vp_p.n11258 vp_p.n11257 13.653
R10421 vp_p.n12696 vp_p.n12695 13.653
R10422 vp_p.n26899 vp_p.n26898 13.653
R10423 vp_p.n25474 vp_p.n25473 13.653
R10424 vp_p.n24052 vp_p.n24051 13.653
R10425 vp_p.n22629 vp_p.n22628 13.653
R10426 vp_p.n21205 vp_p.n21204 13.653
R10427 vp_p.n19780 vp_p.n19779 13.653
R10428 vp_p.n18354 vp_p.n18353 13.653
R10429 vp_p.n16927 vp_p.n16926 13.653
R10430 vp_p.n15499 vp_p.n15498 13.653
R10431 vp_p.n13401 vp_p.n13400 13.653
R10432 vp_p.n13399 vp_p.n13398 13.653
R10433 vp_p.n7349 vp_p.n7348 13.653
R10434 vp_p.n5927 vp_p.n5926 13.653
R10435 vp_p.n4504 vp_p.n4503 13.653
R10436 vp_p.n3080 vp_p.n3079 13.653
R10437 vp_p.n1655 vp_p.n1654 13.653
R10438 vp_p.n171 vp_p.n170 13.653
R10439 vp_p.n8910 vp_p.n8909 13.653
R10440 vp_p.n10412 vp_p.n10411 13.653
R10441 vp_p.n11850 vp_p.n11849 13.653
R10442 vp_p.n26054 vp_p.n26053 13.653
R10443 vp_p.n24628 vp_p.n24627 13.653
R10444 vp_p.n23206 vp_p.n23205 13.653
R10445 vp_p.n21783 vp_p.n21782 13.653
R10446 vp_p.n20359 vp_p.n20358 13.653
R10447 vp_p.n18934 vp_p.n18933 13.653
R10448 vp_p.n17508 vp_p.n17507 13.653
R10449 vp_p.n16081 vp_p.n16080 13.653
R10450 vp_p.n14653 vp_p.n14652 13.653
R10451 vp_p.n13394 vp_p.n13393 13.653
R10452 vp_p.n8209 vp_p.n8208 13.653
R10453 vp_p.n6787 vp_p.n6786 13.653
R10454 vp_p.n5364 vp_p.n5363 13.653
R10455 vp_p.n3940 vp_p.n3939 13.653
R10456 vp_p.n2515 vp_p.n2514 13.653
R10457 vp_p.n1089 vp_p.n1088 13.653
R10458 vp_p.n9835 vp_p.n9834 13.653
R10459 vp_p.n11272 vp_p.n11271 13.653
R10460 vp_p.n12710 vp_p.n12709 13.653
R10461 vp_p.n26913 vp_p.n26912 13.653
R10462 vp_p.n25488 vp_p.n25487 13.653
R10463 vp_p.n24066 vp_p.n24065 13.653
R10464 vp_p.n22643 vp_p.n22642 13.653
R10465 vp_p.n21219 vp_p.n21218 13.653
R10466 vp_p.n19794 vp_p.n19793 13.653
R10467 vp_p.n18368 vp_p.n18367 13.653
R10468 vp_p.n16941 vp_p.n16940 13.653
R10469 vp_p.n15513 vp_p.n15512 13.653
R10470 vp_p.n13391 vp_p.n13390 13.653
R10471 vp_p.n13389 vp_p.n13388 13.653
R10472 vp_p.n7344 vp_p.n7343 13.653
R10473 vp_p.n5922 vp_p.n5921 13.653
R10474 vp_p.n4499 vp_p.n4498 13.653
R10475 vp_p.n3075 vp_p.n3074 13.653
R10476 vp_p.n1650 vp_p.n1649 13.653
R10477 vp_p.n166 vp_p.n165 13.653
R10478 vp_p.n8905 vp_p.n8904 13.653
R10479 vp_p.n10407 vp_p.n10406 13.653
R10480 vp_p.n11845 vp_p.n11844 13.653
R10481 vp_p.n26049 vp_p.n26048 13.653
R10482 vp_p.n24623 vp_p.n24622 13.653
R10483 vp_p.n23201 vp_p.n23200 13.653
R10484 vp_p.n21778 vp_p.n21777 13.653
R10485 vp_p.n20354 vp_p.n20353 13.653
R10486 vp_p.n18929 vp_p.n18928 13.653
R10487 vp_p.n17503 vp_p.n17502 13.653
R10488 vp_p.n16076 vp_p.n16075 13.653
R10489 vp_p.n14648 vp_p.n14647 13.653
R10490 vp_p.n13384 vp_p.n13383 13.653
R10491 vp_p.n8223 vp_p.n8222 13.653
R10492 vp_p.n6801 vp_p.n6800 13.653
R10493 vp_p.n5378 vp_p.n5377 13.653
R10494 vp_p.n3954 vp_p.n3953 13.653
R10495 vp_p.n2529 vp_p.n2528 13.653
R10496 vp_p.n1103 vp_p.n1102 13.653
R10497 vp_p.n9849 vp_p.n9848 13.653
R10498 vp_p.n11286 vp_p.n11285 13.653
R10499 vp_p.n12724 vp_p.n12723 13.653
R10500 vp_p.n26927 vp_p.n26926 13.653
R10501 vp_p.n25502 vp_p.n25501 13.653
R10502 vp_p.n24080 vp_p.n24079 13.653
R10503 vp_p.n22657 vp_p.n22656 13.653
R10504 vp_p.n21233 vp_p.n21232 13.653
R10505 vp_p.n19808 vp_p.n19807 13.653
R10506 vp_p.n18382 vp_p.n18381 13.653
R10507 vp_p.n16955 vp_p.n16954 13.653
R10508 vp_p.n15527 vp_p.n15526 13.653
R10509 vp_p.n13381 vp_p.n13380 13.653
R10510 vp_p.n13379 vp_p.n13378 13.653
R10511 vp_p.n7339 vp_p.n7338 13.653
R10512 vp_p.n5917 vp_p.n5916 13.653
R10513 vp_p.n4494 vp_p.n4493 13.653
R10514 vp_p.n3070 vp_p.n3069 13.653
R10515 vp_p.n1645 vp_p.n1644 13.653
R10516 vp_p.n161 vp_p.n160 13.653
R10517 vp_p.n8900 vp_p.n8899 13.653
R10518 vp_p.n10402 vp_p.n10401 13.653
R10519 vp_p.n11840 vp_p.n11839 13.653
R10520 vp_p.n26044 vp_p.n26043 13.653
R10521 vp_p.n24618 vp_p.n24617 13.653
R10522 vp_p.n23196 vp_p.n23195 13.653
R10523 vp_p.n21773 vp_p.n21772 13.653
R10524 vp_p.n20349 vp_p.n20348 13.653
R10525 vp_p.n18924 vp_p.n18923 13.653
R10526 vp_p.n17498 vp_p.n17497 13.653
R10527 vp_p.n16071 vp_p.n16070 13.653
R10528 vp_p.n14643 vp_p.n14642 13.653
R10529 vp_p.n13374 vp_p.n13373 13.653
R10530 vp_p.n8237 vp_p.n8236 13.653
R10531 vp_p.n6815 vp_p.n6814 13.653
R10532 vp_p.n5392 vp_p.n5391 13.653
R10533 vp_p.n3968 vp_p.n3967 13.653
R10534 vp_p.n2543 vp_p.n2542 13.653
R10535 vp_p.n1117 vp_p.n1116 13.653
R10536 vp_p.n9863 vp_p.n9862 13.653
R10537 vp_p.n11300 vp_p.n11299 13.653
R10538 vp_p.n12738 vp_p.n12737 13.653
R10539 vp_p.n26941 vp_p.n26940 13.653
R10540 vp_p.n25516 vp_p.n25515 13.653
R10541 vp_p.n24094 vp_p.n24093 13.653
R10542 vp_p.n22671 vp_p.n22670 13.653
R10543 vp_p.n21247 vp_p.n21246 13.653
R10544 vp_p.n19822 vp_p.n19821 13.653
R10545 vp_p.n18396 vp_p.n18395 13.653
R10546 vp_p.n16969 vp_p.n16968 13.653
R10547 vp_p.n15541 vp_p.n15540 13.653
R10548 vp_p.n13371 vp_p.n13370 13.653
R10549 vp_p.n13369 vp_p.n13368 13.653
R10550 vp_p.n7334 vp_p.n7333 13.653
R10551 vp_p.n5912 vp_p.n5911 13.653
R10552 vp_p.n4489 vp_p.n4488 13.653
R10553 vp_p.n3065 vp_p.n3064 13.653
R10554 vp_p.n1640 vp_p.n1639 13.653
R10555 vp_p.n156 vp_p.n155 13.653
R10556 vp_p.n8895 vp_p.n8894 13.653
R10557 vp_p.n10397 vp_p.n10396 13.653
R10558 vp_p.n11835 vp_p.n11834 13.653
R10559 vp_p.n26039 vp_p.n26038 13.653
R10560 vp_p.n24613 vp_p.n24612 13.653
R10561 vp_p.n23191 vp_p.n23190 13.653
R10562 vp_p.n21768 vp_p.n21767 13.653
R10563 vp_p.n20344 vp_p.n20343 13.653
R10564 vp_p.n18919 vp_p.n18918 13.653
R10565 vp_p.n17493 vp_p.n17492 13.653
R10566 vp_p.n16066 vp_p.n16065 13.653
R10567 vp_p.n14638 vp_p.n14637 13.653
R10568 vp_p.n13364 vp_p.n13363 13.653
R10569 vp_p.n8251 vp_p.n8250 13.653
R10570 vp_p.n6829 vp_p.n6828 13.653
R10571 vp_p.n5406 vp_p.n5405 13.653
R10572 vp_p.n3982 vp_p.n3981 13.653
R10573 vp_p.n2557 vp_p.n2556 13.653
R10574 vp_p.n1131 vp_p.n1130 13.653
R10575 vp_p.n9877 vp_p.n9876 13.653
R10576 vp_p.n11314 vp_p.n11313 13.653
R10577 vp_p.n12752 vp_p.n12751 13.653
R10578 vp_p.n26955 vp_p.n26954 13.653
R10579 vp_p.n25530 vp_p.n25529 13.653
R10580 vp_p.n24108 vp_p.n24107 13.653
R10581 vp_p.n22685 vp_p.n22684 13.653
R10582 vp_p.n21261 vp_p.n21260 13.653
R10583 vp_p.n19836 vp_p.n19835 13.653
R10584 vp_p.n18410 vp_p.n18409 13.653
R10585 vp_p.n16983 vp_p.n16982 13.653
R10586 vp_p.n15555 vp_p.n15554 13.653
R10587 vp_p.n13361 vp_p.n13360 13.653
R10588 vp_p.n13359 vp_p.n13358 13.653
R10589 vp_p.n7329 vp_p.n7328 13.653
R10590 vp_p.n5907 vp_p.n5906 13.653
R10591 vp_p.n4484 vp_p.n4483 13.653
R10592 vp_p.n3060 vp_p.n3059 13.653
R10593 vp_p.n1635 vp_p.n1634 13.653
R10594 vp_p.n151 vp_p.n150 13.653
R10595 vp_p.n8890 vp_p.n8889 13.653
R10596 vp_p.n10392 vp_p.n10391 13.653
R10597 vp_p.n11830 vp_p.n11829 13.653
R10598 vp_p.n26034 vp_p.n26033 13.653
R10599 vp_p.n24608 vp_p.n24607 13.653
R10600 vp_p.n23186 vp_p.n23185 13.653
R10601 vp_p.n21763 vp_p.n21762 13.653
R10602 vp_p.n20339 vp_p.n20338 13.653
R10603 vp_p.n18914 vp_p.n18913 13.653
R10604 vp_p.n17488 vp_p.n17487 13.653
R10605 vp_p.n16061 vp_p.n16060 13.653
R10606 vp_p.n14633 vp_p.n14632 13.653
R10607 vp_p.n13354 vp_p.n13353 13.653
R10608 vp_p.n8265 vp_p.n8264 13.653
R10609 vp_p.n6843 vp_p.n6842 13.653
R10610 vp_p.n5420 vp_p.n5419 13.653
R10611 vp_p.n3996 vp_p.n3995 13.653
R10612 vp_p.n2571 vp_p.n2570 13.653
R10613 vp_p.n1145 vp_p.n1144 13.653
R10614 vp_p.n9891 vp_p.n9890 13.653
R10615 vp_p.n11328 vp_p.n11327 13.653
R10616 vp_p.n12766 vp_p.n12765 13.653
R10617 vp_p.n26969 vp_p.n26968 13.653
R10618 vp_p.n25544 vp_p.n25543 13.653
R10619 vp_p.n24122 vp_p.n24121 13.653
R10620 vp_p.n22699 vp_p.n22698 13.653
R10621 vp_p.n21275 vp_p.n21274 13.653
R10622 vp_p.n19850 vp_p.n19849 13.653
R10623 vp_p.n18424 vp_p.n18423 13.653
R10624 vp_p.n16997 vp_p.n16996 13.653
R10625 vp_p.n15569 vp_p.n15568 13.653
R10626 vp_p.n13351 vp_p.n13350 13.653
R10627 vp_p.n13349 vp_p.n13348 13.653
R10628 vp_p.n7324 vp_p.n7323 13.653
R10629 vp_p.n5902 vp_p.n5901 13.653
R10630 vp_p.n4479 vp_p.n4478 13.653
R10631 vp_p.n3055 vp_p.n3054 13.653
R10632 vp_p.n1630 vp_p.n1629 13.653
R10633 vp_p.n146 vp_p.n145 13.653
R10634 vp_p.n8885 vp_p.n8884 13.653
R10635 vp_p.n10387 vp_p.n10386 13.653
R10636 vp_p.n11825 vp_p.n11824 13.653
R10637 vp_p.n26029 vp_p.n26028 13.653
R10638 vp_p.n24603 vp_p.n24602 13.653
R10639 vp_p.n23181 vp_p.n23180 13.653
R10640 vp_p.n21758 vp_p.n21757 13.653
R10641 vp_p.n20334 vp_p.n20333 13.653
R10642 vp_p.n18909 vp_p.n18908 13.653
R10643 vp_p.n17483 vp_p.n17482 13.653
R10644 vp_p.n16056 vp_p.n16055 13.653
R10645 vp_p.n14628 vp_p.n14627 13.653
R10646 vp_p.n13344 vp_p.n13343 13.653
R10647 vp_p.n8279 vp_p.n8278 13.653
R10648 vp_p.n6857 vp_p.n6856 13.653
R10649 vp_p.n5434 vp_p.n5433 13.653
R10650 vp_p.n4010 vp_p.n4009 13.653
R10651 vp_p.n2585 vp_p.n2584 13.653
R10652 vp_p.n1159 vp_p.n1158 13.653
R10653 vp_p.n9905 vp_p.n9904 13.653
R10654 vp_p.n11342 vp_p.n11341 13.653
R10655 vp_p.n12780 vp_p.n12779 13.653
R10656 vp_p.n26983 vp_p.n26982 13.653
R10657 vp_p.n25558 vp_p.n25557 13.653
R10658 vp_p.n24136 vp_p.n24135 13.653
R10659 vp_p.n22713 vp_p.n22712 13.653
R10660 vp_p.n21289 vp_p.n21288 13.653
R10661 vp_p.n19864 vp_p.n19863 13.653
R10662 vp_p.n18438 vp_p.n18437 13.653
R10663 vp_p.n17011 vp_p.n17010 13.653
R10664 vp_p.n15583 vp_p.n15582 13.653
R10665 vp_p.n13341 vp_p.n13340 13.653
R10666 vp_p.n13339 vp_p.n13338 13.653
R10667 vp_p.n7319 vp_p.n7318 13.653
R10668 vp_p.n5897 vp_p.n5896 13.653
R10669 vp_p.n4474 vp_p.n4473 13.653
R10670 vp_p.n3050 vp_p.n3049 13.653
R10671 vp_p.n1625 vp_p.n1624 13.653
R10672 vp_p.n141 vp_p.n140 13.653
R10673 vp_p.n8880 vp_p.n8879 13.653
R10674 vp_p.n10382 vp_p.n10381 13.653
R10675 vp_p.n11820 vp_p.n11819 13.653
R10676 vp_p.n26024 vp_p.n26023 13.653
R10677 vp_p.n24598 vp_p.n24597 13.653
R10678 vp_p.n23176 vp_p.n23175 13.653
R10679 vp_p.n21753 vp_p.n21752 13.653
R10680 vp_p.n20329 vp_p.n20328 13.653
R10681 vp_p.n18904 vp_p.n18903 13.653
R10682 vp_p.n17478 vp_p.n17477 13.653
R10683 vp_p.n16051 vp_p.n16050 13.653
R10684 vp_p.n14623 vp_p.n14622 13.653
R10685 vp_p.n13334 vp_p.n13333 13.653
R10686 vp_p.n8293 vp_p.n8292 13.653
R10687 vp_p.n6871 vp_p.n6870 13.653
R10688 vp_p.n5448 vp_p.n5447 13.653
R10689 vp_p.n4024 vp_p.n4023 13.653
R10690 vp_p.n2599 vp_p.n2598 13.653
R10691 vp_p.n1173 vp_p.n1172 13.653
R10692 vp_p.n9919 vp_p.n9918 13.653
R10693 vp_p.n11356 vp_p.n11355 13.653
R10694 vp_p.n12794 vp_p.n12793 13.653
R10695 vp_p.n26997 vp_p.n26996 13.653
R10696 vp_p.n25572 vp_p.n25571 13.653
R10697 vp_p.n24150 vp_p.n24149 13.653
R10698 vp_p.n22727 vp_p.n22726 13.653
R10699 vp_p.n21303 vp_p.n21302 13.653
R10700 vp_p.n19878 vp_p.n19877 13.653
R10701 vp_p.n18452 vp_p.n18451 13.653
R10702 vp_p.n17025 vp_p.n17024 13.653
R10703 vp_p.n15597 vp_p.n15596 13.653
R10704 vp_p.n13331 vp_p.n13330 13.653
R10705 vp_p.n13329 vp_p.n13328 13.653
R10706 vp_p.n7314 vp_p.n7313 13.653
R10707 vp_p.n5892 vp_p.n5891 13.653
R10708 vp_p.n4469 vp_p.n4468 13.653
R10709 vp_p.n3045 vp_p.n3044 13.653
R10710 vp_p.n1620 vp_p.n1619 13.653
R10711 vp_p.n136 vp_p.n135 13.653
R10712 vp_p.n8875 vp_p.n8874 13.653
R10713 vp_p.n10377 vp_p.n10376 13.653
R10714 vp_p.n11815 vp_p.n11814 13.653
R10715 vp_p.n26019 vp_p.n26018 13.653
R10716 vp_p.n24593 vp_p.n24592 13.653
R10717 vp_p.n23171 vp_p.n23170 13.653
R10718 vp_p.n21748 vp_p.n21747 13.653
R10719 vp_p.n20324 vp_p.n20323 13.653
R10720 vp_p.n18899 vp_p.n18898 13.653
R10721 vp_p.n17473 vp_p.n17472 13.653
R10722 vp_p.n16046 vp_p.n16045 13.653
R10723 vp_p.n14618 vp_p.n14617 13.653
R10724 vp_p.n13324 vp_p.n13323 13.653
R10725 vp_p.n8307 vp_p.n8306 13.653
R10726 vp_p.n6885 vp_p.n6884 13.653
R10727 vp_p.n5462 vp_p.n5461 13.653
R10728 vp_p.n4038 vp_p.n4037 13.653
R10729 vp_p.n2613 vp_p.n2612 13.653
R10730 vp_p.n1187 vp_p.n1186 13.653
R10731 vp_p.n9933 vp_p.n9932 13.653
R10732 vp_p.n11370 vp_p.n11369 13.653
R10733 vp_p.n12808 vp_p.n12807 13.653
R10734 vp_p.n27011 vp_p.n27010 13.653
R10735 vp_p.n25586 vp_p.n25585 13.653
R10736 vp_p.n24164 vp_p.n24163 13.653
R10737 vp_p.n22741 vp_p.n22740 13.653
R10738 vp_p.n21317 vp_p.n21316 13.653
R10739 vp_p.n19892 vp_p.n19891 13.653
R10740 vp_p.n18466 vp_p.n18465 13.653
R10741 vp_p.n17039 vp_p.n17038 13.653
R10742 vp_p.n15611 vp_p.n15610 13.653
R10743 vp_p.n13321 vp_p.n13320 13.653
R10744 vp_p.n13319 vp_p.n13318 13.653
R10745 vp_p.n7309 vp_p.n7308 13.653
R10746 vp_p.n5887 vp_p.n5886 13.653
R10747 vp_p.n4464 vp_p.n4463 13.653
R10748 vp_p.n3040 vp_p.n3039 13.653
R10749 vp_p.n1615 vp_p.n1614 13.653
R10750 vp_p.n131 vp_p.n130 13.653
R10751 vp_p.n8870 vp_p.n8869 13.653
R10752 vp_p.n10372 vp_p.n10371 13.653
R10753 vp_p.n11810 vp_p.n11809 13.653
R10754 vp_p.n26014 vp_p.n26013 13.653
R10755 vp_p.n24588 vp_p.n24587 13.653
R10756 vp_p.n23166 vp_p.n23165 13.653
R10757 vp_p.n21743 vp_p.n21742 13.653
R10758 vp_p.n20319 vp_p.n20318 13.653
R10759 vp_p.n18894 vp_p.n18893 13.653
R10760 vp_p.n17468 vp_p.n17467 13.653
R10761 vp_p.n16041 vp_p.n16040 13.653
R10762 vp_p.n14613 vp_p.n14612 13.653
R10763 vp_p.n13314 vp_p.n13313 13.653
R10764 vp_p.n8321 vp_p.n8320 13.653
R10765 vp_p.n6899 vp_p.n6898 13.653
R10766 vp_p.n5476 vp_p.n5475 13.653
R10767 vp_p.n4052 vp_p.n4051 13.653
R10768 vp_p.n2627 vp_p.n2626 13.653
R10769 vp_p.n1201 vp_p.n1200 13.653
R10770 vp_p.n9947 vp_p.n9946 13.653
R10771 vp_p.n11384 vp_p.n11383 13.653
R10772 vp_p.n12822 vp_p.n12821 13.653
R10773 vp_p.n27025 vp_p.n27024 13.653
R10774 vp_p.n25600 vp_p.n25599 13.653
R10775 vp_p.n24178 vp_p.n24177 13.653
R10776 vp_p.n22755 vp_p.n22754 13.653
R10777 vp_p.n21331 vp_p.n21330 13.653
R10778 vp_p.n19906 vp_p.n19905 13.653
R10779 vp_p.n18480 vp_p.n18479 13.653
R10780 vp_p.n17053 vp_p.n17052 13.653
R10781 vp_p.n15625 vp_p.n15624 13.653
R10782 vp_p.n13311 vp_p.n13310 13.653
R10783 vp_p.n13309 vp_p.n13308 13.653
R10784 vp_p.n7304 vp_p.n7303 13.653
R10785 vp_p.n5882 vp_p.n5881 13.653
R10786 vp_p.n4459 vp_p.n4458 13.653
R10787 vp_p.n3035 vp_p.n3034 13.653
R10788 vp_p.n1610 vp_p.n1609 13.653
R10789 vp_p.n126 vp_p.n125 13.653
R10790 vp_p.n8865 vp_p.n8864 13.653
R10791 vp_p.n10367 vp_p.n10366 13.653
R10792 vp_p.n11805 vp_p.n11804 13.653
R10793 vp_p.n26009 vp_p.n26008 13.653
R10794 vp_p.n24583 vp_p.n24582 13.653
R10795 vp_p.n23161 vp_p.n23160 13.653
R10796 vp_p.n21738 vp_p.n21737 13.653
R10797 vp_p.n20314 vp_p.n20313 13.653
R10798 vp_p.n18889 vp_p.n18888 13.653
R10799 vp_p.n17463 vp_p.n17462 13.653
R10800 vp_p.n16036 vp_p.n16035 13.653
R10801 vp_p.n14608 vp_p.n14607 13.653
R10802 vp_p.n13304 vp_p.n13303 13.653
R10803 vp_p.n8335 vp_p.n8334 13.653
R10804 vp_p.n6913 vp_p.n6912 13.653
R10805 vp_p.n5490 vp_p.n5489 13.653
R10806 vp_p.n4066 vp_p.n4065 13.653
R10807 vp_p.n2641 vp_p.n2640 13.653
R10808 vp_p.n1215 vp_p.n1214 13.653
R10809 vp_p.n9961 vp_p.n9960 13.653
R10810 vp_p.n11398 vp_p.n11397 13.653
R10811 vp_p.n12836 vp_p.n12835 13.653
R10812 vp_p.n27039 vp_p.n27038 13.653
R10813 vp_p.n25614 vp_p.n25613 13.653
R10814 vp_p.n24192 vp_p.n24191 13.653
R10815 vp_p.n22769 vp_p.n22768 13.653
R10816 vp_p.n21345 vp_p.n21344 13.653
R10817 vp_p.n19920 vp_p.n19919 13.653
R10818 vp_p.n18494 vp_p.n18493 13.653
R10819 vp_p.n17067 vp_p.n17066 13.653
R10820 vp_p.n15639 vp_p.n15638 13.653
R10821 vp_p.n13301 vp_p.n13300 13.653
R10822 vp_p.n13299 vp_p.n13298 13.653
R10823 vp_p.n7299 vp_p.n7298 13.653
R10824 vp_p.n5877 vp_p.n5876 13.653
R10825 vp_p.n4454 vp_p.n4453 13.653
R10826 vp_p.n3030 vp_p.n3029 13.653
R10827 vp_p.n1605 vp_p.n1604 13.653
R10828 vp_p.n121 vp_p.n120 13.653
R10829 vp_p.n8860 vp_p.n8859 13.653
R10830 vp_p.n10362 vp_p.n10361 13.653
R10831 vp_p.n11800 vp_p.n11799 13.653
R10832 vp_p.n26004 vp_p.n26003 13.653
R10833 vp_p.n24578 vp_p.n24577 13.653
R10834 vp_p.n23156 vp_p.n23155 13.653
R10835 vp_p.n21733 vp_p.n21732 13.653
R10836 vp_p.n20309 vp_p.n20308 13.653
R10837 vp_p.n18884 vp_p.n18883 13.653
R10838 vp_p.n17458 vp_p.n17457 13.653
R10839 vp_p.n16031 vp_p.n16030 13.653
R10840 vp_p.n14603 vp_p.n14602 13.653
R10841 vp_p.n13294 vp_p.n13293 13.653
R10842 vp_p.n8349 vp_p.n8348 13.653
R10843 vp_p.n6927 vp_p.n6926 13.653
R10844 vp_p.n5504 vp_p.n5503 13.653
R10845 vp_p.n4080 vp_p.n4079 13.653
R10846 vp_p.n2655 vp_p.n2654 13.653
R10847 vp_p.n1229 vp_p.n1228 13.653
R10848 vp_p.n9975 vp_p.n9974 13.653
R10849 vp_p.n11412 vp_p.n11411 13.653
R10850 vp_p.n12850 vp_p.n12849 13.653
R10851 vp_p.n27053 vp_p.n27052 13.653
R10852 vp_p.n25628 vp_p.n25627 13.653
R10853 vp_p.n24206 vp_p.n24205 13.653
R10854 vp_p.n22783 vp_p.n22782 13.653
R10855 vp_p.n21359 vp_p.n21358 13.653
R10856 vp_p.n19934 vp_p.n19933 13.653
R10857 vp_p.n18508 vp_p.n18507 13.653
R10858 vp_p.n17081 vp_p.n17080 13.653
R10859 vp_p.n15653 vp_p.n15652 13.653
R10860 vp_p.n13291 vp_p.n13290 13.653
R10861 vp_p.n13289 vp_p.n13288 13.653
R10862 vp_p.n7294 vp_p.n7293 13.653
R10863 vp_p.n5872 vp_p.n5871 13.653
R10864 vp_p.n4449 vp_p.n4448 13.653
R10865 vp_p.n3025 vp_p.n3024 13.653
R10866 vp_p.n1600 vp_p.n1599 13.653
R10867 vp_p.n116 vp_p.n115 13.653
R10868 vp_p.n8855 vp_p.n8854 13.653
R10869 vp_p.n10357 vp_p.n10356 13.653
R10870 vp_p.n11795 vp_p.n11794 13.653
R10871 vp_p.n25999 vp_p.n25998 13.653
R10872 vp_p.n24573 vp_p.n24572 13.653
R10873 vp_p.n23151 vp_p.n23150 13.653
R10874 vp_p.n21728 vp_p.n21727 13.653
R10875 vp_p.n20304 vp_p.n20303 13.653
R10876 vp_p.n18879 vp_p.n18878 13.653
R10877 vp_p.n17453 vp_p.n17452 13.653
R10878 vp_p.n16026 vp_p.n16025 13.653
R10879 vp_p.n14598 vp_p.n14597 13.653
R10880 vp_p.n13284 vp_p.n13283 13.653
R10881 vp_p.n8363 vp_p.n8362 13.653
R10882 vp_p.n6941 vp_p.n6940 13.653
R10883 vp_p.n5518 vp_p.n5517 13.653
R10884 vp_p.n4094 vp_p.n4093 13.653
R10885 vp_p.n2669 vp_p.n2668 13.653
R10886 vp_p.n1243 vp_p.n1242 13.653
R10887 vp_p.n9989 vp_p.n9988 13.653
R10888 vp_p.n11426 vp_p.n11425 13.653
R10889 vp_p.n12864 vp_p.n12863 13.653
R10890 vp_p.n27067 vp_p.n27066 13.653
R10891 vp_p.n25642 vp_p.n25641 13.653
R10892 vp_p.n24220 vp_p.n24219 13.653
R10893 vp_p.n22797 vp_p.n22796 13.653
R10894 vp_p.n21373 vp_p.n21372 13.653
R10895 vp_p.n19948 vp_p.n19947 13.653
R10896 vp_p.n18522 vp_p.n18521 13.653
R10897 vp_p.n17095 vp_p.n17094 13.653
R10898 vp_p.n15667 vp_p.n15666 13.653
R10899 vp_p.n13281 vp_p.n13280 13.653
R10900 vp_p.n13279 vp_p.n13278 13.653
R10901 vp_p.n7289 vp_p.n7288 13.653
R10902 vp_p.n5867 vp_p.n5866 13.653
R10903 vp_p.n4444 vp_p.n4443 13.653
R10904 vp_p.n3020 vp_p.n3019 13.653
R10905 vp_p.n1595 vp_p.n1594 13.653
R10906 vp_p.n111 vp_p.n110 13.653
R10907 vp_p.n8850 vp_p.n8849 13.653
R10908 vp_p.n10352 vp_p.n10351 13.653
R10909 vp_p.n11790 vp_p.n11789 13.653
R10910 vp_p.n25994 vp_p.n25993 13.653
R10911 vp_p.n24568 vp_p.n24567 13.653
R10912 vp_p.n23146 vp_p.n23145 13.653
R10913 vp_p.n21723 vp_p.n21722 13.653
R10914 vp_p.n20299 vp_p.n20298 13.653
R10915 vp_p.n18874 vp_p.n18873 13.653
R10916 vp_p.n17448 vp_p.n17447 13.653
R10917 vp_p.n16021 vp_p.n16020 13.653
R10918 vp_p.n14593 vp_p.n14592 13.653
R10919 vp_p.n13274 vp_p.n13273 13.653
R10920 vp_p.n8377 vp_p.n8376 13.653
R10921 vp_p.n6955 vp_p.n6954 13.653
R10922 vp_p.n5532 vp_p.n5531 13.653
R10923 vp_p.n4108 vp_p.n4107 13.653
R10924 vp_p.n2683 vp_p.n2682 13.653
R10925 vp_p.n1257 vp_p.n1256 13.653
R10926 vp_p.n10003 vp_p.n10002 13.653
R10927 vp_p.n11440 vp_p.n11439 13.653
R10928 vp_p.n12878 vp_p.n12877 13.653
R10929 vp_p.n27081 vp_p.n27080 13.653
R10930 vp_p.n25656 vp_p.n25655 13.653
R10931 vp_p.n24234 vp_p.n24233 13.653
R10932 vp_p.n22811 vp_p.n22810 13.653
R10933 vp_p.n21387 vp_p.n21386 13.653
R10934 vp_p.n19962 vp_p.n19961 13.653
R10935 vp_p.n18536 vp_p.n18535 13.653
R10936 vp_p.n17109 vp_p.n17108 13.653
R10937 vp_p.n15681 vp_p.n15680 13.653
R10938 vp_p.n13271 vp_p.n13270 13.653
R10939 vp_p.n13269 vp_p.n13268 13.653
R10940 vp_p.n7284 vp_p.n7283 13.653
R10941 vp_p.n5862 vp_p.n5861 13.653
R10942 vp_p.n4439 vp_p.n4438 13.653
R10943 vp_p.n3015 vp_p.n3014 13.653
R10944 vp_p.n1590 vp_p.n1589 13.653
R10945 vp_p.n106 vp_p.n105 13.653
R10946 vp_p.n8845 vp_p.n8844 13.653
R10947 vp_p.n10347 vp_p.n10346 13.653
R10948 vp_p.n11785 vp_p.n11784 13.653
R10949 vp_p.n25989 vp_p.n25988 13.653
R10950 vp_p.n24563 vp_p.n24562 13.653
R10951 vp_p.n23141 vp_p.n23140 13.653
R10952 vp_p.n21718 vp_p.n21717 13.653
R10953 vp_p.n20294 vp_p.n20293 13.653
R10954 vp_p.n18869 vp_p.n18868 13.653
R10955 vp_p.n17443 vp_p.n17442 13.653
R10956 vp_p.n16016 vp_p.n16015 13.653
R10957 vp_p.n14588 vp_p.n14587 13.653
R10958 vp_p.n13264 vp_p.n13263 13.653
R10959 vp_p.n8391 vp_p.n8390 13.653
R10960 vp_p.n6969 vp_p.n6968 13.653
R10961 vp_p.n5546 vp_p.n5545 13.653
R10962 vp_p.n4122 vp_p.n4121 13.653
R10963 vp_p.n2697 vp_p.n2696 13.653
R10964 vp_p.n1271 vp_p.n1270 13.653
R10965 vp_p.n10017 vp_p.n10016 13.653
R10966 vp_p.n11454 vp_p.n11453 13.653
R10967 vp_p.n12892 vp_p.n12891 13.653
R10968 vp_p.n27095 vp_p.n27094 13.653
R10969 vp_p.n25670 vp_p.n25669 13.653
R10970 vp_p.n24248 vp_p.n24247 13.653
R10971 vp_p.n22825 vp_p.n22824 13.653
R10972 vp_p.n21401 vp_p.n21400 13.653
R10973 vp_p.n19976 vp_p.n19975 13.653
R10974 vp_p.n18550 vp_p.n18549 13.653
R10975 vp_p.n17123 vp_p.n17122 13.653
R10976 vp_p.n15695 vp_p.n15694 13.653
R10977 vp_p.n13261 vp_p.n13260 13.653
R10978 vp_p.n13259 vp_p.n13258 13.653
R10979 vp_p.n7279 vp_p.n7278 13.653
R10980 vp_p.n5857 vp_p.n5856 13.653
R10981 vp_p.n4434 vp_p.n4433 13.653
R10982 vp_p.n3010 vp_p.n3009 13.653
R10983 vp_p.n1585 vp_p.n1584 13.653
R10984 vp_p.n101 vp_p.n100 13.653
R10985 vp_p.n8840 vp_p.n8839 13.653
R10986 vp_p.n10342 vp_p.n10341 13.653
R10987 vp_p.n11780 vp_p.n11779 13.653
R10988 vp_p.n25984 vp_p.n25983 13.653
R10989 vp_p.n24558 vp_p.n24557 13.653
R10990 vp_p.n23136 vp_p.n23135 13.653
R10991 vp_p.n21713 vp_p.n21712 13.653
R10992 vp_p.n20289 vp_p.n20288 13.653
R10993 vp_p.n18864 vp_p.n18863 13.653
R10994 vp_p.n17438 vp_p.n17437 13.653
R10995 vp_p.n16011 vp_p.n16010 13.653
R10996 vp_p.n14583 vp_p.n14582 13.653
R10997 vp_p.n13254 vp_p.n13253 13.653
R10998 vp_p.n8405 vp_p.n8404 13.653
R10999 vp_p.n6983 vp_p.n6982 13.653
R11000 vp_p.n5560 vp_p.n5559 13.653
R11001 vp_p.n4136 vp_p.n4135 13.653
R11002 vp_p.n2711 vp_p.n2710 13.653
R11003 vp_p.n1285 vp_p.n1284 13.653
R11004 vp_p.n10031 vp_p.n10030 13.653
R11005 vp_p.n11468 vp_p.n11467 13.653
R11006 vp_p.n12906 vp_p.n12905 13.653
R11007 vp_p.n27109 vp_p.n27108 13.653
R11008 vp_p.n25684 vp_p.n25683 13.653
R11009 vp_p.n24262 vp_p.n24261 13.653
R11010 vp_p.n22839 vp_p.n22838 13.653
R11011 vp_p.n21415 vp_p.n21414 13.653
R11012 vp_p.n19990 vp_p.n19989 13.653
R11013 vp_p.n18564 vp_p.n18563 13.653
R11014 vp_p.n17137 vp_p.n17136 13.653
R11015 vp_p.n15709 vp_p.n15708 13.653
R11016 vp_p.n13251 vp_p.n13250 13.653
R11017 vp_p.n13249 vp_p.n13248 13.653
R11018 vp_p.n7274 vp_p.n7273 13.653
R11019 vp_p.n5852 vp_p.n5851 13.653
R11020 vp_p.n4429 vp_p.n4428 13.653
R11021 vp_p.n3005 vp_p.n3004 13.653
R11022 vp_p.n1580 vp_p.n1579 13.653
R11023 vp_p.n96 vp_p.n95 13.653
R11024 vp_p.n8835 vp_p.n8834 13.653
R11025 vp_p.n10337 vp_p.n10336 13.653
R11026 vp_p.n11775 vp_p.n11774 13.653
R11027 vp_p.n25979 vp_p.n25978 13.653
R11028 vp_p.n24553 vp_p.n24552 13.653
R11029 vp_p.n23131 vp_p.n23130 13.653
R11030 vp_p.n21708 vp_p.n21707 13.653
R11031 vp_p.n20284 vp_p.n20283 13.653
R11032 vp_p.n18859 vp_p.n18858 13.653
R11033 vp_p.n17433 vp_p.n17432 13.653
R11034 vp_p.n16006 vp_p.n16005 13.653
R11035 vp_p.n14578 vp_p.n14577 13.653
R11036 vp_p.n13244 vp_p.n13243 13.653
R11037 vp_p.n8419 vp_p.n8418 13.653
R11038 vp_p.n6997 vp_p.n6996 13.653
R11039 vp_p.n5574 vp_p.n5573 13.653
R11040 vp_p.n4150 vp_p.n4149 13.653
R11041 vp_p.n2725 vp_p.n2724 13.653
R11042 vp_p.n1299 vp_p.n1298 13.653
R11043 vp_p.n10045 vp_p.n10044 13.653
R11044 vp_p.n11482 vp_p.n11481 13.653
R11045 vp_p.n12920 vp_p.n12919 13.653
R11046 vp_p.n27123 vp_p.n27122 13.653
R11047 vp_p.n25698 vp_p.n25697 13.653
R11048 vp_p.n24276 vp_p.n24275 13.653
R11049 vp_p.n22853 vp_p.n22852 13.653
R11050 vp_p.n21429 vp_p.n21428 13.653
R11051 vp_p.n20004 vp_p.n20003 13.653
R11052 vp_p.n18578 vp_p.n18577 13.653
R11053 vp_p.n17151 vp_p.n17150 13.653
R11054 vp_p.n15723 vp_p.n15722 13.653
R11055 vp_p.n13241 vp_p.n13240 13.653
R11056 vp_p.n13239 vp_p.n13238 13.653
R11057 vp_p.n7269 vp_p.n7268 13.653
R11058 vp_p.n5847 vp_p.n5846 13.653
R11059 vp_p.n4424 vp_p.n4423 13.653
R11060 vp_p.n3000 vp_p.n2999 13.653
R11061 vp_p.n1575 vp_p.n1574 13.653
R11062 vp_p.n91 vp_p.n90 13.653
R11063 vp_p.n8830 vp_p.n8829 13.653
R11064 vp_p.n10332 vp_p.n10331 13.653
R11065 vp_p.n11770 vp_p.n11769 13.653
R11066 vp_p.n25974 vp_p.n25973 13.653
R11067 vp_p.n24548 vp_p.n24547 13.653
R11068 vp_p.n23126 vp_p.n23125 13.653
R11069 vp_p.n21703 vp_p.n21702 13.653
R11070 vp_p.n20279 vp_p.n20278 13.653
R11071 vp_p.n18854 vp_p.n18853 13.653
R11072 vp_p.n17428 vp_p.n17427 13.653
R11073 vp_p.n16001 vp_p.n16000 13.653
R11074 vp_p.n14573 vp_p.n14572 13.653
R11075 vp_p.n13234 vp_p.n13233 13.653
R11076 vp_p.n8433 vp_p.n8432 13.653
R11077 vp_p.n7011 vp_p.n7010 13.653
R11078 vp_p.n5588 vp_p.n5587 13.653
R11079 vp_p.n4164 vp_p.n4163 13.653
R11080 vp_p.n2739 vp_p.n2738 13.653
R11081 vp_p.n1313 vp_p.n1312 13.653
R11082 vp_p.n10059 vp_p.n10058 13.653
R11083 vp_p.n11496 vp_p.n11495 13.653
R11084 vp_p.n12934 vp_p.n12933 13.653
R11085 vp_p.n27137 vp_p.n27136 13.653
R11086 vp_p.n25712 vp_p.n25711 13.653
R11087 vp_p.n24290 vp_p.n24289 13.653
R11088 vp_p.n22867 vp_p.n22866 13.653
R11089 vp_p.n21443 vp_p.n21442 13.653
R11090 vp_p.n20018 vp_p.n20017 13.653
R11091 vp_p.n18592 vp_p.n18591 13.653
R11092 vp_p.n17165 vp_p.n17164 13.653
R11093 vp_p.n15737 vp_p.n15736 13.653
R11094 vp_p.n13231 vp_p.n13230 13.653
R11095 vp_p.n13229 vp_p.n13228 13.653
R11096 vp_p.n7264 vp_p.n7263 13.653
R11097 vp_p.n5842 vp_p.n5841 13.653
R11098 vp_p.n4419 vp_p.n4418 13.653
R11099 vp_p.n2995 vp_p.n2994 13.653
R11100 vp_p.n1570 vp_p.n1569 13.653
R11101 vp_p.n86 vp_p.n85 13.653
R11102 vp_p.n8825 vp_p.n8824 13.653
R11103 vp_p.n10327 vp_p.n10326 13.653
R11104 vp_p.n11765 vp_p.n11764 13.653
R11105 vp_p.n25969 vp_p.n25968 13.653
R11106 vp_p.n24543 vp_p.n24542 13.653
R11107 vp_p.n23121 vp_p.n23120 13.653
R11108 vp_p.n21698 vp_p.n21697 13.653
R11109 vp_p.n20274 vp_p.n20273 13.653
R11110 vp_p.n18849 vp_p.n18848 13.653
R11111 vp_p.n17423 vp_p.n17422 13.653
R11112 vp_p.n15996 vp_p.n15995 13.653
R11113 vp_p.n14568 vp_p.n14567 13.653
R11114 vp_p.n13224 vp_p.n13223 13.653
R11115 vp_p.n8447 vp_p.n8446 13.653
R11116 vp_p.n7025 vp_p.n7024 13.653
R11117 vp_p.n5602 vp_p.n5601 13.653
R11118 vp_p.n4178 vp_p.n4177 13.653
R11119 vp_p.n2753 vp_p.n2752 13.653
R11120 vp_p.n1327 vp_p.n1326 13.653
R11121 vp_p.n10073 vp_p.n10072 13.653
R11122 vp_p.n11510 vp_p.n11509 13.653
R11123 vp_p.n12948 vp_p.n12947 13.653
R11124 vp_p.n27151 vp_p.n27150 13.653
R11125 vp_p.n25726 vp_p.n25725 13.653
R11126 vp_p.n24304 vp_p.n24303 13.653
R11127 vp_p.n22881 vp_p.n22880 13.653
R11128 vp_p.n21457 vp_p.n21456 13.653
R11129 vp_p.n20032 vp_p.n20031 13.653
R11130 vp_p.n18606 vp_p.n18605 13.653
R11131 vp_p.n17179 vp_p.n17178 13.653
R11132 vp_p.n15751 vp_p.n15750 13.653
R11133 vp_p.n13221 vp_p.n13220 13.653
R11134 vp_p.n13219 vp_p.n13218 13.653
R11135 vp_p.n7259 vp_p.n7258 13.653
R11136 vp_p.n5837 vp_p.n5836 13.653
R11137 vp_p.n4414 vp_p.n4413 13.653
R11138 vp_p.n2990 vp_p.n2989 13.653
R11139 vp_p.n1565 vp_p.n1564 13.653
R11140 vp_p.n81 vp_p.n80 13.653
R11141 vp_p.n8820 vp_p.n8819 13.653
R11142 vp_p.n10322 vp_p.n10321 13.653
R11143 vp_p.n11760 vp_p.n11759 13.653
R11144 vp_p.n25964 vp_p.n25963 13.653
R11145 vp_p.n24538 vp_p.n24537 13.653
R11146 vp_p.n23116 vp_p.n23115 13.653
R11147 vp_p.n21693 vp_p.n21692 13.653
R11148 vp_p.n20269 vp_p.n20268 13.653
R11149 vp_p.n18844 vp_p.n18843 13.653
R11150 vp_p.n17418 vp_p.n17417 13.653
R11151 vp_p.n15991 vp_p.n15990 13.653
R11152 vp_p.n14563 vp_p.n14562 13.653
R11153 vp_p.n13214 vp_p.n13213 13.653
R11154 vp_p.n8461 vp_p.n8460 13.653
R11155 vp_p.n7039 vp_p.n7038 13.653
R11156 vp_p.n5616 vp_p.n5615 13.653
R11157 vp_p.n4192 vp_p.n4191 13.653
R11158 vp_p.n2767 vp_p.n2766 13.653
R11159 vp_p.n1341 vp_p.n1340 13.653
R11160 vp_p.n10087 vp_p.n10086 13.653
R11161 vp_p.n11524 vp_p.n11523 13.653
R11162 vp_p.n12962 vp_p.n12961 13.653
R11163 vp_p.n27165 vp_p.n27164 13.653
R11164 vp_p.n25740 vp_p.n25739 13.653
R11165 vp_p.n24318 vp_p.n24317 13.653
R11166 vp_p.n22895 vp_p.n22894 13.653
R11167 vp_p.n21471 vp_p.n21470 13.653
R11168 vp_p.n20046 vp_p.n20045 13.653
R11169 vp_p.n18620 vp_p.n18619 13.653
R11170 vp_p.n17193 vp_p.n17192 13.653
R11171 vp_p.n15765 vp_p.n15764 13.653
R11172 vp_p.n13211 vp_p.n13210 13.653
R11173 vp_p.n13209 vp_p.n13208 13.653
R11174 vp_p.n7254 vp_p.n7253 13.653
R11175 vp_p.n5832 vp_p.n5831 13.653
R11176 vp_p.n4409 vp_p.n4408 13.653
R11177 vp_p.n2985 vp_p.n2984 13.653
R11178 vp_p.n1560 vp_p.n1559 13.653
R11179 vp_p.n76 vp_p.n75 13.653
R11180 vp_p.n8815 vp_p.n8814 13.653
R11181 vp_p.n10317 vp_p.n10316 13.653
R11182 vp_p.n11755 vp_p.n11754 13.653
R11183 vp_p.n25959 vp_p.n25958 13.653
R11184 vp_p.n24533 vp_p.n24532 13.653
R11185 vp_p.n23111 vp_p.n23110 13.653
R11186 vp_p.n21688 vp_p.n21687 13.653
R11187 vp_p.n20264 vp_p.n20263 13.653
R11188 vp_p.n18839 vp_p.n18838 13.653
R11189 vp_p.n17413 vp_p.n17412 13.653
R11190 vp_p.n15986 vp_p.n15985 13.653
R11191 vp_p.n14558 vp_p.n14557 13.653
R11192 vp_p.n13204 vp_p.n13203 13.653
R11193 vp_p.n8475 vp_p.n8474 13.653
R11194 vp_p.n7053 vp_p.n7052 13.653
R11195 vp_p.n5630 vp_p.n5629 13.653
R11196 vp_p.n4206 vp_p.n4205 13.653
R11197 vp_p.n2781 vp_p.n2780 13.653
R11198 vp_p.n1355 vp_p.n1354 13.653
R11199 vp_p.n10101 vp_p.n10100 13.653
R11200 vp_p.n11538 vp_p.n11537 13.653
R11201 vp_p.n12976 vp_p.n12975 13.653
R11202 vp_p.n27179 vp_p.n27178 13.653
R11203 vp_p.n25754 vp_p.n25753 13.653
R11204 vp_p.n24332 vp_p.n24331 13.653
R11205 vp_p.n22909 vp_p.n22908 13.653
R11206 vp_p.n21485 vp_p.n21484 13.653
R11207 vp_p.n20060 vp_p.n20059 13.653
R11208 vp_p.n18634 vp_p.n18633 13.653
R11209 vp_p.n17207 vp_p.n17206 13.653
R11210 vp_p.n15779 vp_p.n15778 13.653
R11211 vp_p.n13201 vp_p.n13200 13.653
R11212 vp_p.n13199 vp_p.n13198 13.653
R11213 vp_p.n7249 vp_p.n7248 13.653
R11214 vp_p.n5827 vp_p.n5826 13.653
R11215 vp_p.n4404 vp_p.n4403 13.653
R11216 vp_p.n2980 vp_p.n2979 13.653
R11217 vp_p.n1555 vp_p.n1554 13.653
R11218 vp_p.n71 vp_p.n70 13.653
R11219 vp_p.n8810 vp_p.n8809 13.653
R11220 vp_p.n10312 vp_p.n10311 13.653
R11221 vp_p.n11750 vp_p.n11749 13.653
R11222 vp_p.n25954 vp_p.n25953 13.653
R11223 vp_p.n24528 vp_p.n24527 13.653
R11224 vp_p.n23106 vp_p.n23105 13.653
R11225 vp_p.n21683 vp_p.n21682 13.653
R11226 vp_p.n20259 vp_p.n20258 13.653
R11227 vp_p.n18834 vp_p.n18833 13.653
R11228 vp_p.n17408 vp_p.n17407 13.653
R11229 vp_p.n15981 vp_p.n15980 13.653
R11230 vp_p.n14553 vp_p.n14552 13.653
R11231 vp_p.n13194 vp_p.n13193 13.653
R11232 vp_p.n8489 vp_p.n8488 13.653
R11233 vp_p.n7067 vp_p.n7066 13.653
R11234 vp_p.n5644 vp_p.n5643 13.653
R11235 vp_p.n4220 vp_p.n4219 13.653
R11236 vp_p.n2795 vp_p.n2794 13.653
R11237 vp_p.n1369 vp_p.n1368 13.653
R11238 vp_p.n10115 vp_p.n10114 13.653
R11239 vp_p.n11552 vp_p.n11551 13.653
R11240 vp_p.n12990 vp_p.n12989 13.653
R11241 vp_p.n27193 vp_p.n27192 13.653
R11242 vp_p.n25768 vp_p.n25767 13.653
R11243 vp_p.n24346 vp_p.n24345 13.653
R11244 vp_p.n22923 vp_p.n22922 13.653
R11245 vp_p.n21499 vp_p.n21498 13.653
R11246 vp_p.n20074 vp_p.n20073 13.653
R11247 vp_p.n18648 vp_p.n18647 13.653
R11248 vp_p.n17221 vp_p.n17220 13.653
R11249 vp_p.n15793 vp_p.n15792 13.653
R11250 vp_p.n13191 vp_p.n13190 13.653
R11251 vp_p.n13189 vp_p.n13188 13.653
R11252 vp_p.n7244 vp_p.n7243 13.653
R11253 vp_p.n5822 vp_p.n5821 13.653
R11254 vp_p.n4399 vp_p.n4398 13.653
R11255 vp_p.n2975 vp_p.n2974 13.653
R11256 vp_p.n1550 vp_p.n1549 13.653
R11257 vp_p.n66 vp_p.n65 13.653
R11258 vp_p.n8805 vp_p.n8804 13.653
R11259 vp_p.n10307 vp_p.n10306 13.653
R11260 vp_p.n11745 vp_p.n11744 13.653
R11261 vp_p.n25949 vp_p.n25948 13.653
R11262 vp_p.n24523 vp_p.n24522 13.653
R11263 vp_p.n23101 vp_p.n23100 13.653
R11264 vp_p.n21678 vp_p.n21677 13.653
R11265 vp_p.n20254 vp_p.n20253 13.653
R11266 vp_p.n18829 vp_p.n18828 13.653
R11267 vp_p.n17403 vp_p.n17402 13.653
R11268 vp_p.n15976 vp_p.n15975 13.653
R11269 vp_p.n14548 vp_p.n14547 13.653
R11270 vp_p.n13184 vp_p.n13183 13.653
R11271 vp_p.n8503 vp_p.n8502 13.653
R11272 vp_p.n7081 vp_p.n7080 13.653
R11273 vp_p.n5658 vp_p.n5657 13.653
R11274 vp_p.n4234 vp_p.n4233 13.653
R11275 vp_p.n2809 vp_p.n2808 13.653
R11276 vp_p.n1383 vp_p.n1382 13.653
R11277 vp_p.n10129 vp_p.n10128 13.653
R11278 vp_p.n11566 vp_p.n11565 13.653
R11279 vp_p.n13004 vp_p.n13003 13.653
R11280 vp_p.n27207 vp_p.n27206 13.653
R11281 vp_p.n25782 vp_p.n25781 13.653
R11282 vp_p.n24360 vp_p.n24359 13.653
R11283 vp_p.n22937 vp_p.n22936 13.653
R11284 vp_p.n21513 vp_p.n21512 13.653
R11285 vp_p.n20088 vp_p.n20087 13.653
R11286 vp_p.n18662 vp_p.n18661 13.653
R11287 vp_p.n17235 vp_p.n17234 13.653
R11288 vp_p.n15807 vp_p.n15806 13.653
R11289 vp_p.n13181 vp_p.n13180 13.653
R11290 vp_p.n13179 vp_p.n13178 13.653
R11291 vp_p.n13186 vp_p.n13185 13.653
R11292 vp_p.n13196 vp_p.n13195 13.653
R11293 vp_p.n13206 vp_p.n13205 13.653
R11294 vp_p.n13216 vp_p.n13215 13.653
R11295 vp_p.n13226 vp_p.n13225 13.653
R11296 vp_p.n13236 vp_p.n13235 13.653
R11297 vp_p.n13246 vp_p.n13245 13.653
R11298 vp_p.n13256 vp_p.n13255 13.653
R11299 vp_p.n13266 vp_p.n13265 13.653
R11300 vp_p.n13276 vp_p.n13275 13.653
R11301 vp_p.n13286 vp_p.n13285 13.653
R11302 vp_p.n13296 vp_p.n13295 13.653
R11303 vp_p.n13306 vp_p.n13305 13.653
R11304 vp_p.n13316 vp_p.n13315 13.653
R11305 vp_p.n13326 vp_p.n13325 13.653
R11306 vp_p.n13336 vp_p.n13335 13.653
R11307 vp_p.n13346 vp_p.n13345 13.653
R11308 vp_p.n13356 vp_p.n13355 13.653
R11309 vp_p.n13366 vp_p.n13365 13.653
R11310 vp_p.n13376 vp_p.n13375 13.653
R11311 vp_p.n13386 vp_p.n13385 13.653
R11312 vp_p.n13396 vp_p.n13395 13.653
R11313 vp_p.n13406 vp_p.n13405 13.653
R11314 vp_p.n13416 vp_p.n13415 13.653
R11315 vp_p.n13426 vp_p.n13425 13.653
R11316 vp_p.n13436 vp_p.n13435 13.653
R11317 vp_p.n13446 vp_p.n13445 13.653
R11318 vp_p.n13456 vp_p.n13455 13.653
R11319 vp_p.n13466 vp_p.n13465 13.653
R11320 vp_p.n13476 vp_p.n13475 13.653
R11321 vp_p.n13486 vp_p.n13485 13.653
R11322 vp_p.n13496 vp_p.n13495 13.653
R11323 vp_p.n13506 vp_p.n13505 13.653
R11324 vp_p.n13516 vp_p.n13515 13.653
R11325 vp_p.n13526 vp_p.n13525 13.653
R11326 vp_p.n13536 vp_p.n13535 13.653
R11327 vp_p.n13546 vp_p.n13545 13.653
R11328 vp_p.n13556 vp_p.n13555 13.653
R11329 vp_p.n13566 vp_p.n13565 13.653
R11330 vp_p.n13576 vp_p.n13575 13.653
R11331 vp_p.n13586 vp_p.n13585 13.653
R11332 vp_p.n13596 vp_p.n13595 13.653
R11333 vp_p.n13606 vp_p.n13605 13.653
R11334 vp_p.n13616 vp_p.n13615 13.653
R11335 vp_p.n13626 vp_p.n13625 13.653
R11336 vp_p.n13636 vp_p.n13635 13.653
R11337 vp_p.n13646 vp_p.n13645 13.653
R11338 vp_p.n13656 vp_p.n13655 13.653
R11339 vp_p.n13666 vp_p.n13665 13.653
R11340 vp_p.n13676 vp_p.n13675 13.653
R11341 vp_p.n13686 vp_p.n13685 13.653
R11342 vp_p.n13696 vp_p.n13695 13.653
R11343 vp_p.n13706 vp_p.n13705 13.653
R11344 vp_p.n13716 vp_p.n13715 13.653
R11345 vp_p.n13726 vp_p.n13725 13.653
R11346 vp_p.n13736 vp_p.n13735 13.653
R11347 vp_p.n13746 vp_p.n13745 13.653
R11348 vp_p.n13756 vp_p.n13755 13.653
R11349 vp_p.n13766 vp_p.n13765 13.653
R11350 vp_p.n13776 vp_p.n13775 13.653
R11351 vp_p.n13786 vp_p.n13785 13.653
R11352 vp_p.n13796 vp_p.n13795 13.653
R11353 vp_p.n13806 vp_p.n13805 13.653
R11354 vp_p.n13816 vp_p.n13815 13.653
R11355 vp_p.n13826 vp_p.n13825 13.653
R11356 vp_p.n25944 vp_p.n25943 13.653
R11357 vp_p.n24518 vp_p.n24517 13.653
R11358 vp_p.n23096 vp_p.n23095 13.653
R11359 vp_p.n21673 vp_p.n21672 13.653
R11360 vp_p.n20249 vp_p.n20248 13.653
R11361 vp_p.n18824 vp_p.n18823 13.653
R11362 vp_p.n17398 vp_p.n17397 13.653
R11363 vp_p.n15971 vp_p.n15970 13.653
R11364 vp_p.n14543 vp_p.n14542 13.653
R11365 vp_p.n14382 vp_p.n14381 13.653
R11366 vp_p.n14380 vp_p.n14379 13.653
R11367 vp_p.n11740 vp_p.n11739 13.653
R11368 vp_p.n11742 vp_p.n11741 13.653
R11369 vp_p.n13002 vp_p.n13001 13.653
R11370 vp_p.n11747 vp_p.n11746 13.653
R11371 vp_p.n12988 vp_p.n12987 13.653
R11372 vp_p.n11752 vp_p.n11751 13.653
R11373 vp_p.n12974 vp_p.n12973 13.653
R11374 vp_p.n11757 vp_p.n11756 13.653
R11375 vp_p.n12960 vp_p.n12959 13.653
R11376 vp_p.n11762 vp_p.n11761 13.653
R11377 vp_p.n12946 vp_p.n12945 13.653
R11378 vp_p.n11767 vp_p.n11766 13.653
R11379 vp_p.n12932 vp_p.n12931 13.653
R11380 vp_p.n11772 vp_p.n11771 13.653
R11381 vp_p.n12918 vp_p.n12917 13.653
R11382 vp_p.n11777 vp_p.n11776 13.653
R11383 vp_p.n12904 vp_p.n12903 13.653
R11384 vp_p.n11782 vp_p.n11781 13.653
R11385 vp_p.n12890 vp_p.n12889 13.653
R11386 vp_p.n11787 vp_p.n11786 13.653
R11387 vp_p.n12876 vp_p.n12875 13.653
R11388 vp_p.n11792 vp_p.n11791 13.653
R11389 vp_p.n12862 vp_p.n12861 13.653
R11390 vp_p.n11797 vp_p.n11796 13.653
R11391 vp_p.n12848 vp_p.n12847 13.653
R11392 vp_p.n11802 vp_p.n11801 13.653
R11393 vp_p.n12834 vp_p.n12833 13.653
R11394 vp_p.n11807 vp_p.n11806 13.653
R11395 vp_p.n12820 vp_p.n12819 13.653
R11396 vp_p.n11812 vp_p.n11811 13.653
R11397 vp_p.n12806 vp_p.n12805 13.653
R11398 vp_p.n11817 vp_p.n11816 13.653
R11399 vp_p.n12792 vp_p.n12791 13.653
R11400 vp_p.n11822 vp_p.n11821 13.653
R11401 vp_p.n12778 vp_p.n12777 13.653
R11402 vp_p.n11827 vp_p.n11826 13.653
R11403 vp_p.n12764 vp_p.n12763 13.653
R11404 vp_p.n11832 vp_p.n11831 13.653
R11405 vp_p.n12750 vp_p.n12749 13.653
R11406 vp_p.n11837 vp_p.n11836 13.653
R11407 vp_p.n12736 vp_p.n12735 13.653
R11408 vp_p.n11842 vp_p.n11841 13.653
R11409 vp_p.n12722 vp_p.n12721 13.653
R11410 vp_p.n11847 vp_p.n11846 13.653
R11411 vp_p.n12708 vp_p.n12707 13.653
R11412 vp_p.n11852 vp_p.n11851 13.653
R11413 vp_p.n12694 vp_p.n12693 13.653
R11414 vp_p.n11857 vp_p.n11856 13.653
R11415 vp_p.n12680 vp_p.n12679 13.653
R11416 vp_p.n11862 vp_p.n11861 13.653
R11417 vp_p.n12666 vp_p.n12665 13.653
R11418 vp_p.n11867 vp_p.n11866 13.653
R11419 vp_p.n12652 vp_p.n12651 13.653
R11420 vp_p.n11872 vp_p.n11871 13.653
R11421 vp_p.n12638 vp_p.n12637 13.653
R11422 vp_p.n11877 vp_p.n11876 13.653
R11423 vp_p.n12624 vp_p.n12623 13.653
R11424 vp_p.n11882 vp_p.n11881 13.653
R11425 vp_p.n12610 vp_p.n12609 13.653
R11426 vp_p.n11887 vp_p.n11886 13.653
R11427 vp_p.n12596 vp_p.n12595 13.653
R11428 vp_p.n11892 vp_p.n11891 13.653
R11429 vp_p.n12582 vp_p.n12581 13.653
R11430 vp_p.n11897 vp_p.n11896 13.653
R11431 vp_p.n12568 vp_p.n12567 13.653
R11432 vp_p.n11902 vp_p.n11901 13.653
R11433 vp_p.n12554 vp_p.n12553 13.653
R11434 vp_p.n11907 vp_p.n11906 13.653
R11435 vp_p.n12540 vp_p.n12539 13.653
R11436 vp_p.n11912 vp_p.n11911 13.653
R11437 vp_p.n12526 vp_p.n12525 13.653
R11438 vp_p.n11917 vp_p.n11916 13.653
R11439 vp_p.n12512 vp_p.n12511 13.653
R11440 vp_p.n11922 vp_p.n11921 13.653
R11441 vp_p.n12498 vp_p.n12497 13.653
R11442 vp_p.n11927 vp_p.n11926 13.653
R11443 vp_p.n12484 vp_p.n12483 13.653
R11444 vp_p.n11932 vp_p.n11931 13.653
R11445 vp_p.n12470 vp_p.n12469 13.653
R11446 vp_p.n11937 vp_p.n11936 13.653
R11447 vp_p.n12456 vp_p.n12455 13.653
R11448 vp_p.n11942 vp_p.n11941 13.653
R11449 vp_p.n12442 vp_p.n12441 13.653
R11450 vp_p.n11947 vp_p.n11946 13.653
R11451 vp_p.n12428 vp_p.n12427 13.653
R11452 vp_p.n11952 vp_p.n11951 13.653
R11453 vp_p.n12414 vp_p.n12413 13.653
R11454 vp_p.n11957 vp_p.n11956 13.653
R11455 vp_p.n12400 vp_p.n12399 13.653
R11456 vp_p.n11962 vp_p.n11961 13.653
R11457 vp_p.n12386 vp_p.n12385 13.653
R11458 vp_p.n11967 vp_p.n11966 13.653
R11459 vp_p.n12372 vp_p.n12371 13.653
R11460 vp_p.n11972 vp_p.n11971 13.653
R11461 vp_p.n12358 vp_p.n12357 13.653
R11462 vp_p.n11977 vp_p.n11976 13.653
R11463 vp_p.n12344 vp_p.n12343 13.653
R11464 vp_p.n11982 vp_p.n11981 13.653
R11465 vp_p.n12330 vp_p.n12329 13.653
R11466 vp_p.n11987 vp_p.n11986 13.653
R11467 vp_p.n12316 vp_p.n12315 13.653
R11468 vp_p.n11992 vp_p.n11991 13.653
R11469 vp_p.n12302 vp_p.n12301 13.653
R11470 vp_p.n11997 vp_p.n11996 13.653
R11471 vp_p.n12288 vp_p.n12287 13.653
R11472 vp_p.n12002 vp_p.n12001 13.653
R11473 vp_p.n12274 vp_p.n12273 13.653
R11474 vp_p.n12007 vp_p.n12006 13.653
R11475 vp_p.n12260 vp_p.n12259 13.653
R11476 vp_p.n12012 vp_p.n12011 13.653
R11477 vp_p.n12246 vp_p.n12245 13.653
R11478 vp_p.n12017 vp_p.n12016 13.653
R11479 vp_p.n12232 vp_p.n12231 13.653
R11480 vp_p.n12022 vp_p.n12021 13.653
R11481 vp_p.n12218 vp_p.n12217 13.653
R11482 vp_p.n12027 vp_p.n12026 13.653
R11483 vp_p.n12204 vp_p.n12203 13.653
R11484 vp_p.n12032 vp_p.n12031 13.653
R11485 vp_p.n12190 vp_p.n12189 13.653
R11486 vp_p.n12037 vp_p.n12036 13.653
R11487 vp_p.n12176 vp_p.n12175 13.653
R11488 vp_p.n12042 vp_p.n12041 13.653
R11489 vp_p.n12162 vp_p.n12161 13.653
R11490 vp_p.n12047 vp_p.n12046 13.653
R11491 vp_p.n12148 vp_p.n12147 13.653
R11492 vp_p.n12052 vp_p.n12051 13.653
R11493 vp_p.n12134 vp_p.n12133 13.653
R11494 vp_p.n12057 vp_p.n12056 13.653
R11495 vp_p.n12120 vp_p.n12119 13.653
R11496 vp_p.n12062 vp_p.n12061 13.653
R11497 vp_p.n12106 vp_p.n12105 13.653
R11498 vp_p.n12067 vp_p.n12066 13.653
R11499 vp_p.n12092 vp_p.n12091 13.653
R11500 vp_p.n8517 vp_p.n8516 13.653
R11501 vp_p.n7095 vp_p.n7094 13.653
R11502 vp_p.n5672 vp_p.n5671 13.653
R11503 vp_p.n4248 vp_p.n4247 13.653
R11504 vp_p.n2823 vp_p.n2822 13.653
R11505 vp_p.n1397 vp_p.n1396 13.653
R11506 vp_p.n10143 vp_p.n10142 13.653
R11507 vp_p.n11580 vp_p.n11579 13.653
R11508 vp_p.n13016 vp_p.n13015 13.653
R11509 vp_p.n13018 vp_p.n13017 13.653
R11510 vp_p.n13174 vp_p.n13173 13.653
R11511 vp_p.n13176 vp_p.n13175 13.653
R11512 vp_p.n27221 vp_p.n27220 13.653
R11513 vp_p.n25796 vp_p.n25795 13.653
R11514 vp_p.n24374 vp_p.n24373 13.653
R11515 vp_p.n22951 vp_p.n22950 13.653
R11516 vp_p.n21527 vp_p.n21526 13.653
R11517 vp_p.n20102 vp_p.n20101 13.653
R11518 vp_p.n18676 vp_p.n18675 13.653
R11519 vp_p.n17249 vp_p.n17248 13.653
R11520 vp_p.n14540 vp_p.n14539 13.653
R11521 vp_p.n14538 vp_p.n14537 13.653
R11522 vp_p.n14545 vp_p.n14544 13.653
R11523 vp_p.n15805 vp_p.n15804 13.653
R11524 vp_p.n14550 vp_p.n14549 13.653
R11525 vp_p.n15791 vp_p.n15790 13.653
R11526 vp_p.n14555 vp_p.n14554 13.653
R11527 vp_p.n15777 vp_p.n15776 13.653
R11528 vp_p.n14560 vp_p.n14559 13.653
R11529 vp_p.n15763 vp_p.n15762 13.653
R11530 vp_p.n14565 vp_p.n14564 13.653
R11531 vp_p.n15749 vp_p.n15748 13.653
R11532 vp_p.n14570 vp_p.n14569 13.653
R11533 vp_p.n15735 vp_p.n15734 13.653
R11534 vp_p.n14575 vp_p.n14574 13.653
R11535 vp_p.n15721 vp_p.n15720 13.653
R11536 vp_p.n14580 vp_p.n14579 13.653
R11537 vp_p.n15707 vp_p.n15706 13.653
R11538 vp_p.n14585 vp_p.n14584 13.653
R11539 vp_p.n15693 vp_p.n15692 13.653
R11540 vp_p.n14590 vp_p.n14589 13.653
R11541 vp_p.n15679 vp_p.n15678 13.653
R11542 vp_p.n14595 vp_p.n14594 13.653
R11543 vp_p.n15665 vp_p.n15664 13.653
R11544 vp_p.n14600 vp_p.n14599 13.653
R11545 vp_p.n15651 vp_p.n15650 13.653
R11546 vp_p.n14605 vp_p.n14604 13.653
R11547 vp_p.n15637 vp_p.n15636 13.653
R11548 vp_p.n14610 vp_p.n14609 13.653
R11549 vp_p.n15623 vp_p.n15622 13.653
R11550 vp_p.n14615 vp_p.n14614 13.653
R11551 vp_p.n15609 vp_p.n15608 13.653
R11552 vp_p.n14620 vp_p.n14619 13.653
R11553 vp_p.n15595 vp_p.n15594 13.653
R11554 vp_p.n14625 vp_p.n14624 13.653
R11555 vp_p.n15581 vp_p.n15580 13.653
R11556 vp_p.n14630 vp_p.n14629 13.653
R11557 vp_p.n15567 vp_p.n15566 13.653
R11558 vp_p.n14635 vp_p.n14634 13.653
R11559 vp_p.n15553 vp_p.n15552 13.653
R11560 vp_p.n14640 vp_p.n14639 13.653
R11561 vp_p.n15539 vp_p.n15538 13.653
R11562 vp_p.n14645 vp_p.n14644 13.653
R11563 vp_p.n15525 vp_p.n15524 13.653
R11564 vp_p.n14650 vp_p.n14649 13.653
R11565 vp_p.n15511 vp_p.n15510 13.653
R11566 vp_p.n14655 vp_p.n14654 13.653
R11567 vp_p.n15497 vp_p.n15496 13.653
R11568 vp_p.n14660 vp_p.n14659 13.653
R11569 vp_p.n15483 vp_p.n15482 13.653
R11570 vp_p.n14665 vp_p.n14664 13.653
R11571 vp_p.n15469 vp_p.n15468 13.653
R11572 vp_p.n14670 vp_p.n14669 13.653
R11573 vp_p.n15455 vp_p.n15454 13.653
R11574 vp_p.n14675 vp_p.n14674 13.653
R11575 vp_p.n15441 vp_p.n15440 13.653
R11576 vp_p.n14680 vp_p.n14679 13.653
R11577 vp_p.n15427 vp_p.n15426 13.653
R11578 vp_p.n14685 vp_p.n14684 13.653
R11579 vp_p.n15413 vp_p.n15412 13.653
R11580 vp_p.n14690 vp_p.n14689 13.653
R11581 vp_p.n15399 vp_p.n15398 13.653
R11582 vp_p.n14695 vp_p.n14694 13.653
R11583 vp_p.n15385 vp_p.n15384 13.653
R11584 vp_p.n14700 vp_p.n14699 13.653
R11585 vp_p.n15371 vp_p.n15370 13.653
R11586 vp_p.n14705 vp_p.n14704 13.653
R11587 vp_p.n15357 vp_p.n15356 13.653
R11588 vp_p.n14710 vp_p.n14709 13.653
R11589 vp_p.n15343 vp_p.n15342 13.653
R11590 vp_p.n14715 vp_p.n14714 13.653
R11591 vp_p.n15329 vp_p.n15328 13.653
R11592 vp_p.n14720 vp_p.n14719 13.653
R11593 vp_p.n15315 vp_p.n15314 13.653
R11594 vp_p.n14725 vp_p.n14724 13.653
R11595 vp_p.n15301 vp_p.n15300 13.653
R11596 vp_p.n14730 vp_p.n14729 13.653
R11597 vp_p.n15287 vp_p.n15286 13.653
R11598 vp_p.n14735 vp_p.n14734 13.653
R11599 vp_p.n15273 vp_p.n15272 13.653
R11600 vp_p.n14740 vp_p.n14739 13.653
R11601 vp_p.n15259 vp_p.n15258 13.653
R11602 vp_p.n14745 vp_p.n14744 13.653
R11603 vp_p.n15245 vp_p.n15244 13.653
R11604 vp_p.n14750 vp_p.n14749 13.653
R11605 vp_p.n15231 vp_p.n15230 13.653
R11606 vp_p.n14755 vp_p.n14754 13.653
R11607 vp_p.n15217 vp_p.n15216 13.653
R11608 vp_p.n14760 vp_p.n14759 13.653
R11609 vp_p.n15203 vp_p.n15202 13.653
R11610 vp_p.n14765 vp_p.n14764 13.653
R11611 vp_p.n15189 vp_p.n15188 13.653
R11612 vp_p.n14770 vp_p.n14769 13.653
R11613 vp_p.n15175 vp_p.n15174 13.653
R11614 vp_p.n14775 vp_p.n14774 13.653
R11615 vp_p.n15161 vp_p.n15160 13.653
R11616 vp_p.n14780 vp_p.n14779 13.653
R11617 vp_p.n15147 vp_p.n15146 13.653
R11618 vp_p.n14785 vp_p.n14784 13.653
R11619 vp_p.n15133 vp_p.n15132 13.653
R11620 vp_p.n14790 vp_p.n14789 13.653
R11621 vp_p.n15119 vp_p.n15118 13.653
R11622 vp_p.n14795 vp_p.n14794 13.653
R11623 vp_p.n15105 vp_p.n15104 13.653
R11624 vp_p.n14800 vp_p.n14799 13.653
R11625 vp_p.n15091 vp_p.n15090 13.653
R11626 vp_p.n14805 vp_p.n14804 13.653
R11627 vp_p.n15077 vp_p.n15076 13.653
R11628 vp_p.n14810 vp_p.n14809 13.653
R11629 vp_p.n15063 vp_p.n15062 13.653
R11630 vp_p.n14815 vp_p.n14814 13.653
R11631 vp_p.n15049 vp_p.n15048 13.653
R11632 vp_p.n14820 vp_p.n14819 13.653
R11633 vp_p.n15035 vp_p.n15034 13.653
R11634 vp_p.n14825 vp_p.n14824 13.653
R11635 vp_p.n15021 vp_p.n15020 13.653
R11636 vp_p.n14830 vp_p.n14829 13.653
R11637 vp_p.n15007 vp_p.n15006 13.653
R11638 vp_p.n14835 vp_p.n14834 13.653
R11639 vp_p.n14993 vp_p.n14992 13.653
R11640 vp_p.n14840 vp_p.n14839 13.653
R11641 vp_p.n14979 vp_p.n14978 13.653
R11642 vp_p.n14845 vp_p.n14844 13.653
R11643 vp_p.n14965 vp_p.n14964 13.653
R11644 vp_p.n14850 vp_p.n14849 13.653
R11645 vp_p.n14951 vp_p.n14950 13.653
R11646 vp_p.n14855 vp_p.n14854 13.653
R11647 vp_p.n14937 vp_p.n14936 13.653
R11648 vp_p.n14860 vp_p.n14859 13.653
R11649 vp_p.n14923 vp_p.n14922 13.653
R11650 vp_p.n14865 vp_p.n14864 13.653
R11651 vp_p.n14909 vp_p.n14908 13.653
R11652 vp_p.n14870 vp_p.n14869 13.653
R11653 vp_p.n14895 vp_p.n14894 13.653
R11654 vp_p.n25939 vp_p.n25938 13.653
R11655 vp_p.n24513 vp_p.n24512 13.653
R11656 vp_p.n23091 vp_p.n23090 13.653
R11657 vp_p.n21668 vp_p.n21667 13.653
R11658 vp_p.n20244 vp_p.n20243 13.653
R11659 vp_p.n18819 vp_p.n18818 13.653
R11660 vp_p.n17393 vp_p.n17392 13.653
R11661 vp_p.n15966 vp_p.n15965 13.653
R11662 vp_p.n15825 vp_p.n15824 13.653
R11663 vp_p.n15823 vp_p.n15822 13.653
R11664 vp_p.n13169 vp_p.n13168 13.653
R11665 vp_p.n13171 vp_p.n13170 13.653
R11666 vp_p.n11735 vp_p.n11734 13.653
R11667 vp_p.n11737 vp_p.n11736 13.653
R11668 vp_p.n10297 vp_p.n10296 13.653
R11669 vp_p.n10299 vp_p.n10298 13.653
R11670 vp_p.n11578 vp_p.n11577 13.653
R11671 vp_p.n10304 vp_p.n10303 13.653
R11672 vp_p.n11564 vp_p.n11563 13.653
R11673 vp_p.n10309 vp_p.n10308 13.653
R11674 vp_p.n11550 vp_p.n11549 13.653
R11675 vp_p.n10314 vp_p.n10313 13.653
R11676 vp_p.n11536 vp_p.n11535 13.653
R11677 vp_p.n10319 vp_p.n10318 13.653
R11678 vp_p.n11522 vp_p.n11521 13.653
R11679 vp_p.n10324 vp_p.n10323 13.653
R11680 vp_p.n11508 vp_p.n11507 13.653
R11681 vp_p.n10329 vp_p.n10328 13.653
R11682 vp_p.n11494 vp_p.n11493 13.653
R11683 vp_p.n10334 vp_p.n10333 13.653
R11684 vp_p.n11480 vp_p.n11479 13.653
R11685 vp_p.n10339 vp_p.n10338 13.653
R11686 vp_p.n11466 vp_p.n11465 13.653
R11687 vp_p.n10344 vp_p.n10343 13.653
R11688 vp_p.n11452 vp_p.n11451 13.653
R11689 vp_p.n10349 vp_p.n10348 13.653
R11690 vp_p.n11438 vp_p.n11437 13.653
R11691 vp_p.n10354 vp_p.n10353 13.653
R11692 vp_p.n11424 vp_p.n11423 13.653
R11693 vp_p.n10359 vp_p.n10358 13.653
R11694 vp_p.n11410 vp_p.n11409 13.653
R11695 vp_p.n10364 vp_p.n10363 13.653
R11696 vp_p.n11396 vp_p.n11395 13.653
R11697 vp_p.n10369 vp_p.n10368 13.653
R11698 vp_p.n11382 vp_p.n11381 13.653
R11699 vp_p.n10374 vp_p.n10373 13.653
R11700 vp_p.n11368 vp_p.n11367 13.653
R11701 vp_p.n10379 vp_p.n10378 13.653
R11702 vp_p.n11354 vp_p.n11353 13.653
R11703 vp_p.n10384 vp_p.n10383 13.653
R11704 vp_p.n11340 vp_p.n11339 13.653
R11705 vp_p.n10389 vp_p.n10388 13.653
R11706 vp_p.n11326 vp_p.n11325 13.653
R11707 vp_p.n10394 vp_p.n10393 13.653
R11708 vp_p.n11312 vp_p.n11311 13.653
R11709 vp_p.n10399 vp_p.n10398 13.653
R11710 vp_p.n11298 vp_p.n11297 13.653
R11711 vp_p.n10404 vp_p.n10403 13.653
R11712 vp_p.n11284 vp_p.n11283 13.653
R11713 vp_p.n10409 vp_p.n10408 13.653
R11714 vp_p.n11270 vp_p.n11269 13.653
R11715 vp_p.n10414 vp_p.n10413 13.653
R11716 vp_p.n11256 vp_p.n11255 13.653
R11717 vp_p.n10419 vp_p.n10418 13.653
R11718 vp_p.n11242 vp_p.n11241 13.653
R11719 vp_p.n10424 vp_p.n10423 13.653
R11720 vp_p.n11228 vp_p.n11227 13.653
R11721 vp_p.n10429 vp_p.n10428 13.653
R11722 vp_p.n11214 vp_p.n11213 13.653
R11723 vp_p.n10434 vp_p.n10433 13.653
R11724 vp_p.n11200 vp_p.n11199 13.653
R11725 vp_p.n10439 vp_p.n10438 13.653
R11726 vp_p.n11186 vp_p.n11185 13.653
R11727 vp_p.n10444 vp_p.n10443 13.653
R11728 vp_p.n11172 vp_p.n11171 13.653
R11729 vp_p.n10449 vp_p.n10448 13.653
R11730 vp_p.n11158 vp_p.n11157 13.653
R11731 vp_p.n10454 vp_p.n10453 13.653
R11732 vp_p.n11144 vp_p.n11143 13.653
R11733 vp_p.n10459 vp_p.n10458 13.653
R11734 vp_p.n11130 vp_p.n11129 13.653
R11735 vp_p.n10464 vp_p.n10463 13.653
R11736 vp_p.n11116 vp_p.n11115 13.653
R11737 vp_p.n10469 vp_p.n10468 13.653
R11738 vp_p.n11102 vp_p.n11101 13.653
R11739 vp_p.n10474 vp_p.n10473 13.653
R11740 vp_p.n11088 vp_p.n11087 13.653
R11741 vp_p.n10479 vp_p.n10478 13.653
R11742 vp_p.n11074 vp_p.n11073 13.653
R11743 vp_p.n10484 vp_p.n10483 13.653
R11744 vp_p.n11060 vp_p.n11059 13.653
R11745 vp_p.n10489 vp_p.n10488 13.653
R11746 vp_p.n11046 vp_p.n11045 13.653
R11747 vp_p.n10494 vp_p.n10493 13.653
R11748 vp_p.n11032 vp_p.n11031 13.653
R11749 vp_p.n10499 vp_p.n10498 13.653
R11750 vp_p.n11018 vp_p.n11017 13.653
R11751 vp_p.n10504 vp_p.n10503 13.653
R11752 vp_p.n11004 vp_p.n11003 13.653
R11753 vp_p.n10509 vp_p.n10508 13.653
R11754 vp_p.n10990 vp_p.n10989 13.653
R11755 vp_p.n10514 vp_p.n10513 13.653
R11756 vp_p.n10976 vp_p.n10975 13.653
R11757 vp_p.n10519 vp_p.n10518 13.653
R11758 vp_p.n10962 vp_p.n10961 13.653
R11759 vp_p.n10524 vp_p.n10523 13.653
R11760 vp_p.n10948 vp_p.n10947 13.653
R11761 vp_p.n10529 vp_p.n10528 13.653
R11762 vp_p.n10934 vp_p.n10933 13.653
R11763 vp_p.n10534 vp_p.n10533 13.653
R11764 vp_p.n10920 vp_p.n10919 13.653
R11765 vp_p.n10539 vp_p.n10538 13.653
R11766 vp_p.n10906 vp_p.n10905 13.653
R11767 vp_p.n10544 vp_p.n10543 13.653
R11768 vp_p.n10892 vp_p.n10891 13.653
R11769 vp_p.n10549 vp_p.n10548 13.653
R11770 vp_p.n10878 vp_p.n10877 13.653
R11771 vp_p.n10554 vp_p.n10553 13.653
R11772 vp_p.n10864 vp_p.n10863 13.653
R11773 vp_p.n10559 vp_p.n10558 13.653
R11774 vp_p.n10850 vp_p.n10849 13.653
R11775 vp_p.n10564 vp_p.n10563 13.653
R11776 vp_p.n10836 vp_p.n10835 13.653
R11777 vp_p.n10569 vp_p.n10568 13.653
R11778 vp_p.n10822 vp_p.n10821 13.653
R11779 vp_p.n10574 vp_p.n10573 13.653
R11780 vp_p.n10808 vp_p.n10807 13.653
R11781 vp_p.n10579 vp_p.n10578 13.653
R11782 vp_p.n10794 vp_p.n10793 13.653
R11783 vp_p.n10584 vp_p.n10583 13.653
R11784 vp_p.n10780 vp_p.n10779 13.653
R11785 vp_p.n10589 vp_p.n10588 13.653
R11786 vp_p.n10766 vp_p.n10765 13.653
R11787 vp_p.n10594 vp_p.n10593 13.653
R11788 vp_p.n10752 vp_p.n10751 13.653
R11789 vp_p.n10599 vp_p.n10598 13.653
R11790 vp_p.n10738 vp_p.n10737 13.653
R11791 vp_p.n10604 vp_p.n10603 13.653
R11792 vp_p.n10724 vp_p.n10723 13.653
R11793 vp_p.n10609 vp_p.n10608 13.653
R11794 vp_p.n10710 vp_p.n10709 13.653
R11795 vp_p.n10614 vp_p.n10613 13.653
R11796 vp_p.n10696 vp_p.n10695 13.653
R11797 vp_p.n10619 vp_p.n10618 13.653
R11798 vp_p.n10682 vp_p.n10681 13.653
R11799 vp_p.n10624 vp_p.n10623 13.653
R11800 vp_p.n10668 vp_p.n10667 13.653
R11801 vp_p.n10629 vp_p.n10628 13.653
R11802 vp_p.n10654 vp_p.n10653 13.653
R11803 vp_p.n8531 vp_p.n8530 13.653
R11804 vp_p.n7109 vp_p.n7108 13.653
R11805 vp_p.n5686 vp_p.n5685 13.653
R11806 vp_p.n4262 vp_p.n4261 13.653
R11807 vp_p.n2837 vp_p.n2836 13.653
R11808 vp_p.n1411 vp_p.n1410 13.653
R11809 vp_p.n10157 vp_p.n10156 13.653
R11810 vp_p.n11592 vp_p.n11591 13.653
R11811 vp_p.n11594 vp_p.n11593 13.653
R11812 vp_p.n11730 vp_p.n11729 13.653
R11813 vp_p.n11732 vp_p.n11731 13.653
R11814 vp_p.n13164 vp_p.n13163 13.653
R11815 vp_p.n13166 vp_p.n13165 13.653
R11816 vp_p.n14533 vp_p.n14532 13.653
R11817 vp_p.n14535 vp_p.n14534 13.653
R11818 vp_p.n27235 vp_p.n27234 13.653
R11819 vp_p.n25810 vp_p.n25809 13.653
R11820 vp_p.n24388 vp_p.n24387 13.653
R11821 vp_p.n22965 vp_p.n22964 13.653
R11822 vp_p.n21541 vp_p.n21540 13.653
R11823 vp_p.n20116 vp_p.n20115 13.653
R11824 vp_p.n18690 vp_p.n18689 13.653
R11825 vp_p.n15963 vp_p.n15962 13.653
R11826 vp_p.n15961 vp_p.n15960 13.653
R11827 vp_p.n15968 vp_p.n15967 13.653
R11828 vp_p.n17247 vp_p.n17246 13.653
R11829 vp_p.n15973 vp_p.n15972 13.653
R11830 vp_p.n17233 vp_p.n17232 13.653
R11831 vp_p.n15978 vp_p.n15977 13.653
R11832 vp_p.n17219 vp_p.n17218 13.653
R11833 vp_p.n15983 vp_p.n15982 13.653
R11834 vp_p.n17205 vp_p.n17204 13.653
R11835 vp_p.n15988 vp_p.n15987 13.653
R11836 vp_p.n17191 vp_p.n17190 13.653
R11837 vp_p.n15993 vp_p.n15992 13.653
R11838 vp_p.n17177 vp_p.n17176 13.653
R11839 vp_p.n15998 vp_p.n15997 13.653
R11840 vp_p.n17163 vp_p.n17162 13.653
R11841 vp_p.n16003 vp_p.n16002 13.653
R11842 vp_p.n17149 vp_p.n17148 13.653
R11843 vp_p.n16008 vp_p.n16007 13.653
R11844 vp_p.n17135 vp_p.n17134 13.653
R11845 vp_p.n16013 vp_p.n16012 13.653
R11846 vp_p.n17121 vp_p.n17120 13.653
R11847 vp_p.n16018 vp_p.n16017 13.653
R11848 vp_p.n17107 vp_p.n17106 13.653
R11849 vp_p.n16023 vp_p.n16022 13.653
R11850 vp_p.n17093 vp_p.n17092 13.653
R11851 vp_p.n16028 vp_p.n16027 13.653
R11852 vp_p.n17079 vp_p.n17078 13.653
R11853 vp_p.n16033 vp_p.n16032 13.653
R11854 vp_p.n17065 vp_p.n17064 13.653
R11855 vp_p.n16038 vp_p.n16037 13.653
R11856 vp_p.n17051 vp_p.n17050 13.653
R11857 vp_p.n16043 vp_p.n16042 13.653
R11858 vp_p.n17037 vp_p.n17036 13.653
R11859 vp_p.n16048 vp_p.n16047 13.653
R11860 vp_p.n17023 vp_p.n17022 13.653
R11861 vp_p.n16053 vp_p.n16052 13.653
R11862 vp_p.n17009 vp_p.n17008 13.653
R11863 vp_p.n16058 vp_p.n16057 13.653
R11864 vp_p.n16995 vp_p.n16994 13.653
R11865 vp_p.n16063 vp_p.n16062 13.653
R11866 vp_p.n16981 vp_p.n16980 13.653
R11867 vp_p.n16068 vp_p.n16067 13.653
R11868 vp_p.n16967 vp_p.n16966 13.653
R11869 vp_p.n16073 vp_p.n16072 13.653
R11870 vp_p.n16953 vp_p.n16952 13.653
R11871 vp_p.n16078 vp_p.n16077 13.653
R11872 vp_p.n16939 vp_p.n16938 13.653
R11873 vp_p.n16083 vp_p.n16082 13.653
R11874 vp_p.n16925 vp_p.n16924 13.653
R11875 vp_p.n16088 vp_p.n16087 13.653
R11876 vp_p.n16911 vp_p.n16910 13.653
R11877 vp_p.n16093 vp_p.n16092 13.653
R11878 vp_p.n16897 vp_p.n16896 13.653
R11879 vp_p.n16098 vp_p.n16097 13.653
R11880 vp_p.n16883 vp_p.n16882 13.653
R11881 vp_p.n16103 vp_p.n16102 13.653
R11882 vp_p.n16869 vp_p.n16868 13.653
R11883 vp_p.n16108 vp_p.n16107 13.653
R11884 vp_p.n16855 vp_p.n16854 13.653
R11885 vp_p.n16113 vp_p.n16112 13.653
R11886 vp_p.n16841 vp_p.n16840 13.653
R11887 vp_p.n16118 vp_p.n16117 13.653
R11888 vp_p.n16827 vp_p.n16826 13.653
R11889 vp_p.n16123 vp_p.n16122 13.653
R11890 vp_p.n16813 vp_p.n16812 13.653
R11891 vp_p.n16128 vp_p.n16127 13.653
R11892 vp_p.n16799 vp_p.n16798 13.653
R11893 vp_p.n16133 vp_p.n16132 13.653
R11894 vp_p.n16785 vp_p.n16784 13.653
R11895 vp_p.n16138 vp_p.n16137 13.653
R11896 vp_p.n16771 vp_p.n16770 13.653
R11897 vp_p.n16143 vp_p.n16142 13.653
R11898 vp_p.n16757 vp_p.n16756 13.653
R11899 vp_p.n16148 vp_p.n16147 13.653
R11900 vp_p.n16743 vp_p.n16742 13.653
R11901 vp_p.n16153 vp_p.n16152 13.653
R11902 vp_p.n16729 vp_p.n16728 13.653
R11903 vp_p.n16158 vp_p.n16157 13.653
R11904 vp_p.n16715 vp_p.n16714 13.653
R11905 vp_p.n16163 vp_p.n16162 13.653
R11906 vp_p.n16701 vp_p.n16700 13.653
R11907 vp_p.n16168 vp_p.n16167 13.653
R11908 vp_p.n16687 vp_p.n16686 13.653
R11909 vp_p.n16173 vp_p.n16172 13.653
R11910 vp_p.n16673 vp_p.n16672 13.653
R11911 vp_p.n16178 vp_p.n16177 13.653
R11912 vp_p.n16659 vp_p.n16658 13.653
R11913 vp_p.n16183 vp_p.n16182 13.653
R11914 vp_p.n16645 vp_p.n16644 13.653
R11915 vp_p.n16188 vp_p.n16187 13.653
R11916 vp_p.n16631 vp_p.n16630 13.653
R11917 vp_p.n16193 vp_p.n16192 13.653
R11918 vp_p.n16617 vp_p.n16616 13.653
R11919 vp_p.n16198 vp_p.n16197 13.653
R11920 vp_p.n16603 vp_p.n16602 13.653
R11921 vp_p.n16203 vp_p.n16202 13.653
R11922 vp_p.n16589 vp_p.n16588 13.653
R11923 vp_p.n16208 vp_p.n16207 13.653
R11924 vp_p.n16575 vp_p.n16574 13.653
R11925 vp_p.n16213 vp_p.n16212 13.653
R11926 vp_p.n16561 vp_p.n16560 13.653
R11927 vp_p.n16218 vp_p.n16217 13.653
R11928 vp_p.n16547 vp_p.n16546 13.653
R11929 vp_p.n16223 vp_p.n16222 13.653
R11930 vp_p.n16533 vp_p.n16532 13.653
R11931 vp_p.n16228 vp_p.n16227 13.653
R11932 vp_p.n16519 vp_p.n16518 13.653
R11933 vp_p.n16233 vp_p.n16232 13.653
R11934 vp_p.n16505 vp_p.n16504 13.653
R11935 vp_p.n16238 vp_p.n16237 13.653
R11936 vp_p.n16491 vp_p.n16490 13.653
R11937 vp_p.n16243 vp_p.n16242 13.653
R11938 vp_p.n16477 vp_p.n16476 13.653
R11939 vp_p.n16248 vp_p.n16247 13.653
R11940 vp_p.n16463 vp_p.n16462 13.653
R11941 vp_p.n16253 vp_p.n16252 13.653
R11942 vp_p.n16449 vp_p.n16448 13.653
R11943 vp_p.n16258 vp_p.n16257 13.653
R11944 vp_p.n16435 vp_p.n16434 13.653
R11945 vp_p.n16263 vp_p.n16262 13.653
R11946 vp_p.n16421 vp_p.n16420 13.653
R11947 vp_p.n16268 vp_p.n16267 13.653
R11948 vp_p.n16407 vp_p.n16406 13.653
R11949 vp_p.n16273 vp_p.n16272 13.653
R11950 vp_p.n16393 vp_p.n16392 13.653
R11951 vp_p.n16278 vp_p.n16277 13.653
R11952 vp_p.n16379 vp_p.n16378 13.653
R11953 vp_p.n16283 vp_p.n16282 13.653
R11954 vp_p.n16365 vp_p.n16364 13.653
R11955 vp_p.n16288 vp_p.n16287 13.653
R11956 vp_p.n16351 vp_p.n16350 13.653
R11957 vp_p.n16293 vp_p.n16292 13.653
R11958 vp_p.n16337 vp_p.n16336 13.653
R11959 vp_p.n16298 vp_p.n16297 13.653
R11960 vp_p.n16323 vp_p.n16322 13.653
R11961 vp_p.n25934 vp_p.n25933 13.653
R11962 vp_p.n24508 vp_p.n24507 13.653
R11963 vp_p.n23086 vp_p.n23085 13.653
R11964 vp_p.n21663 vp_p.n21662 13.653
R11965 vp_p.n20239 vp_p.n20238 13.653
R11966 vp_p.n18814 vp_p.n18813 13.653
R11967 vp_p.n17388 vp_p.n17387 13.653
R11968 vp_p.n17267 vp_p.n17266 13.653
R11969 vp_p.n17265 vp_p.n17264 13.653
R11970 vp_p.n14528 vp_p.n14527 13.653
R11971 vp_p.n14530 vp_p.n14529 13.653
R11972 vp_p.n13159 vp_p.n13158 13.653
R11973 vp_p.n13161 vp_p.n13160 13.653
R11974 vp_p.n11725 vp_p.n11724 13.653
R11975 vp_p.n11727 vp_p.n11726 13.653
R11976 vp_p.n10292 vp_p.n10291 13.653
R11977 vp_p.n10294 vp_p.n10293 13.653
R11978 vp_p.n8790 vp_p.n8789 13.653
R11979 vp_p.n8792 vp_p.n8791 13.653
R11980 vp_p.n10155 vp_p.n10154 13.653
R11981 vp_p.n8797 vp_p.n8796 13.653
R11982 vp_p.n10141 vp_p.n10140 13.653
R11983 vp_p.n8802 vp_p.n8801 13.653
R11984 vp_p.n10127 vp_p.n10126 13.653
R11985 vp_p.n8807 vp_p.n8806 13.653
R11986 vp_p.n10113 vp_p.n10112 13.653
R11987 vp_p.n8812 vp_p.n8811 13.653
R11988 vp_p.n10099 vp_p.n10098 13.653
R11989 vp_p.n8817 vp_p.n8816 13.653
R11990 vp_p.n10085 vp_p.n10084 13.653
R11991 vp_p.n8822 vp_p.n8821 13.653
R11992 vp_p.n10071 vp_p.n10070 13.653
R11993 vp_p.n8827 vp_p.n8826 13.653
R11994 vp_p.n10057 vp_p.n10056 13.653
R11995 vp_p.n8832 vp_p.n8831 13.653
R11996 vp_p.n10043 vp_p.n10042 13.653
R11997 vp_p.n8837 vp_p.n8836 13.653
R11998 vp_p.n10029 vp_p.n10028 13.653
R11999 vp_p.n8842 vp_p.n8841 13.653
R12000 vp_p.n10015 vp_p.n10014 13.653
R12001 vp_p.n8847 vp_p.n8846 13.653
R12002 vp_p.n10001 vp_p.n10000 13.653
R12003 vp_p.n8852 vp_p.n8851 13.653
R12004 vp_p.n9987 vp_p.n9986 13.653
R12005 vp_p.n8857 vp_p.n8856 13.653
R12006 vp_p.n9973 vp_p.n9972 13.653
R12007 vp_p.n8862 vp_p.n8861 13.653
R12008 vp_p.n9959 vp_p.n9958 13.653
R12009 vp_p.n8867 vp_p.n8866 13.653
R12010 vp_p.n9945 vp_p.n9944 13.653
R12011 vp_p.n8872 vp_p.n8871 13.653
R12012 vp_p.n9931 vp_p.n9930 13.653
R12013 vp_p.n8877 vp_p.n8876 13.653
R12014 vp_p.n9917 vp_p.n9916 13.653
R12015 vp_p.n8882 vp_p.n8881 13.653
R12016 vp_p.n9903 vp_p.n9902 13.653
R12017 vp_p.n8887 vp_p.n8886 13.653
R12018 vp_p.n9889 vp_p.n9888 13.653
R12019 vp_p.n8892 vp_p.n8891 13.653
R12020 vp_p.n9875 vp_p.n9874 13.653
R12021 vp_p.n8897 vp_p.n8896 13.653
R12022 vp_p.n9861 vp_p.n9860 13.653
R12023 vp_p.n8902 vp_p.n8901 13.653
R12024 vp_p.n9847 vp_p.n9846 13.653
R12025 vp_p.n8907 vp_p.n8906 13.653
R12026 vp_p.n9833 vp_p.n9832 13.653
R12027 vp_p.n8912 vp_p.n8911 13.653
R12028 vp_p.n9819 vp_p.n9818 13.653
R12029 vp_p.n8917 vp_p.n8916 13.653
R12030 vp_p.n9805 vp_p.n9804 13.653
R12031 vp_p.n8922 vp_p.n8921 13.653
R12032 vp_p.n9791 vp_p.n9790 13.653
R12033 vp_p.n8927 vp_p.n8926 13.653
R12034 vp_p.n9777 vp_p.n9776 13.653
R12035 vp_p.n8932 vp_p.n8931 13.653
R12036 vp_p.n9763 vp_p.n9762 13.653
R12037 vp_p.n8937 vp_p.n8936 13.653
R12038 vp_p.n9749 vp_p.n9748 13.653
R12039 vp_p.n8942 vp_p.n8941 13.653
R12040 vp_p.n9735 vp_p.n9734 13.653
R12041 vp_p.n8947 vp_p.n8946 13.653
R12042 vp_p.n9721 vp_p.n9720 13.653
R12043 vp_p.n8952 vp_p.n8951 13.653
R12044 vp_p.n9707 vp_p.n9706 13.653
R12045 vp_p.n8957 vp_p.n8956 13.653
R12046 vp_p.n9693 vp_p.n9692 13.653
R12047 vp_p.n8962 vp_p.n8961 13.653
R12048 vp_p.n9679 vp_p.n9678 13.653
R12049 vp_p.n8967 vp_p.n8966 13.653
R12050 vp_p.n9665 vp_p.n9664 13.653
R12051 vp_p.n8972 vp_p.n8971 13.653
R12052 vp_p.n9651 vp_p.n9650 13.653
R12053 vp_p.n8977 vp_p.n8976 13.653
R12054 vp_p.n9637 vp_p.n9636 13.653
R12055 vp_p.n8982 vp_p.n8981 13.653
R12056 vp_p.n9623 vp_p.n9622 13.653
R12057 vp_p.n8987 vp_p.n8986 13.653
R12058 vp_p.n9609 vp_p.n9608 13.653
R12059 vp_p.n8992 vp_p.n8991 13.653
R12060 vp_p.n9595 vp_p.n9594 13.653
R12061 vp_p.n8997 vp_p.n8996 13.653
R12062 vp_p.n9581 vp_p.n9580 13.653
R12063 vp_p.n9002 vp_p.n9001 13.653
R12064 vp_p.n9567 vp_p.n9566 13.653
R12065 vp_p.n9007 vp_p.n9006 13.653
R12066 vp_p.n9553 vp_p.n9552 13.653
R12067 vp_p.n9012 vp_p.n9011 13.653
R12068 vp_p.n9539 vp_p.n9538 13.653
R12069 vp_p.n9017 vp_p.n9016 13.653
R12070 vp_p.n9525 vp_p.n9524 13.653
R12071 vp_p.n9022 vp_p.n9021 13.653
R12072 vp_p.n9511 vp_p.n9510 13.653
R12073 vp_p.n9027 vp_p.n9026 13.653
R12074 vp_p.n9497 vp_p.n9496 13.653
R12075 vp_p.n9032 vp_p.n9031 13.653
R12076 vp_p.n9483 vp_p.n9482 13.653
R12077 vp_p.n9037 vp_p.n9036 13.653
R12078 vp_p.n9469 vp_p.n9468 13.653
R12079 vp_p.n9042 vp_p.n9041 13.653
R12080 vp_p.n9455 vp_p.n9454 13.653
R12081 vp_p.n9047 vp_p.n9046 13.653
R12082 vp_p.n9441 vp_p.n9440 13.653
R12083 vp_p.n9052 vp_p.n9051 13.653
R12084 vp_p.n9427 vp_p.n9426 13.653
R12085 vp_p.n9057 vp_p.n9056 13.653
R12086 vp_p.n9413 vp_p.n9412 13.653
R12087 vp_p.n9062 vp_p.n9061 13.653
R12088 vp_p.n9399 vp_p.n9398 13.653
R12089 vp_p.n9067 vp_p.n9066 13.653
R12090 vp_p.n9385 vp_p.n9384 13.653
R12091 vp_p.n9072 vp_p.n9071 13.653
R12092 vp_p.n9371 vp_p.n9370 13.653
R12093 vp_p.n9077 vp_p.n9076 13.653
R12094 vp_p.n9357 vp_p.n9356 13.653
R12095 vp_p.n9082 vp_p.n9081 13.653
R12096 vp_p.n9343 vp_p.n9342 13.653
R12097 vp_p.n9087 vp_p.n9086 13.653
R12098 vp_p.n9329 vp_p.n9328 13.653
R12099 vp_p.n9092 vp_p.n9091 13.653
R12100 vp_p.n9315 vp_p.n9314 13.653
R12101 vp_p.n9097 vp_p.n9096 13.653
R12102 vp_p.n9301 vp_p.n9300 13.653
R12103 vp_p.n9102 vp_p.n9101 13.653
R12104 vp_p.n9287 vp_p.n9286 13.653
R12105 vp_p.n9107 vp_p.n9106 13.653
R12106 vp_p.n9273 vp_p.n9272 13.653
R12107 vp_p.n9112 vp_p.n9111 13.653
R12108 vp_p.n9259 vp_p.n9258 13.653
R12109 vp_p.n9117 vp_p.n9116 13.653
R12110 vp_p.n9245 vp_p.n9244 13.653
R12111 vp_p.n9122 vp_p.n9121 13.653
R12112 vp_p.n9231 vp_p.n9230 13.653
R12113 vp_p.n9127 vp_p.n9126 13.653
R12114 vp_p.n9217 vp_p.n9216 13.653
R12115 vp_p.n8545 vp_p.n8544 13.653
R12116 vp_p.n7123 vp_p.n7122 13.653
R12117 vp_p.n5700 vp_p.n5699 13.653
R12118 vp_p.n4276 vp_p.n4275 13.653
R12119 vp_p.n2851 vp_p.n2850 13.653
R12120 vp_p.n1425 vp_p.n1424 13.653
R12121 vp_p.n10169 vp_p.n10168 13.653
R12122 vp_p.n10171 vp_p.n10170 13.653
R12123 vp_p.n10287 vp_p.n10286 13.653
R12124 vp_p.n10289 vp_p.n10288 13.653
R12125 vp_p.n11720 vp_p.n11719 13.653
R12126 vp_p.n11722 vp_p.n11721 13.653
R12127 vp_p.n13154 vp_p.n13153 13.653
R12128 vp_p.n13156 vp_p.n13155 13.653
R12129 vp_p.n14523 vp_p.n14522 13.653
R12130 vp_p.n14525 vp_p.n14524 13.653
R12131 vp_p.n15956 vp_p.n15955 13.653
R12132 vp_p.n15958 vp_p.n15957 13.653
R12133 vp_p.n27249 vp_p.n27248 13.653
R12134 vp_p.n25824 vp_p.n25823 13.653
R12135 vp_p.n24402 vp_p.n24401 13.653
R12136 vp_p.n22979 vp_p.n22978 13.653
R12137 vp_p.n21555 vp_p.n21554 13.653
R12138 vp_p.n20130 vp_p.n20129 13.653
R12139 vp_p.n17385 vp_p.n17384 13.653
R12140 vp_p.n17383 vp_p.n17382 13.653
R12141 vp_p.n17390 vp_p.n17389 13.653
R12142 vp_p.n18688 vp_p.n18687 13.653
R12143 vp_p.n17395 vp_p.n17394 13.653
R12144 vp_p.n18674 vp_p.n18673 13.653
R12145 vp_p.n17400 vp_p.n17399 13.653
R12146 vp_p.n18660 vp_p.n18659 13.653
R12147 vp_p.n17405 vp_p.n17404 13.653
R12148 vp_p.n18646 vp_p.n18645 13.653
R12149 vp_p.n17410 vp_p.n17409 13.653
R12150 vp_p.n18632 vp_p.n18631 13.653
R12151 vp_p.n17415 vp_p.n17414 13.653
R12152 vp_p.n18618 vp_p.n18617 13.653
R12153 vp_p.n17420 vp_p.n17419 13.653
R12154 vp_p.n18604 vp_p.n18603 13.653
R12155 vp_p.n17425 vp_p.n17424 13.653
R12156 vp_p.n18590 vp_p.n18589 13.653
R12157 vp_p.n17430 vp_p.n17429 13.653
R12158 vp_p.n18576 vp_p.n18575 13.653
R12159 vp_p.n17435 vp_p.n17434 13.653
R12160 vp_p.n18562 vp_p.n18561 13.653
R12161 vp_p.n17440 vp_p.n17439 13.653
R12162 vp_p.n18548 vp_p.n18547 13.653
R12163 vp_p.n17445 vp_p.n17444 13.653
R12164 vp_p.n18534 vp_p.n18533 13.653
R12165 vp_p.n17450 vp_p.n17449 13.653
R12166 vp_p.n18520 vp_p.n18519 13.653
R12167 vp_p.n17455 vp_p.n17454 13.653
R12168 vp_p.n18506 vp_p.n18505 13.653
R12169 vp_p.n17460 vp_p.n17459 13.653
R12170 vp_p.n18492 vp_p.n18491 13.653
R12171 vp_p.n17465 vp_p.n17464 13.653
R12172 vp_p.n18478 vp_p.n18477 13.653
R12173 vp_p.n17470 vp_p.n17469 13.653
R12174 vp_p.n18464 vp_p.n18463 13.653
R12175 vp_p.n17475 vp_p.n17474 13.653
R12176 vp_p.n18450 vp_p.n18449 13.653
R12177 vp_p.n17480 vp_p.n17479 13.653
R12178 vp_p.n18436 vp_p.n18435 13.653
R12179 vp_p.n17485 vp_p.n17484 13.653
R12180 vp_p.n18422 vp_p.n18421 13.653
R12181 vp_p.n17490 vp_p.n17489 13.653
R12182 vp_p.n18408 vp_p.n18407 13.653
R12183 vp_p.n17495 vp_p.n17494 13.653
R12184 vp_p.n18394 vp_p.n18393 13.653
R12185 vp_p.n17500 vp_p.n17499 13.653
R12186 vp_p.n18380 vp_p.n18379 13.653
R12187 vp_p.n17505 vp_p.n17504 13.653
R12188 vp_p.n18366 vp_p.n18365 13.653
R12189 vp_p.n17510 vp_p.n17509 13.653
R12190 vp_p.n18352 vp_p.n18351 13.653
R12191 vp_p.n17515 vp_p.n17514 13.653
R12192 vp_p.n18338 vp_p.n18337 13.653
R12193 vp_p.n17520 vp_p.n17519 13.653
R12194 vp_p.n18324 vp_p.n18323 13.653
R12195 vp_p.n17525 vp_p.n17524 13.653
R12196 vp_p.n18310 vp_p.n18309 13.653
R12197 vp_p.n17530 vp_p.n17529 13.653
R12198 vp_p.n18296 vp_p.n18295 13.653
R12199 vp_p.n17535 vp_p.n17534 13.653
R12200 vp_p.n18282 vp_p.n18281 13.653
R12201 vp_p.n17540 vp_p.n17539 13.653
R12202 vp_p.n18268 vp_p.n18267 13.653
R12203 vp_p.n17545 vp_p.n17544 13.653
R12204 vp_p.n18254 vp_p.n18253 13.653
R12205 vp_p.n17550 vp_p.n17549 13.653
R12206 vp_p.n18240 vp_p.n18239 13.653
R12207 vp_p.n17555 vp_p.n17554 13.653
R12208 vp_p.n18226 vp_p.n18225 13.653
R12209 vp_p.n17560 vp_p.n17559 13.653
R12210 vp_p.n18212 vp_p.n18211 13.653
R12211 vp_p.n17565 vp_p.n17564 13.653
R12212 vp_p.n18198 vp_p.n18197 13.653
R12213 vp_p.n17570 vp_p.n17569 13.653
R12214 vp_p.n18184 vp_p.n18183 13.653
R12215 vp_p.n17575 vp_p.n17574 13.653
R12216 vp_p.n18170 vp_p.n18169 13.653
R12217 vp_p.n17580 vp_p.n17579 13.653
R12218 vp_p.n18156 vp_p.n18155 13.653
R12219 vp_p.n17585 vp_p.n17584 13.653
R12220 vp_p.n18142 vp_p.n18141 13.653
R12221 vp_p.n17590 vp_p.n17589 13.653
R12222 vp_p.n18128 vp_p.n18127 13.653
R12223 vp_p.n17595 vp_p.n17594 13.653
R12224 vp_p.n18114 vp_p.n18113 13.653
R12225 vp_p.n17600 vp_p.n17599 13.653
R12226 vp_p.n18100 vp_p.n18099 13.653
R12227 vp_p.n17605 vp_p.n17604 13.653
R12228 vp_p.n18086 vp_p.n18085 13.653
R12229 vp_p.n17610 vp_p.n17609 13.653
R12230 vp_p.n18072 vp_p.n18071 13.653
R12231 vp_p.n17615 vp_p.n17614 13.653
R12232 vp_p.n18058 vp_p.n18057 13.653
R12233 vp_p.n17620 vp_p.n17619 13.653
R12234 vp_p.n18044 vp_p.n18043 13.653
R12235 vp_p.n17625 vp_p.n17624 13.653
R12236 vp_p.n18030 vp_p.n18029 13.653
R12237 vp_p.n17630 vp_p.n17629 13.653
R12238 vp_p.n18016 vp_p.n18015 13.653
R12239 vp_p.n17635 vp_p.n17634 13.653
R12240 vp_p.n18002 vp_p.n18001 13.653
R12241 vp_p.n17640 vp_p.n17639 13.653
R12242 vp_p.n17988 vp_p.n17987 13.653
R12243 vp_p.n17645 vp_p.n17644 13.653
R12244 vp_p.n17974 vp_p.n17973 13.653
R12245 vp_p.n17650 vp_p.n17649 13.653
R12246 vp_p.n17960 vp_p.n17959 13.653
R12247 vp_p.n17655 vp_p.n17654 13.653
R12248 vp_p.n17946 vp_p.n17945 13.653
R12249 vp_p.n17660 vp_p.n17659 13.653
R12250 vp_p.n17932 vp_p.n17931 13.653
R12251 vp_p.n17665 vp_p.n17664 13.653
R12252 vp_p.n17918 vp_p.n17917 13.653
R12253 vp_p.n17670 vp_p.n17669 13.653
R12254 vp_p.n17904 vp_p.n17903 13.653
R12255 vp_p.n17675 vp_p.n17674 13.653
R12256 vp_p.n17890 vp_p.n17889 13.653
R12257 vp_p.n17680 vp_p.n17679 13.653
R12258 vp_p.n17876 vp_p.n17875 13.653
R12259 vp_p.n17685 vp_p.n17684 13.653
R12260 vp_p.n17862 vp_p.n17861 13.653
R12261 vp_p.n17690 vp_p.n17689 13.653
R12262 vp_p.n17848 vp_p.n17847 13.653
R12263 vp_p.n17695 vp_p.n17694 13.653
R12264 vp_p.n17834 vp_p.n17833 13.653
R12265 vp_p.n17700 vp_p.n17699 13.653
R12266 vp_p.n17820 vp_p.n17819 13.653
R12267 vp_p.n17705 vp_p.n17704 13.653
R12268 vp_p.n17806 vp_p.n17805 13.653
R12269 vp_p.n17710 vp_p.n17709 13.653
R12270 vp_p.n17792 vp_p.n17791 13.653
R12271 vp_p.n17715 vp_p.n17714 13.653
R12272 vp_p.n17778 vp_p.n17777 13.653
R12273 vp_p.n17720 vp_p.n17719 13.653
R12274 vp_p.n17764 vp_p.n17763 13.653
R12275 vp_p.n17725 vp_p.n17724 13.653
R12276 vp_p.n17750 vp_p.n17749 13.653
R12277 vp_p.n25929 vp_p.n25928 13.653
R12278 vp_p.n24503 vp_p.n24502 13.653
R12279 vp_p.n23081 vp_p.n23080 13.653
R12280 vp_p.n21658 vp_p.n21657 13.653
R12281 vp_p.n20234 vp_p.n20233 13.653
R12282 vp_p.n18809 vp_p.n18808 13.653
R12283 vp_p.n18708 vp_p.n18707 13.653
R12284 vp_p.n18706 vp_p.n18705 13.653
R12285 vp_p.n15951 vp_p.n15950 13.653
R12286 vp_p.n15953 vp_p.n15952 13.653
R12287 vp_p.n14518 vp_p.n14517 13.653
R12288 vp_p.n14520 vp_p.n14519 13.653
R12289 vp_p.n13149 vp_p.n13148 13.653
R12290 vp_p.n13151 vp_p.n13150 13.653
R12291 vp_p.n11715 vp_p.n11714 13.653
R12292 vp_p.n11717 vp_p.n11716 13.653
R12293 vp_p.n10282 vp_p.n10281 13.653
R12294 vp_p.n10284 vp_p.n10283 13.653
R12295 vp_p.n8785 vp_p.n8784 13.653
R12296 vp_p.n8787 vp_p.n8786 13.653
R12297 vp_p.n46 vp_p.n45 13.653
R12298 vp_p.n48 vp_p.n47 13.653
R12299 vp_p.n1423 vp_p.n1422 13.653
R12300 vp_p.n53 vp_p.n52 13.653
R12301 vp_p.n1409 vp_p.n1408 13.653
R12302 vp_p.n58 vp_p.n57 13.653
R12303 vp_p.n1395 vp_p.n1394 13.653
R12304 vp_p.n63 vp_p.n62 13.653
R12305 vp_p.n1381 vp_p.n1380 13.653
R12306 vp_p.n68 vp_p.n67 13.653
R12307 vp_p.n1367 vp_p.n1366 13.653
R12308 vp_p.n73 vp_p.n72 13.653
R12309 vp_p.n1353 vp_p.n1352 13.653
R12310 vp_p.n78 vp_p.n77 13.653
R12311 vp_p.n1339 vp_p.n1338 13.653
R12312 vp_p.n83 vp_p.n82 13.653
R12313 vp_p.n1325 vp_p.n1324 13.653
R12314 vp_p.n88 vp_p.n87 13.653
R12315 vp_p.n1311 vp_p.n1310 13.653
R12316 vp_p.n93 vp_p.n92 13.653
R12317 vp_p.n1297 vp_p.n1296 13.653
R12318 vp_p.n98 vp_p.n97 13.653
R12319 vp_p.n1283 vp_p.n1282 13.653
R12320 vp_p.n103 vp_p.n102 13.653
R12321 vp_p.n1269 vp_p.n1268 13.653
R12322 vp_p.n108 vp_p.n107 13.653
R12323 vp_p.n1255 vp_p.n1254 13.653
R12324 vp_p.n113 vp_p.n112 13.653
R12325 vp_p.n1241 vp_p.n1240 13.653
R12326 vp_p.n118 vp_p.n117 13.653
R12327 vp_p.n1227 vp_p.n1226 13.653
R12328 vp_p.n123 vp_p.n122 13.653
R12329 vp_p.n1213 vp_p.n1212 13.653
R12330 vp_p.n128 vp_p.n127 13.653
R12331 vp_p.n1199 vp_p.n1198 13.653
R12332 vp_p.n133 vp_p.n132 13.653
R12333 vp_p.n1185 vp_p.n1184 13.653
R12334 vp_p.n138 vp_p.n137 13.653
R12335 vp_p.n1171 vp_p.n1170 13.653
R12336 vp_p.n143 vp_p.n142 13.653
R12337 vp_p.n1157 vp_p.n1156 13.653
R12338 vp_p.n148 vp_p.n147 13.653
R12339 vp_p.n1143 vp_p.n1142 13.653
R12340 vp_p.n153 vp_p.n152 13.653
R12341 vp_p.n1129 vp_p.n1128 13.653
R12342 vp_p.n158 vp_p.n157 13.653
R12343 vp_p.n1115 vp_p.n1114 13.653
R12344 vp_p.n163 vp_p.n162 13.653
R12345 vp_p.n1101 vp_p.n1100 13.653
R12346 vp_p.n168 vp_p.n167 13.653
R12347 vp_p.n1087 vp_p.n1086 13.653
R12348 vp_p.n173 vp_p.n172 13.653
R12349 vp_p.n1073 vp_p.n1072 13.653
R12350 vp_p.n178 vp_p.n177 13.653
R12351 vp_p.n1059 vp_p.n1058 13.653
R12352 vp_p.n183 vp_p.n182 13.653
R12353 vp_p.n1045 vp_p.n1044 13.653
R12354 vp_p.n188 vp_p.n187 13.653
R12355 vp_p.n1031 vp_p.n1030 13.653
R12356 vp_p.n193 vp_p.n192 13.653
R12357 vp_p.n1017 vp_p.n1016 13.653
R12358 vp_p.n198 vp_p.n197 13.653
R12359 vp_p.n1003 vp_p.n1002 13.653
R12360 vp_p.n203 vp_p.n202 13.653
R12361 vp_p.n989 vp_p.n988 13.653
R12362 vp_p.n208 vp_p.n207 13.653
R12363 vp_p.n975 vp_p.n974 13.653
R12364 vp_p.n213 vp_p.n212 13.653
R12365 vp_p.n961 vp_p.n960 13.653
R12366 vp_p.n218 vp_p.n217 13.653
R12367 vp_p.n947 vp_p.n946 13.653
R12368 vp_p.n223 vp_p.n222 13.653
R12369 vp_p.n933 vp_p.n932 13.653
R12370 vp_p.n228 vp_p.n227 13.653
R12371 vp_p.n919 vp_p.n918 13.653
R12372 vp_p.n233 vp_p.n232 13.653
R12373 vp_p.n905 vp_p.n904 13.653
R12374 vp_p.n238 vp_p.n237 13.653
R12375 vp_p.n891 vp_p.n890 13.653
R12376 vp_p.n243 vp_p.n242 13.653
R12377 vp_p.n877 vp_p.n876 13.653
R12378 vp_p.n248 vp_p.n247 13.653
R12379 vp_p.n863 vp_p.n862 13.653
R12380 vp_p.n253 vp_p.n252 13.653
R12381 vp_p.n849 vp_p.n848 13.653
R12382 vp_p.n258 vp_p.n257 13.653
R12383 vp_p.n835 vp_p.n834 13.653
R12384 vp_p.n263 vp_p.n262 13.653
R12385 vp_p.n821 vp_p.n820 13.653
R12386 vp_p.n268 vp_p.n267 13.653
R12387 vp_p.n807 vp_p.n806 13.653
R12388 vp_p.n273 vp_p.n272 13.653
R12389 vp_p.n793 vp_p.n792 13.653
R12390 vp_p.n278 vp_p.n277 13.653
R12391 vp_p.n779 vp_p.n778 13.653
R12392 vp_p.n283 vp_p.n282 13.653
R12393 vp_p.n765 vp_p.n764 13.653
R12394 vp_p.n288 vp_p.n287 13.653
R12395 vp_p.n751 vp_p.n750 13.653
R12396 vp_p.n293 vp_p.n292 13.653
R12397 vp_p.n737 vp_p.n736 13.653
R12398 vp_p.n298 vp_p.n297 13.653
R12399 vp_p.n723 vp_p.n722 13.653
R12400 vp_p.n303 vp_p.n302 13.653
R12401 vp_p.n709 vp_p.n708 13.653
R12402 vp_p.n308 vp_p.n307 13.653
R12403 vp_p.n695 vp_p.n694 13.653
R12404 vp_p.n313 vp_p.n312 13.653
R12405 vp_p.n681 vp_p.n680 13.653
R12406 vp_p.n318 vp_p.n317 13.653
R12407 vp_p.n667 vp_p.n666 13.653
R12408 vp_p.n323 vp_p.n322 13.653
R12409 vp_p.n653 vp_p.n652 13.653
R12410 vp_p.n328 vp_p.n327 13.653
R12411 vp_p.n639 vp_p.n638 13.653
R12412 vp_p.n333 vp_p.n332 13.653
R12413 vp_p.n625 vp_p.n624 13.653
R12414 vp_p.n338 vp_p.n337 13.653
R12415 vp_p.n611 vp_p.n610 13.653
R12416 vp_p.n343 vp_p.n342 13.653
R12417 vp_p.n597 vp_p.n596 13.653
R12418 vp_p.n348 vp_p.n347 13.653
R12419 vp_p.n583 vp_p.n582 13.653
R12420 vp_p.n353 vp_p.n352 13.653
R12421 vp_p.n569 vp_p.n568 13.653
R12422 vp_p.n358 vp_p.n357 13.653
R12423 vp_p.n555 vp_p.n554 13.653
R12424 vp_p.n363 vp_p.n362 13.653
R12425 vp_p.n541 vp_p.n540 13.653
R12426 vp_p.n368 vp_p.n367 13.653
R12427 vp_p.n527 vp_p.n526 13.653
R12428 vp_p.n373 vp_p.n372 13.653
R12429 vp_p.n513 vp_p.n512 13.653
R12430 vp_p.n378 vp_p.n377 13.653
R12431 vp_p.n499 vp_p.n498 13.653
R12432 vp_p.n383 vp_p.n382 13.653
R12433 vp_p.n485 vp_p.n484 13.653
R12434 vp_p.n388 vp_p.n387 13.653
R12435 vp_p.n471 vp_p.n470 13.653
R12436 vp_p.n8559 vp_p.n8558 13.653
R12437 vp_p.n7137 vp_p.n7136 13.653
R12438 vp_p.n5714 vp_p.n5713 13.653
R12439 vp_p.n4290 vp_p.n4289 13.653
R12440 vp_p.n2865 vp_p.n2864 13.653
R12441 vp_p.n1437 vp_p.n1436 13.653
R12442 vp_p.n1439 vp_p.n1438 13.653
R12443 vp_p.n8780 vp_p.n8779 13.653
R12444 vp_p.n8782 vp_p.n8781 13.653
R12445 vp_p.n10277 vp_p.n10276 13.653
R12446 vp_p.n10279 vp_p.n10278 13.653
R12447 vp_p.n11710 vp_p.n11709 13.653
R12448 vp_p.n11712 vp_p.n11711 13.653
R12449 vp_p.n13144 vp_p.n13143 13.653
R12450 vp_p.n13146 vp_p.n13145 13.653
R12451 vp_p.n14513 vp_p.n14512 13.653
R12452 vp_p.n14515 vp_p.n14514 13.653
R12453 vp_p.n15946 vp_p.n15945 13.653
R12454 vp_p.n15948 vp_p.n15947 13.653
R12455 vp_p.n17378 vp_p.n17377 13.653
R12456 vp_p.n17380 vp_p.n17379 13.653
R12457 vp_p.n27263 vp_p.n27262 13.653
R12458 vp_p.n25838 vp_p.n25837 13.653
R12459 vp_p.n24416 vp_p.n24415 13.653
R12460 vp_p.n22993 vp_p.n22992 13.653
R12461 vp_p.n21569 vp_p.n21568 13.653
R12462 vp_p.n18806 vp_p.n18805 13.653
R12463 vp_p.n18804 vp_p.n18803 13.653
R12464 vp_p.n18811 vp_p.n18810 13.653
R12465 vp_p.n20128 vp_p.n20127 13.653
R12466 vp_p.n18816 vp_p.n18815 13.653
R12467 vp_p.n20114 vp_p.n20113 13.653
R12468 vp_p.n18821 vp_p.n18820 13.653
R12469 vp_p.n20100 vp_p.n20099 13.653
R12470 vp_p.n18826 vp_p.n18825 13.653
R12471 vp_p.n20086 vp_p.n20085 13.653
R12472 vp_p.n18831 vp_p.n18830 13.653
R12473 vp_p.n20072 vp_p.n20071 13.653
R12474 vp_p.n18836 vp_p.n18835 13.653
R12475 vp_p.n20058 vp_p.n20057 13.653
R12476 vp_p.n18841 vp_p.n18840 13.653
R12477 vp_p.n20044 vp_p.n20043 13.653
R12478 vp_p.n18846 vp_p.n18845 13.653
R12479 vp_p.n20030 vp_p.n20029 13.653
R12480 vp_p.n18851 vp_p.n18850 13.653
R12481 vp_p.n20016 vp_p.n20015 13.653
R12482 vp_p.n18856 vp_p.n18855 13.653
R12483 vp_p.n20002 vp_p.n20001 13.653
R12484 vp_p.n18861 vp_p.n18860 13.653
R12485 vp_p.n19988 vp_p.n19987 13.653
R12486 vp_p.n18866 vp_p.n18865 13.653
R12487 vp_p.n19974 vp_p.n19973 13.653
R12488 vp_p.n18871 vp_p.n18870 13.653
R12489 vp_p.n19960 vp_p.n19959 13.653
R12490 vp_p.n18876 vp_p.n18875 13.653
R12491 vp_p.n19946 vp_p.n19945 13.653
R12492 vp_p.n18881 vp_p.n18880 13.653
R12493 vp_p.n19932 vp_p.n19931 13.653
R12494 vp_p.n18886 vp_p.n18885 13.653
R12495 vp_p.n19918 vp_p.n19917 13.653
R12496 vp_p.n18891 vp_p.n18890 13.653
R12497 vp_p.n19904 vp_p.n19903 13.653
R12498 vp_p.n18896 vp_p.n18895 13.653
R12499 vp_p.n19890 vp_p.n19889 13.653
R12500 vp_p.n18901 vp_p.n18900 13.653
R12501 vp_p.n19876 vp_p.n19875 13.653
R12502 vp_p.n18906 vp_p.n18905 13.653
R12503 vp_p.n19862 vp_p.n19861 13.653
R12504 vp_p.n18911 vp_p.n18910 13.653
R12505 vp_p.n19848 vp_p.n19847 13.653
R12506 vp_p.n18916 vp_p.n18915 13.653
R12507 vp_p.n19834 vp_p.n19833 13.653
R12508 vp_p.n18921 vp_p.n18920 13.653
R12509 vp_p.n19820 vp_p.n19819 13.653
R12510 vp_p.n18926 vp_p.n18925 13.653
R12511 vp_p.n19806 vp_p.n19805 13.653
R12512 vp_p.n18931 vp_p.n18930 13.653
R12513 vp_p.n19792 vp_p.n19791 13.653
R12514 vp_p.n18936 vp_p.n18935 13.653
R12515 vp_p.n19778 vp_p.n19777 13.653
R12516 vp_p.n18941 vp_p.n18940 13.653
R12517 vp_p.n19764 vp_p.n19763 13.653
R12518 vp_p.n18946 vp_p.n18945 13.653
R12519 vp_p.n19750 vp_p.n19749 13.653
R12520 vp_p.n18951 vp_p.n18950 13.653
R12521 vp_p.n19736 vp_p.n19735 13.653
R12522 vp_p.n18956 vp_p.n18955 13.653
R12523 vp_p.n19722 vp_p.n19721 13.653
R12524 vp_p.n18961 vp_p.n18960 13.653
R12525 vp_p.n19708 vp_p.n19707 13.653
R12526 vp_p.n18966 vp_p.n18965 13.653
R12527 vp_p.n19694 vp_p.n19693 13.653
R12528 vp_p.n18971 vp_p.n18970 13.653
R12529 vp_p.n19680 vp_p.n19679 13.653
R12530 vp_p.n18976 vp_p.n18975 13.653
R12531 vp_p.n19666 vp_p.n19665 13.653
R12532 vp_p.n18981 vp_p.n18980 13.653
R12533 vp_p.n19652 vp_p.n19651 13.653
R12534 vp_p.n18986 vp_p.n18985 13.653
R12535 vp_p.n19638 vp_p.n19637 13.653
R12536 vp_p.n18991 vp_p.n18990 13.653
R12537 vp_p.n19624 vp_p.n19623 13.653
R12538 vp_p.n18996 vp_p.n18995 13.653
R12539 vp_p.n19610 vp_p.n19609 13.653
R12540 vp_p.n19001 vp_p.n19000 13.653
R12541 vp_p.n19596 vp_p.n19595 13.653
R12542 vp_p.n19006 vp_p.n19005 13.653
R12543 vp_p.n19582 vp_p.n19581 13.653
R12544 vp_p.n19011 vp_p.n19010 13.653
R12545 vp_p.n19568 vp_p.n19567 13.653
R12546 vp_p.n19016 vp_p.n19015 13.653
R12547 vp_p.n19554 vp_p.n19553 13.653
R12548 vp_p.n19021 vp_p.n19020 13.653
R12549 vp_p.n19540 vp_p.n19539 13.653
R12550 vp_p.n19026 vp_p.n19025 13.653
R12551 vp_p.n19526 vp_p.n19525 13.653
R12552 vp_p.n19031 vp_p.n19030 13.653
R12553 vp_p.n19512 vp_p.n19511 13.653
R12554 vp_p.n19036 vp_p.n19035 13.653
R12555 vp_p.n19498 vp_p.n19497 13.653
R12556 vp_p.n19041 vp_p.n19040 13.653
R12557 vp_p.n19484 vp_p.n19483 13.653
R12558 vp_p.n19046 vp_p.n19045 13.653
R12559 vp_p.n19470 vp_p.n19469 13.653
R12560 vp_p.n19051 vp_p.n19050 13.653
R12561 vp_p.n19456 vp_p.n19455 13.653
R12562 vp_p.n19056 vp_p.n19055 13.653
R12563 vp_p.n19442 vp_p.n19441 13.653
R12564 vp_p.n19061 vp_p.n19060 13.653
R12565 vp_p.n19428 vp_p.n19427 13.653
R12566 vp_p.n19066 vp_p.n19065 13.653
R12567 vp_p.n19414 vp_p.n19413 13.653
R12568 vp_p.n19071 vp_p.n19070 13.653
R12569 vp_p.n19400 vp_p.n19399 13.653
R12570 vp_p.n19076 vp_p.n19075 13.653
R12571 vp_p.n19386 vp_p.n19385 13.653
R12572 vp_p.n19081 vp_p.n19080 13.653
R12573 vp_p.n19372 vp_p.n19371 13.653
R12574 vp_p.n19086 vp_p.n19085 13.653
R12575 vp_p.n19358 vp_p.n19357 13.653
R12576 vp_p.n19091 vp_p.n19090 13.653
R12577 vp_p.n19344 vp_p.n19343 13.653
R12578 vp_p.n19096 vp_p.n19095 13.653
R12579 vp_p.n19330 vp_p.n19329 13.653
R12580 vp_p.n19101 vp_p.n19100 13.653
R12581 vp_p.n19316 vp_p.n19315 13.653
R12582 vp_p.n19106 vp_p.n19105 13.653
R12583 vp_p.n19302 vp_p.n19301 13.653
R12584 vp_p.n19111 vp_p.n19110 13.653
R12585 vp_p.n19288 vp_p.n19287 13.653
R12586 vp_p.n19116 vp_p.n19115 13.653
R12587 vp_p.n19274 vp_p.n19273 13.653
R12588 vp_p.n19121 vp_p.n19120 13.653
R12589 vp_p.n19260 vp_p.n19259 13.653
R12590 vp_p.n19126 vp_p.n19125 13.653
R12591 vp_p.n19246 vp_p.n19245 13.653
R12592 vp_p.n19131 vp_p.n19130 13.653
R12593 vp_p.n19232 vp_p.n19231 13.653
R12594 vp_p.n19136 vp_p.n19135 13.653
R12595 vp_p.n19218 vp_p.n19217 13.653
R12596 vp_p.n19141 vp_p.n19140 13.653
R12597 vp_p.n19204 vp_p.n19203 13.653
R12598 vp_p.n19146 vp_p.n19145 13.653
R12599 vp_p.n19190 vp_p.n19189 13.653
R12600 vp_p.n19151 vp_p.n19150 13.653
R12601 vp_p.n19176 vp_p.n19175 13.653
R12602 vp_p.n25924 vp_p.n25923 13.653
R12603 vp_p.n24498 vp_p.n24497 13.653
R12604 vp_p.n23076 vp_p.n23075 13.653
R12605 vp_p.n21653 vp_p.n21652 13.653
R12606 vp_p.n20229 vp_p.n20228 13.653
R12607 vp_p.n20148 vp_p.n20147 13.653
R12608 vp_p.n20146 vp_p.n20145 13.653
R12609 vp_p.n17373 vp_p.n17372 13.653
R12610 vp_p.n17375 vp_p.n17374 13.653
R12611 vp_p.n15941 vp_p.n15940 13.653
R12612 vp_p.n15943 vp_p.n15942 13.653
R12613 vp_p.n14508 vp_p.n14507 13.653
R12614 vp_p.n14510 vp_p.n14509 13.653
R12615 vp_p.n13139 vp_p.n13138 13.653
R12616 vp_p.n13141 vp_p.n13140 13.653
R12617 vp_p.n11705 vp_p.n11704 13.653
R12618 vp_p.n11707 vp_p.n11706 13.653
R12619 vp_p.n10272 vp_p.n10271 13.653
R12620 vp_p.n10274 vp_p.n10273 13.653
R12621 vp_p.n8775 vp_p.n8774 13.653
R12622 vp_p.n8777 vp_p.n8776 13.653
R12623 vp_p.n41 vp_p.n40 13.653
R12624 vp_p.n43 vp_p.n42 13.653
R12625 vp_p.n1525 vp_p.n1524 13.653
R12626 vp_p.n1527 vp_p.n1526 13.653
R12627 vp_p.n2863 vp_p.n2862 13.653
R12628 vp_p.n1532 vp_p.n1531 13.653
R12629 vp_p.n2849 vp_p.n2848 13.653
R12630 vp_p.n1537 vp_p.n1536 13.653
R12631 vp_p.n2835 vp_p.n2834 13.653
R12632 vp_p.n1542 vp_p.n1541 13.653
R12633 vp_p.n2821 vp_p.n2820 13.653
R12634 vp_p.n1547 vp_p.n1546 13.653
R12635 vp_p.n2807 vp_p.n2806 13.653
R12636 vp_p.n1552 vp_p.n1551 13.653
R12637 vp_p.n2793 vp_p.n2792 13.653
R12638 vp_p.n1557 vp_p.n1556 13.653
R12639 vp_p.n2779 vp_p.n2778 13.653
R12640 vp_p.n1562 vp_p.n1561 13.653
R12641 vp_p.n2765 vp_p.n2764 13.653
R12642 vp_p.n1567 vp_p.n1566 13.653
R12643 vp_p.n2751 vp_p.n2750 13.653
R12644 vp_p.n1572 vp_p.n1571 13.653
R12645 vp_p.n2737 vp_p.n2736 13.653
R12646 vp_p.n1577 vp_p.n1576 13.653
R12647 vp_p.n2723 vp_p.n2722 13.653
R12648 vp_p.n1582 vp_p.n1581 13.653
R12649 vp_p.n2709 vp_p.n2708 13.653
R12650 vp_p.n1587 vp_p.n1586 13.653
R12651 vp_p.n2695 vp_p.n2694 13.653
R12652 vp_p.n1592 vp_p.n1591 13.653
R12653 vp_p.n2681 vp_p.n2680 13.653
R12654 vp_p.n1597 vp_p.n1596 13.653
R12655 vp_p.n2667 vp_p.n2666 13.653
R12656 vp_p.n1602 vp_p.n1601 13.653
R12657 vp_p.n2653 vp_p.n2652 13.653
R12658 vp_p.n1607 vp_p.n1606 13.653
R12659 vp_p.n2639 vp_p.n2638 13.653
R12660 vp_p.n1612 vp_p.n1611 13.653
R12661 vp_p.n2625 vp_p.n2624 13.653
R12662 vp_p.n1617 vp_p.n1616 13.653
R12663 vp_p.n2611 vp_p.n2610 13.653
R12664 vp_p.n1622 vp_p.n1621 13.653
R12665 vp_p.n2597 vp_p.n2596 13.653
R12666 vp_p.n1627 vp_p.n1626 13.653
R12667 vp_p.n2583 vp_p.n2582 13.653
R12668 vp_p.n1632 vp_p.n1631 13.653
R12669 vp_p.n2569 vp_p.n2568 13.653
R12670 vp_p.n1637 vp_p.n1636 13.653
R12671 vp_p.n2555 vp_p.n2554 13.653
R12672 vp_p.n1642 vp_p.n1641 13.653
R12673 vp_p.n2541 vp_p.n2540 13.653
R12674 vp_p.n1647 vp_p.n1646 13.653
R12675 vp_p.n2527 vp_p.n2526 13.653
R12676 vp_p.n1652 vp_p.n1651 13.653
R12677 vp_p.n2513 vp_p.n2512 13.653
R12678 vp_p.n1657 vp_p.n1656 13.653
R12679 vp_p.n2499 vp_p.n2498 13.653
R12680 vp_p.n1662 vp_p.n1661 13.653
R12681 vp_p.n2485 vp_p.n2484 13.653
R12682 vp_p.n1667 vp_p.n1666 13.653
R12683 vp_p.n2471 vp_p.n2470 13.653
R12684 vp_p.n1672 vp_p.n1671 13.653
R12685 vp_p.n2457 vp_p.n2456 13.653
R12686 vp_p.n1677 vp_p.n1676 13.653
R12687 vp_p.n2443 vp_p.n2442 13.653
R12688 vp_p.n1682 vp_p.n1681 13.653
R12689 vp_p.n2429 vp_p.n2428 13.653
R12690 vp_p.n1687 vp_p.n1686 13.653
R12691 vp_p.n2415 vp_p.n2414 13.653
R12692 vp_p.n1692 vp_p.n1691 13.653
R12693 vp_p.n2401 vp_p.n2400 13.653
R12694 vp_p.n1697 vp_p.n1696 13.653
R12695 vp_p.n2387 vp_p.n2386 13.653
R12696 vp_p.n1702 vp_p.n1701 13.653
R12697 vp_p.n2373 vp_p.n2372 13.653
R12698 vp_p.n1707 vp_p.n1706 13.653
R12699 vp_p.n2359 vp_p.n2358 13.653
R12700 vp_p.n1712 vp_p.n1711 13.653
R12701 vp_p.n2345 vp_p.n2344 13.653
R12702 vp_p.n1717 vp_p.n1716 13.653
R12703 vp_p.n2331 vp_p.n2330 13.653
R12704 vp_p.n1722 vp_p.n1721 13.653
R12705 vp_p.n2317 vp_p.n2316 13.653
R12706 vp_p.n1727 vp_p.n1726 13.653
R12707 vp_p.n2303 vp_p.n2302 13.653
R12708 vp_p.n1732 vp_p.n1731 13.653
R12709 vp_p.n2289 vp_p.n2288 13.653
R12710 vp_p.n1737 vp_p.n1736 13.653
R12711 vp_p.n2275 vp_p.n2274 13.653
R12712 vp_p.n1742 vp_p.n1741 13.653
R12713 vp_p.n2261 vp_p.n2260 13.653
R12714 vp_p.n1747 vp_p.n1746 13.653
R12715 vp_p.n2247 vp_p.n2246 13.653
R12716 vp_p.n1752 vp_p.n1751 13.653
R12717 vp_p.n2233 vp_p.n2232 13.653
R12718 vp_p.n1757 vp_p.n1756 13.653
R12719 vp_p.n2219 vp_p.n2218 13.653
R12720 vp_p.n1762 vp_p.n1761 13.653
R12721 vp_p.n2205 vp_p.n2204 13.653
R12722 vp_p.n1767 vp_p.n1766 13.653
R12723 vp_p.n2191 vp_p.n2190 13.653
R12724 vp_p.n1772 vp_p.n1771 13.653
R12725 vp_p.n2177 vp_p.n2176 13.653
R12726 vp_p.n1777 vp_p.n1776 13.653
R12727 vp_p.n2163 vp_p.n2162 13.653
R12728 vp_p.n1782 vp_p.n1781 13.653
R12729 vp_p.n2149 vp_p.n2148 13.653
R12730 vp_p.n1787 vp_p.n1786 13.653
R12731 vp_p.n2135 vp_p.n2134 13.653
R12732 vp_p.n1792 vp_p.n1791 13.653
R12733 vp_p.n2121 vp_p.n2120 13.653
R12734 vp_p.n1797 vp_p.n1796 13.653
R12735 vp_p.n2107 vp_p.n2106 13.653
R12736 vp_p.n1802 vp_p.n1801 13.653
R12737 vp_p.n2093 vp_p.n2092 13.653
R12738 vp_p.n1807 vp_p.n1806 13.653
R12739 vp_p.n2079 vp_p.n2078 13.653
R12740 vp_p.n1812 vp_p.n1811 13.653
R12741 vp_p.n2065 vp_p.n2064 13.653
R12742 vp_p.n1817 vp_p.n1816 13.653
R12743 vp_p.n2051 vp_p.n2050 13.653
R12744 vp_p.n1822 vp_p.n1821 13.653
R12745 vp_p.n2037 vp_p.n2036 13.653
R12746 vp_p.n1827 vp_p.n1826 13.653
R12747 vp_p.n2023 vp_p.n2022 13.653
R12748 vp_p.n1832 vp_p.n1831 13.653
R12749 vp_p.n2009 vp_p.n2008 13.653
R12750 vp_p.n1837 vp_p.n1836 13.653
R12751 vp_p.n1995 vp_p.n1994 13.653
R12752 vp_p.n1842 vp_p.n1841 13.653
R12753 vp_p.n1981 vp_p.n1980 13.653
R12754 vp_p.n1847 vp_p.n1846 13.653
R12755 vp_p.n1967 vp_p.n1966 13.653
R12756 vp_p.n1852 vp_p.n1851 13.653
R12757 vp_p.n1953 vp_p.n1952 13.653
R12758 vp_p.n1857 vp_p.n1856 13.653
R12759 vp_p.n1939 vp_p.n1938 13.653
R12760 vp_p.n1862 vp_p.n1861 13.653
R12761 vp_p.n1925 vp_p.n1924 13.653
R12762 vp_p.n1867 vp_p.n1866 13.653
R12763 vp_p.n1911 vp_p.n1910 13.653
R12764 vp_p.n1872 vp_p.n1871 13.653
R12765 vp_p.n1897 vp_p.n1896 13.653
R12766 vp_p.n8573 vp_p.n8572 13.653
R12767 vp_p.n7151 vp_p.n7150 13.653
R12768 vp_p.n5728 vp_p.n5727 13.653
R12769 vp_p.n4304 vp_p.n4303 13.653
R12770 vp_p.n2877 vp_p.n2876 13.653
R12771 vp_p.n2879 vp_p.n2878 13.653
R12772 vp_p.n36 vp_p.n35 13.653
R12773 vp_p.n38 vp_p.n37 13.653
R12774 vp_p.n8770 vp_p.n8769 13.653
R12775 vp_p.n8772 vp_p.n8771 13.653
R12776 vp_p.n10267 vp_p.n10266 13.653
R12777 vp_p.n10269 vp_p.n10268 13.653
R12778 vp_p.n11700 vp_p.n11699 13.653
R12779 vp_p.n11702 vp_p.n11701 13.653
R12780 vp_p.n13134 vp_p.n13133 13.653
R12781 vp_p.n13136 vp_p.n13135 13.653
R12782 vp_p.n14503 vp_p.n14502 13.653
R12783 vp_p.n14505 vp_p.n14504 13.653
R12784 vp_p.n15936 vp_p.n15935 13.653
R12785 vp_p.n15938 vp_p.n15937 13.653
R12786 vp_p.n17368 vp_p.n17367 13.653
R12787 vp_p.n17370 vp_p.n17369 13.653
R12788 vp_p.n18799 vp_p.n18798 13.653
R12789 vp_p.n18801 vp_p.n18800 13.653
R12790 vp_p.n27277 vp_p.n27276 13.653
R12791 vp_p.n25852 vp_p.n25851 13.653
R12792 vp_p.n24430 vp_p.n24429 13.653
R12793 vp_p.n23007 vp_p.n23006 13.653
R12794 vp_p.n20226 vp_p.n20225 13.653
R12795 vp_p.n20224 vp_p.n20223 13.653
R12796 vp_p.n20231 vp_p.n20230 13.653
R12797 vp_p.n21567 vp_p.n21566 13.653
R12798 vp_p.n20236 vp_p.n20235 13.653
R12799 vp_p.n21553 vp_p.n21552 13.653
R12800 vp_p.n20241 vp_p.n20240 13.653
R12801 vp_p.n21539 vp_p.n21538 13.653
R12802 vp_p.n20246 vp_p.n20245 13.653
R12803 vp_p.n21525 vp_p.n21524 13.653
R12804 vp_p.n20251 vp_p.n20250 13.653
R12805 vp_p.n21511 vp_p.n21510 13.653
R12806 vp_p.n20256 vp_p.n20255 13.653
R12807 vp_p.n21497 vp_p.n21496 13.653
R12808 vp_p.n20261 vp_p.n20260 13.653
R12809 vp_p.n21483 vp_p.n21482 13.653
R12810 vp_p.n20266 vp_p.n20265 13.653
R12811 vp_p.n21469 vp_p.n21468 13.653
R12812 vp_p.n20271 vp_p.n20270 13.653
R12813 vp_p.n21455 vp_p.n21454 13.653
R12814 vp_p.n20276 vp_p.n20275 13.653
R12815 vp_p.n21441 vp_p.n21440 13.653
R12816 vp_p.n20281 vp_p.n20280 13.653
R12817 vp_p.n21427 vp_p.n21426 13.653
R12818 vp_p.n20286 vp_p.n20285 13.653
R12819 vp_p.n21413 vp_p.n21412 13.653
R12820 vp_p.n20291 vp_p.n20290 13.653
R12821 vp_p.n21399 vp_p.n21398 13.653
R12822 vp_p.n20296 vp_p.n20295 13.653
R12823 vp_p.n21385 vp_p.n21384 13.653
R12824 vp_p.n20301 vp_p.n20300 13.653
R12825 vp_p.n21371 vp_p.n21370 13.653
R12826 vp_p.n20306 vp_p.n20305 13.653
R12827 vp_p.n21357 vp_p.n21356 13.653
R12828 vp_p.n20311 vp_p.n20310 13.653
R12829 vp_p.n21343 vp_p.n21342 13.653
R12830 vp_p.n20316 vp_p.n20315 13.653
R12831 vp_p.n21329 vp_p.n21328 13.653
R12832 vp_p.n20321 vp_p.n20320 13.653
R12833 vp_p.n21315 vp_p.n21314 13.653
R12834 vp_p.n20326 vp_p.n20325 13.653
R12835 vp_p.n21301 vp_p.n21300 13.653
R12836 vp_p.n20331 vp_p.n20330 13.653
R12837 vp_p.n21287 vp_p.n21286 13.653
R12838 vp_p.n20336 vp_p.n20335 13.653
R12839 vp_p.n21273 vp_p.n21272 13.653
R12840 vp_p.n20341 vp_p.n20340 13.653
R12841 vp_p.n21259 vp_p.n21258 13.653
R12842 vp_p.n20346 vp_p.n20345 13.653
R12843 vp_p.n21245 vp_p.n21244 13.653
R12844 vp_p.n20351 vp_p.n20350 13.653
R12845 vp_p.n21231 vp_p.n21230 13.653
R12846 vp_p.n20356 vp_p.n20355 13.653
R12847 vp_p.n21217 vp_p.n21216 13.653
R12848 vp_p.n20361 vp_p.n20360 13.653
R12849 vp_p.n21203 vp_p.n21202 13.653
R12850 vp_p.n20366 vp_p.n20365 13.653
R12851 vp_p.n21189 vp_p.n21188 13.653
R12852 vp_p.n20371 vp_p.n20370 13.653
R12853 vp_p.n21175 vp_p.n21174 13.653
R12854 vp_p.n20376 vp_p.n20375 13.653
R12855 vp_p.n21161 vp_p.n21160 13.653
R12856 vp_p.n20381 vp_p.n20380 13.653
R12857 vp_p.n21147 vp_p.n21146 13.653
R12858 vp_p.n20386 vp_p.n20385 13.653
R12859 vp_p.n21133 vp_p.n21132 13.653
R12860 vp_p.n20391 vp_p.n20390 13.653
R12861 vp_p.n21119 vp_p.n21118 13.653
R12862 vp_p.n20396 vp_p.n20395 13.653
R12863 vp_p.n21105 vp_p.n21104 13.653
R12864 vp_p.n20401 vp_p.n20400 13.653
R12865 vp_p.n21091 vp_p.n21090 13.653
R12866 vp_p.n20406 vp_p.n20405 13.653
R12867 vp_p.n21077 vp_p.n21076 13.653
R12868 vp_p.n20411 vp_p.n20410 13.653
R12869 vp_p.n21063 vp_p.n21062 13.653
R12870 vp_p.n20416 vp_p.n20415 13.653
R12871 vp_p.n21049 vp_p.n21048 13.653
R12872 vp_p.n20421 vp_p.n20420 13.653
R12873 vp_p.n21035 vp_p.n21034 13.653
R12874 vp_p.n20426 vp_p.n20425 13.653
R12875 vp_p.n21021 vp_p.n21020 13.653
R12876 vp_p.n20431 vp_p.n20430 13.653
R12877 vp_p.n21007 vp_p.n21006 13.653
R12878 vp_p.n20436 vp_p.n20435 13.653
R12879 vp_p.n20993 vp_p.n20992 13.653
R12880 vp_p.n20441 vp_p.n20440 13.653
R12881 vp_p.n20979 vp_p.n20978 13.653
R12882 vp_p.n20446 vp_p.n20445 13.653
R12883 vp_p.n20965 vp_p.n20964 13.653
R12884 vp_p.n20451 vp_p.n20450 13.653
R12885 vp_p.n20951 vp_p.n20950 13.653
R12886 vp_p.n20456 vp_p.n20455 13.653
R12887 vp_p.n20937 vp_p.n20936 13.653
R12888 vp_p.n20461 vp_p.n20460 13.653
R12889 vp_p.n20923 vp_p.n20922 13.653
R12890 vp_p.n20466 vp_p.n20465 13.653
R12891 vp_p.n20909 vp_p.n20908 13.653
R12892 vp_p.n20471 vp_p.n20470 13.653
R12893 vp_p.n20895 vp_p.n20894 13.653
R12894 vp_p.n20476 vp_p.n20475 13.653
R12895 vp_p.n20881 vp_p.n20880 13.653
R12896 vp_p.n20481 vp_p.n20480 13.653
R12897 vp_p.n20867 vp_p.n20866 13.653
R12898 vp_p.n20486 vp_p.n20485 13.653
R12899 vp_p.n20853 vp_p.n20852 13.653
R12900 vp_p.n20491 vp_p.n20490 13.653
R12901 vp_p.n20839 vp_p.n20838 13.653
R12902 vp_p.n20496 vp_p.n20495 13.653
R12903 vp_p.n20825 vp_p.n20824 13.653
R12904 vp_p.n20501 vp_p.n20500 13.653
R12905 vp_p.n20811 vp_p.n20810 13.653
R12906 vp_p.n20506 vp_p.n20505 13.653
R12907 vp_p.n20797 vp_p.n20796 13.653
R12908 vp_p.n20511 vp_p.n20510 13.653
R12909 vp_p.n20783 vp_p.n20782 13.653
R12910 vp_p.n20516 vp_p.n20515 13.653
R12911 vp_p.n20769 vp_p.n20768 13.653
R12912 vp_p.n20521 vp_p.n20520 13.653
R12913 vp_p.n20755 vp_p.n20754 13.653
R12914 vp_p.n20526 vp_p.n20525 13.653
R12915 vp_p.n20741 vp_p.n20740 13.653
R12916 vp_p.n20531 vp_p.n20530 13.653
R12917 vp_p.n20727 vp_p.n20726 13.653
R12918 vp_p.n20536 vp_p.n20535 13.653
R12919 vp_p.n20713 vp_p.n20712 13.653
R12920 vp_p.n20541 vp_p.n20540 13.653
R12921 vp_p.n20699 vp_p.n20698 13.653
R12922 vp_p.n20546 vp_p.n20545 13.653
R12923 vp_p.n20685 vp_p.n20684 13.653
R12924 vp_p.n20551 vp_p.n20550 13.653
R12925 vp_p.n20671 vp_p.n20670 13.653
R12926 vp_p.n20556 vp_p.n20555 13.653
R12927 vp_p.n20657 vp_p.n20656 13.653
R12928 vp_p.n20561 vp_p.n20560 13.653
R12929 vp_p.n20643 vp_p.n20642 13.653
R12930 vp_p.n20566 vp_p.n20565 13.653
R12931 vp_p.n20629 vp_p.n20628 13.653
R12932 vp_p.n20571 vp_p.n20570 13.653
R12933 vp_p.n20615 vp_p.n20614 13.653
R12934 vp_p.n20576 vp_p.n20575 13.653
R12935 vp_p.n20601 vp_p.n20600 13.653
R12936 vp_p.n25919 vp_p.n25918 13.653
R12937 vp_p.n24493 vp_p.n24492 13.653
R12938 vp_p.n23071 vp_p.n23070 13.653
R12939 vp_p.n21648 vp_p.n21647 13.653
R12940 vp_p.n21587 vp_p.n21586 13.653
R12941 vp_p.n21585 vp_p.n21584 13.653
R12942 vp_p.n18794 vp_p.n18793 13.653
R12943 vp_p.n18796 vp_p.n18795 13.653
R12944 vp_p.n17363 vp_p.n17362 13.653
R12945 vp_p.n17365 vp_p.n17364 13.653
R12946 vp_p.n15931 vp_p.n15930 13.653
R12947 vp_p.n15933 vp_p.n15932 13.653
R12948 vp_p.n14498 vp_p.n14497 13.653
R12949 vp_p.n14500 vp_p.n14499 13.653
R12950 vp_p.n13129 vp_p.n13128 13.653
R12951 vp_p.n13131 vp_p.n13130 13.653
R12952 vp_p.n11695 vp_p.n11694 13.653
R12953 vp_p.n11697 vp_p.n11696 13.653
R12954 vp_p.n10262 vp_p.n10261 13.653
R12955 vp_p.n10264 vp_p.n10263 13.653
R12956 vp_p.n8765 vp_p.n8764 13.653
R12957 vp_p.n8767 vp_p.n8766 13.653
R12958 vp_p.n31 vp_p.n30 13.653
R12959 vp_p.n33 vp_p.n32 13.653
R12960 vp_p.n1520 vp_p.n1519 13.653
R12961 vp_p.n1522 vp_p.n1521 13.653
R12962 vp_p.n2945 vp_p.n2944 13.653
R12963 vp_p.n2947 vp_p.n2946 13.653
R12964 vp_p.n4302 vp_p.n4301 13.653
R12965 vp_p.n2952 vp_p.n2951 13.653
R12966 vp_p.n4288 vp_p.n4287 13.653
R12967 vp_p.n2957 vp_p.n2956 13.653
R12968 vp_p.n4274 vp_p.n4273 13.653
R12969 vp_p.n2962 vp_p.n2961 13.653
R12970 vp_p.n4260 vp_p.n4259 13.653
R12971 vp_p.n2967 vp_p.n2966 13.653
R12972 vp_p.n4246 vp_p.n4245 13.653
R12973 vp_p.n2972 vp_p.n2971 13.653
R12974 vp_p.n4232 vp_p.n4231 13.653
R12975 vp_p.n2977 vp_p.n2976 13.653
R12976 vp_p.n4218 vp_p.n4217 13.653
R12977 vp_p.n2982 vp_p.n2981 13.653
R12978 vp_p.n4204 vp_p.n4203 13.653
R12979 vp_p.n2987 vp_p.n2986 13.653
R12980 vp_p.n4190 vp_p.n4189 13.653
R12981 vp_p.n2992 vp_p.n2991 13.653
R12982 vp_p.n4176 vp_p.n4175 13.653
R12983 vp_p.n2997 vp_p.n2996 13.653
R12984 vp_p.n4162 vp_p.n4161 13.653
R12985 vp_p.n3002 vp_p.n3001 13.653
R12986 vp_p.n4148 vp_p.n4147 13.653
R12987 vp_p.n3007 vp_p.n3006 13.653
R12988 vp_p.n4134 vp_p.n4133 13.653
R12989 vp_p.n3012 vp_p.n3011 13.653
R12990 vp_p.n4120 vp_p.n4119 13.653
R12991 vp_p.n3017 vp_p.n3016 13.653
R12992 vp_p.n4106 vp_p.n4105 13.653
R12993 vp_p.n3022 vp_p.n3021 13.653
R12994 vp_p.n4092 vp_p.n4091 13.653
R12995 vp_p.n3027 vp_p.n3026 13.653
R12996 vp_p.n4078 vp_p.n4077 13.653
R12997 vp_p.n3032 vp_p.n3031 13.653
R12998 vp_p.n4064 vp_p.n4063 13.653
R12999 vp_p.n3037 vp_p.n3036 13.653
R13000 vp_p.n4050 vp_p.n4049 13.653
R13001 vp_p.n3042 vp_p.n3041 13.653
R13002 vp_p.n4036 vp_p.n4035 13.653
R13003 vp_p.n3047 vp_p.n3046 13.653
R13004 vp_p.n4022 vp_p.n4021 13.653
R13005 vp_p.n3052 vp_p.n3051 13.653
R13006 vp_p.n4008 vp_p.n4007 13.653
R13007 vp_p.n3057 vp_p.n3056 13.653
R13008 vp_p.n3994 vp_p.n3993 13.653
R13009 vp_p.n3062 vp_p.n3061 13.653
R13010 vp_p.n3980 vp_p.n3979 13.653
R13011 vp_p.n3067 vp_p.n3066 13.653
R13012 vp_p.n3966 vp_p.n3965 13.653
R13013 vp_p.n3072 vp_p.n3071 13.653
R13014 vp_p.n3952 vp_p.n3951 13.653
R13015 vp_p.n3077 vp_p.n3076 13.653
R13016 vp_p.n3938 vp_p.n3937 13.653
R13017 vp_p.n3082 vp_p.n3081 13.653
R13018 vp_p.n3924 vp_p.n3923 13.653
R13019 vp_p.n3087 vp_p.n3086 13.653
R13020 vp_p.n3910 vp_p.n3909 13.653
R13021 vp_p.n3092 vp_p.n3091 13.653
R13022 vp_p.n3896 vp_p.n3895 13.653
R13023 vp_p.n3097 vp_p.n3096 13.653
R13024 vp_p.n3882 vp_p.n3881 13.653
R13025 vp_p.n3102 vp_p.n3101 13.653
R13026 vp_p.n3868 vp_p.n3867 13.653
R13027 vp_p.n3107 vp_p.n3106 13.653
R13028 vp_p.n3854 vp_p.n3853 13.653
R13029 vp_p.n3112 vp_p.n3111 13.653
R13030 vp_p.n3840 vp_p.n3839 13.653
R13031 vp_p.n3117 vp_p.n3116 13.653
R13032 vp_p.n3826 vp_p.n3825 13.653
R13033 vp_p.n3122 vp_p.n3121 13.653
R13034 vp_p.n3812 vp_p.n3811 13.653
R13035 vp_p.n3127 vp_p.n3126 13.653
R13036 vp_p.n3798 vp_p.n3797 13.653
R13037 vp_p.n3132 vp_p.n3131 13.653
R13038 vp_p.n3784 vp_p.n3783 13.653
R13039 vp_p.n3137 vp_p.n3136 13.653
R13040 vp_p.n3770 vp_p.n3769 13.653
R13041 vp_p.n3142 vp_p.n3141 13.653
R13042 vp_p.n3756 vp_p.n3755 13.653
R13043 vp_p.n3147 vp_p.n3146 13.653
R13044 vp_p.n3742 vp_p.n3741 13.653
R13045 vp_p.n3152 vp_p.n3151 13.653
R13046 vp_p.n3728 vp_p.n3727 13.653
R13047 vp_p.n3157 vp_p.n3156 13.653
R13048 vp_p.n3714 vp_p.n3713 13.653
R13049 vp_p.n3162 vp_p.n3161 13.653
R13050 vp_p.n3700 vp_p.n3699 13.653
R13051 vp_p.n3167 vp_p.n3166 13.653
R13052 vp_p.n3686 vp_p.n3685 13.653
R13053 vp_p.n3172 vp_p.n3171 13.653
R13054 vp_p.n3672 vp_p.n3671 13.653
R13055 vp_p.n3177 vp_p.n3176 13.653
R13056 vp_p.n3658 vp_p.n3657 13.653
R13057 vp_p.n3182 vp_p.n3181 13.653
R13058 vp_p.n3644 vp_p.n3643 13.653
R13059 vp_p.n3187 vp_p.n3186 13.653
R13060 vp_p.n3630 vp_p.n3629 13.653
R13061 vp_p.n3192 vp_p.n3191 13.653
R13062 vp_p.n3616 vp_p.n3615 13.653
R13063 vp_p.n3197 vp_p.n3196 13.653
R13064 vp_p.n3602 vp_p.n3601 13.653
R13065 vp_p.n3202 vp_p.n3201 13.653
R13066 vp_p.n3588 vp_p.n3587 13.653
R13067 vp_p.n3207 vp_p.n3206 13.653
R13068 vp_p.n3574 vp_p.n3573 13.653
R13069 vp_p.n3212 vp_p.n3211 13.653
R13070 vp_p.n3560 vp_p.n3559 13.653
R13071 vp_p.n3217 vp_p.n3216 13.653
R13072 vp_p.n3546 vp_p.n3545 13.653
R13073 vp_p.n3222 vp_p.n3221 13.653
R13074 vp_p.n3532 vp_p.n3531 13.653
R13075 vp_p.n3227 vp_p.n3226 13.653
R13076 vp_p.n3518 vp_p.n3517 13.653
R13077 vp_p.n3232 vp_p.n3231 13.653
R13078 vp_p.n3504 vp_p.n3503 13.653
R13079 vp_p.n3237 vp_p.n3236 13.653
R13080 vp_p.n3490 vp_p.n3489 13.653
R13081 vp_p.n3242 vp_p.n3241 13.653
R13082 vp_p.n3476 vp_p.n3475 13.653
R13083 vp_p.n3247 vp_p.n3246 13.653
R13084 vp_p.n3462 vp_p.n3461 13.653
R13085 vp_p.n3252 vp_p.n3251 13.653
R13086 vp_p.n3448 vp_p.n3447 13.653
R13087 vp_p.n3257 vp_p.n3256 13.653
R13088 vp_p.n3434 vp_p.n3433 13.653
R13089 vp_p.n3262 vp_p.n3261 13.653
R13090 vp_p.n3420 vp_p.n3419 13.653
R13091 vp_p.n3267 vp_p.n3266 13.653
R13092 vp_p.n3406 vp_p.n3405 13.653
R13093 vp_p.n3272 vp_p.n3271 13.653
R13094 vp_p.n3392 vp_p.n3391 13.653
R13095 vp_p.n3277 vp_p.n3276 13.653
R13096 vp_p.n3378 vp_p.n3377 13.653
R13097 vp_p.n3282 vp_p.n3281 13.653
R13098 vp_p.n3364 vp_p.n3363 13.653
R13099 vp_p.n3287 vp_p.n3286 13.653
R13100 vp_p.n3350 vp_p.n3349 13.653
R13101 vp_p.n3292 vp_p.n3291 13.653
R13102 vp_p.n3336 vp_p.n3335 13.653
R13103 vp_p.n3297 vp_p.n3296 13.653
R13104 vp_p.n3322 vp_p.n3321 13.653
R13105 vp_p.n8587 vp_p.n8586 13.653
R13106 vp_p.n7165 vp_p.n7164 13.653
R13107 vp_p.n5742 vp_p.n5741 13.653
R13108 vp_p.n4316 vp_p.n4315 13.653
R13109 vp_p.n4318 vp_p.n4317 13.653
R13110 vp_p.n1515 vp_p.n1514 13.653
R13111 vp_p.n1517 vp_p.n1516 13.653
R13112 vp_p.n26 vp_p.n25 13.653
R13113 vp_p.n28 vp_p.n27 13.653
R13114 vp_p.n8760 vp_p.n8759 13.653
R13115 vp_p.n8762 vp_p.n8761 13.653
R13116 vp_p.n10257 vp_p.n10256 13.653
R13117 vp_p.n10259 vp_p.n10258 13.653
R13118 vp_p.n11690 vp_p.n11689 13.653
R13119 vp_p.n11692 vp_p.n11691 13.653
R13120 vp_p.n13124 vp_p.n13123 13.653
R13121 vp_p.n13126 vp_p.n13125 13.653
R13122 vp_p.n14493 vp_p.n14492 13.653
R13123 vp_p.n14495 vp_p.n14494 13.653
R13124 vp_p.n15926 vp_p.n15925 13.653
R13125 vp_p.n15928 vp_p.n15927 13.653
R13126 vp_p.n17358 vp_p.n17357 13.653
R13127 vp_p.n17360 vp_p.n17359 13.653
R13128 vp_p.n18789 vp_p.n18788 13.653
R13129 vp_p.n18791 vp_p.n18790 13.653
R13130 vp_p.n20219 vp_p.n20218 13.653
R13131 vp_p.n20221 vp_p.n20220 13.653
R13132 vp_p.n27291 vp_p.n27290 13.653
R13133 vp_p.n25866 vp_p.n25865 13.653
R13134 vp_p.n24444 vp_p.n24443 13.653
R13135 vp_p.n21645 vp_p.n21644 13.653
R13136 vp_p.n21643 vp_p.n21642 13.653
R13137 vp_p.n21650 vp_p.n21649 13.653
R13138 vp_p.n23005 vp_p.n23004 13.653
R13139 vp_p.n21655 vp_p.n21654 13.653
R13140 vp_p.n22991 vp_p.n22990 13.653
R13141 vp_p.n21660 vp_p.n21659 13.653
R13142 vp_p.n22977 vp_p.n22976 13.653
R13143 vp_p.n21665 vp_p.n21664 13.653
R13144 vp_p.n22963 vp_p.n22962 13.653
R13145 vp_p.n21670 vp_p.n21669 13.653
R13146 vp_p.n22949 vp_p.n22948 13.653
R13147 vp_p.n21675 vp_p.n21674 13.653
R13148 vp_p.n22935 vp_p.n22934 13.653
R13149 vp_p.n21680 vp_p.n21679 13.653
R13150 vp_p.n22921 vp_p.n22920 13.653
R13151 vp_p.n21685 vp_p.n21684 13.653
R13152 vp_p.n22907 vp_p.n22906 13.653
R13153 vp_p.n21690 vp_p.n21689 13.653
R13154 vp_p.n22893 vp_p.n22892 13.653
R13155 vp_p.n21695 vp_p.n21694 13.653
R13156 vp_p.n22879 vp_p.n22878 13.653
R13157 vp_p.n21700 vp_p.n21699 13.653
R13158 vp_p.n22865 vp_p.n22864 13.653
R13159 vp_p.n21705 vp_p.n21704 13.653
R13160 vp_p.n22851 vp_p.n22850 13.653
R13161 vp_p.n21710 vp_p.n21709 13.653
R13162 vp_p.n22837 vp_p.n22836 13.653
R13163 vp_p.n21715 vp_p.n21714 13.653
R13164 vp_p.n22823 vp_p.n22822 13.653
R13165 vp_p.n21720 vp_p.n21719 13.653
R13166 vp_p.n22809 vp_p.n22808 13.653
R13167 vp_p.n21725 vp_p.n21724 13.653
R13168 vp_p.n22795 vp_p.n22794 13.653
R13169 vp_p.n21730 vp_p.n21729 13.653
R13170 vp_p.n22781 vp_p.n22780 13.653
R13171 vp_p.n21735 vp_p.n21734 13.653
R13172 vp_p.n22767 vp_p.n22766 13.653
R13173 vp_p.n21740 vp_p.n21739 13.653
R13174 vp_p.n22753 vp_p.n22752 13.653
R13175 vp_p.n21745 vp_p.n21744 13.653
R13176 vp_p.n22739 vp_p.n22738 13.653
R13177 vp_p.n21750 vp_p.n21749 13.653
R13178 vp_p.n22725 vp_p.n22724 13.653
R13179 vp_p.n21755 vp_p.n21754 13.653
R13180 vp_p.n22711 vp_p.n22710 13.653
R13181 vp_p.n21760 vp_p.n21759 13.653
R13182 vp_p.n22697 vp_p.n22696 13.653
R13183 vp_p.n21765 vp_p.n21764 13.653
R13184 vp_p.n22683 vp_p.n22682 13.653
R13185 vp_p.n21770 vp_p.n21769 13.653
R13186 vp_p.n22669 vp_p.n22668 13.653
R13187 vp_p.n21775 vp_p.n21774 13.653
R13188 vp_p.n22655 vp_p.n22654 13.653
R13189 vp_p.n21780 vp_p.n21779 13.653
R13190 vp_p.n22641 vp_p.n22640 13.653
R13191 vp_p.n21785 vp_p.n21784 13.653
R13192 vp_p.n22627 vp_p.n22626 13.653
R13193 vp_p.n21790 vp_p.n21789 13.653
R13194 vp_p.n22613 vp_p.n22612 13.653
R13195 vp_p.n21795 vp_p.n21794 13.653
R13196 vp_p.n22599 vp_p.n22598 13.653
R13197 vp_p.n21800 vp_p.n21799 13.653
R13198 vp_p.n22585 vp_p.n22584 13.653
R13199 vp_p.n21805 vp_p.n21804 13.653
R13200 vp_p.n22571 vp_p.n22570 13.653
R13201 vp_p.n21810 vp_p.n21809 13.653
R13202 vp_p.n22557 vp_p.n22556 13.653
R13203 vp_p.n21815 vp_p.n21814 13.653
R13204 vp_p.n22543 vp_p.n22542 13.653
R13205 vp_p.n21820 vp_p.n21819 13.653
R13206 vp_p.n22529 vp_p.n22528 13.653
R13207 vp_p.n21825 vp_p.n21824 13.653
R13208 vp_p.n22515 vp_p.n22514 13.653
R13209 vp_p.n21830 vp_p.n21829 13.653
R13210 vp_p.n22501 vp_p.n22500 13.653
R13211 vp_p.n21835 vp_p.n21834 13.653
R13212 vp_p.n22487 vp_p.n22486 13.653
R13213 vp_p.n21840 vp_p.n21839 13.653
R13214 vp_p.n22473 vp_p.n22472 13.653
R13215 vp_p.n21845 vp_p.n21844 13.653
R13216 vp_p.n22459 vp_p.n22458 13.653
R13217 vp_p.n21850 vp_p.n21849 13.653
R13218 vp_p.n22445 vp_p.n22444 13.653
R13219 vp_p.n21855 vp_p.n21854 13.653
R13220 vp_p.n22431 vp_p.n22430 13.653
R13221 vp_p.n21860 vp_p.n21859 13.653
R13222 vp_p.n22417 vp_p.n22416 13.653
R13223 vp_p.n21865 vp_p.n21864 13.653
R13224 vp_p.n22403 vp_p.n22402 13.653
R13225 vp_p.n21870 vp_p.n21869 13.653
R13226 vp_p.n22389 vp_p.n22388 13.653
R13227 vp_p.n21875 vp_p.n21874 13.653
R13228 vp_p.n22375 vp_p.n22374 13.653
R13229 vp_p.n21880 vp_p.n21879 13.653
R13230 vp_p.n22361 vp_p.n22360 13.653
R13231 vp_p.n21885 vp_p.n21884 13.653
R13232 vp_p.n22347 vp_p.n22346 13.653
R13233 vp_p.n21890 vp_p.n21889 13.653
R13234 vp_p.n22333 vp_p.n22332 13.653
R13235 vp_p.n21895 vp_p.n21894 13.653
R13236 vp_p.n22319 vp_p.n22318 13.653
R13237 vp_p.n21900 vp_p.n21899 13.653
R13238 vp_p.n22305 vp_p.n22304 13.653
R13239 vp_p.n21905 vp_p.n21904 13.653
R13240 vp_p.n22291 vp_p.n22290 13.653
R13241 vp_p.n21910 vp_p.n21909 13.653
R13242 vp_p.n22277 vp_p.n22276 13.653
R13243 vp_p.n21915 vp_p.n21914 13.653
R13244 vp_p.n22263 vp_p.n22262 13.653
R13245 vp_p.n21920 vp_p.n21919 13.653
R13246 vp_p.n22249 vp_p.n22248 13.653
R13247 vp_p.n21925 vp_p.n21924 13.653
R13248 vp_p.n22235 vp_p.n22234 13.653
R13249 vp_p.n21930 vp_p.n21929 13.653
R13250 vp_p.n22221 vp_p.n22220 13.653
R13251 vp_p.n21935 vp_p.n21934 13.653
R13252 vp_p.n22207 vp_p.n22206 13.653
R13253 vp_p.n21940 vp_p.n21939 13.653
R13254 vp_p.n22193 vp_p.n22192 13.653
R13255 vp_p.n21945 vp_p.n21944 13.653
R13256 vp_p.n22179 vp_p.n22178 13.653
R13257 vp_p.n21950 vp_p.n21949 13.653
R13258 vp_p.n22165 vp_p.n22164 13.653
R13259 vp_p.n21955 vp_p.n21954 13.653
R13260 vp_p.n22151 vp_p.n22150 13.653
R13261 vp_p.n21960 vp_p.n21959 13.653
R13262 vp_p.n22137 vp_p.n22136 13.653
R13263 vp_p.n21965 vp_p.n21964 13.653
R13264 vp_p.n22123 vp_p.n22122 13.653
R13265 vp_p.n21970 vp_p.n21969 13.653
R13266 vp_p.n22109 vp_p.n22108 13.653
R13267 vp_p.n21975 vp_p.n21974 13.653
R13268 vp_p.n22095 vp_p.n22094 13.653
R13269 vp_p.n21980 vp_p.n21979 13.653
R13270 vp_p.n22081 vp_p.n22080 13.653
R13271 vp_p.n21985 vp_p.n21984 13.653
R13272 vp_p.n22067 vp_p.n22066 13.653
R13273 vp_p.n21990 vp_p.n21989 13.653
R13274 vp_p.n22053 vp_p.n22052 13.653
R13275 vp_p.n21995 vp_p.n21994 13.653
R13276 vp_p.n22039 vp_p.n22038 13.653
R13277 vp_p.n22000 vp_p.n21999 13.653
R13278 vp_p.n22025 vp_p.n22024 13.653
R13279 vp_p.n25914 vp_p.n25913 13.653
R13280 vp_p.n24488 vp_p.n24487 13.653
R13281 vp_p.n23066 vp_p.n23065 13.653
R13282 vp_p.n23025 vp_p.n23024 13.653
R13283 vp_p.n23023 vp_p.n23022 13.653
R13284 vp_p.n20214 vp_p.n20213 13.653
R13285 vp_p.n20216 vp_p.n20215 13.653
R13286 vp_p.n18784 vp_p.n18783 13.653
R13287 vp_p.n18786 vp_p.n18785 13.653
R13288 vp_p.n17353 vp_p.n17352 13.653
R13289 vp_p.n17355 vp_p.n17354 13.653
R13290 vp_p.n15921 vp_p.n15920 13.653
R13291 vp_p.n15923 vp_p.n15922 13.653
R13292 vp_p.n14488 vp_p.n14487 13.653
R13293 vp_p.n14490 vp_p.n14489 13.653
R13294 vp_p.n13119 vp_p.n13118 13.653
R13295 vp_p.n13121 vp_p.n13120 13.653
R13296 vp_p.n11685 vp_p.n11684 13.653
R13297 vp_p.n11687 vp_p.n11686 13.653
R13298 vp_p.n10252 vp_p.n10251 13.653
R13299 vp_p.n10254 vp_p.n10253 13.653
R13300 vp_p.n8755 vp_p.n8754 13.653
R13301 vp_p.n8757 vp_p.n8756 13.653
R13302 vp_p.n21 vp_p.n20 13.653
R13303 vp_p.n23 vp_p.n22 13.653
R13304 vp_p.n1510 vp_p.n1509 13.653
R13305 vp_p.n1512 vp_p.n1511 13.653
R13306 vp_p.n2940 vp_p.n2939 13.653
R13307 vp_p.n2942 vp_p.n2941 13.653
R13308 vp_p.n4364 vp_p.n4363 13.653
R13309 vp_p.n4366 vp_p.n4365 13.653
R13310 vp_p.n5740 vp_p.n5739 13.653
R13311 vp_p.n4371 vp_p.n4370 13.653
R13312 vp_p.n5726 vp_p.n5725 13.653
R13313 vp_p.n4376 vp_p.n4375 13.653
R13314 vp_p.n5712 vp_p.n5711 13.653
R13315 vp_p.n4381 vp_p.n4380 13.653
R13316 vp_p.n5698 vp_p.n5697 13.653
R13317 vp_p.n4386 vp_p.n4385 13.653
R13318 vp_p.n5684 vp_p.n5683 13.653
R13319 vp_p.n4391 vp_p.n4390 13.653
R13320 vp_p.n5670 vp_p.n5669 13.653
R13321 vp_p.n4396 vp_p.n4395 13.653
R13322 vp_p.n5656 vp_p.n5655 13.653
R13323 vp_p.n4401 vp_p.n4400 13.653
R13324 vp_p.n5642 vp_p.n5641 13.653
R13325 vp_p.n4406 vp_p.n4405 13.653
R13326 vp_p.n5628 vp_p.n5627 13.653
R13327 vp_p.n4411 vp_p.n4410 13.653
R13328 vp_p.n5614 vp_p.n5613 13.653
R13329 vp_p.n4416 vp_p.n4415 13.653
R13330 vp_p.n5600 vp_p.n5599 13.653
R13331 vp_p.n4421 vp_p.n4420 13.653
R13332 vp_p.n5586 vp_p.n5585 13.653
R13333 vp_p.n4426 vp_p.n4425 13.653
R13334 vp_p.n5572 vp_p.n5571 13.653
R13335 vp_p.n4431 vp_p.n4430 13.653
R13336 vp_p.n5558 vp_p.n5557 13.653
R13337 vp_p.n4436 vp_p.n4435 13.653
R13338 vp_p.n5544 vp_p.n5543 13.653
R13339 vp_p.n4441 vp_p.n4440 13.653
R13340 vp_p.n5530 vp_p.n5529 13.653
R13341 vp_p.n4446 vp_p.n4445 13.653
R13342 vp_p.n5516 vp_p.n5515 13.653
R13343 vp_p.n4451 vp_p.n4450 13.653
R13344 vp_p.n5502 vp_p.n5501 13.653
R13345 vp_p.n4456 vp_p.n4455 13.653
R13346 vp_p.n5488 vp_p.n5487 13.653
R13347 vp_p.n4461 vp_p.n4460 13.653
R13348 vp_p.n5474 vp_p.n5473 13.653
R13349 vp_p.n4466 vp_p.n4465 13.653
R13350 vp_p.n5460 vp_p.n5459 13.653
R13351 vp_p.n4471 vp_p.n4470 13.653
R13352 vp_p.n5446 vp_p.n5445 13.653
R13353 vp_p.n4476 vp_p.n4475 13.653
R13354 vp_p.n5432 vp_p.n5431 13.653
R13355 vp_p.n4481 vp_p.n4480 13.653
R13356 vp_p.n5418 vp_p.n5417 13.653
R13357 vp_p.n4486 vp_p.n4485 13.653
R13358 vp_p.n5404 vp_p.n5403 13.653
R13359 vp_p.n4491 vp_p.n4490 13.653
R13360 vp_p.n5390 vp_p.n5389 13.653
R13361 vp_p.n4496 vp_p.n4495 13.653
R13362 vp_p.n5376 vp_p.n5375 13.653
R13363 vp_p.n4501 vp_p.n4500 13.653
R13364 vp_p.n5362 vp_p.n5361 13.653
R13365 vp_p.n4506 vp_p.n4505 13.653
R13366 vp_p.n5348 vp_p.n5347 13.653
R13367 vp_p.n4511 vp_p.n4510 13.653
R13368 vp_p.n5334 vp_p.n5333 13.653
R13369 vp_p.n4516 vp_p.n4515 13.653
R13370 vp_p.n5320 vp_p.n5319 13.653
R13371 vp_p.n4521 vp_p.n4520 13.653
R13372 vp_p.n5306 vp_p.n5305 13.653
R13373 vp_p.n4526 vp_p.n4525 13.653
R13374 vp_p.n5292 vp_p.n5291 13.653
R13375 vp_p.n4531 vp_p.n4530 13.653
R13376 vp_p.n5278 vp_p.n5277 13.653
R13377 vp_p.n4536 vp_p.n4535 13.653
R13378 vp_p.n5264 vp_p.n5263 13.653
R13379 vp_p.n4541 vp_p.n4540 13.653
R13380 vp_p.n5250 vp_p.n5249 13.653
R13381 vp_p.n4546 vp_p.n4545 13.653
R13382 vp_p.n5236 vp_p.n5235 13.653
R13383 vp_p.n4551 vp_p.n4550 13.653
R13384 vp_p.n5222 vp_p.n5221 13.653
R13385 vp_p.n4556 vp_p.n4555 13.653
R13386 vp_p.n5208 vp_p.n5207 13.653
R13387 vp_p.n4561 vp_p.n4560 13.653
R13388 vp_p.n5194 vp_p.n5193 13.653
R13389 vp_p.n4566 vp_p.n4565 13.653
R13390 vp_p.n5180 vp_p.n5179 13.653
R13391 vp_p.n4571 vp_p.n4570 13.653
R13392 vp_p.n5166 vp_p.n5165 13.653
R13393 vp_p.n4576 vp_p.n4575 13.653
R13394 vp_p.n5152 vp_p.n5151 13.653
R13395 vp_p.n4581 vp_p.n4580 13.653
R13396 vp_p.n5138 vp_p.n5137 13.653
R13397 vp_p.n4586 vp_p.n4585 13.653
R13398 vp_p.n5124 vp_p.n5123 13.653
R13399 vp_p.n4591 vp_p.n4590 13.653
R13400 vp_p.n5110 vp_p.n5109 13.653
R13401 vp_p.n4596 vp_p.n4595 13.653
R13402 vp_p.n5096 vp_p.n5095 13.653
R13403 vp_p.n4601 vp_p.n4600 13.653
R13404 vp_p.n5082 vp_p.n5081 13.653
R13405 vp_p.n4606 vp_p.n4605 13.653
R13406 vp_p.n5068 vp_p.n5067 13.653
R13407 vp_p.n4611 vp_p.n4610 13.653
R13408 vp_p.n5054 vp_p.n5053 13.653
R13409 vp_p.n4616 vp_p.n4615 13.653
R13410 vp_p.n5040 vp_p.n5039 13.653
R13411 vp_p.n4621 vp_p.n4620 13.653
R13412 vp_p.n5026 vp_p.n5025 13.653
R13413 vp_p.n4626 vp_p.n4625 13.653
R13414 vp_p.n5012 vp_p.n5011 13.653
R13415 vp_p.n4631 vp_p.n4630 13.653
R13416 vp_p.n4998 vp_p.n4997 13.653
R13417 vp_p.n4636 vp_p.n4635 13.653
R13418 vp_p.n4984 vp_p.n4983 13.653
R13419 vp_p.n4641 vp_p.n4640 13.653
R13420 vp_p.n4970 vp_p.n4969 13.653
R13421 vp_p.n4646 vp_p.n4645 13.653
R13422 vp_p.n4956 vp_p.n4955 13.653
R13423 vp_p.n4651 vp_p.n4650 13.653
R13424 vp_p.n4942 vp_p.n4941 13.653
R13425 vp_p.n4656 vp_p.n4655 13.653
R13426 vp_p.n4928 vp_p.n4927 13.653
R13427 vp_p.n4661 vp_p.n4660 13.653
R13428 vp_p.n4914 vp_p.n4913 13.653
R13429 vp_p.n4666 vp_p.n4665 13.653
R13430 vp_p.n4900 vp_p.n4899 13.653
R13431 vp_p.n4671 vp_p.n4670 13.653
R13432 vp_p.n4886 vp_p.n4885 13.653
R13433 vp_p.n4676 vp_p.n4675 13.653
R13434 vp_p.n4872 vp_p.n4871 13.653
R13435 vp_p.n4681 vp_p.n4680 13.653
R13436 vp_p.n4858 vp_p.n4857 13.653
R13437 vp_p.n4686 vp_p.n4685 13.653
R13438 vp_p.n4844 vp_p.n4843 13.653
R13439 vp_p.n4691 vp_p.n4690 13.653
R13440 vp_p.n4830 vp_p.n4829 13.653
R13441 vp_p.n4696 vp_p.n4695 13.653
R13442 vp_p.n4816 vp_p.n4815 13.653
R13443 vp_p.n4701 vp_p.n4700 13.653
R13444 vp_p.n4802 vp_p.n4801 13.653
R13445 vp_p.n4706 vp_p.n4705 13.653
R13446 vp_p.n4788 vp_p.n4787 13.653
R13447 vp_p.n4711 vp_p.n4710 13.653
R13448 vp_p.n4774 vp_p.n4773 13.653
R13449 vp_p.n4716 vp_p.n4715 13.653
R13450 vp_p.n4760 vp_p.n4759 13.653
R13451 vp_p.n4721 vp_p.n4720 13.653
R13452 vp_p.n4746 vp_p.n4745 13.653
R13453 vp_p.n8601 vp_p.n8600 13.653
R13454 vp_p.n7179 vp_p.n7178 13.653
R13455 vp_p.n5754 vp_p.n5753 13.653
R13456 vp_p.n5756 vp_p.n5755 13.653
R13457 vp_p.n2935 vp_p.n2934 13.653
R13458 vp_p.n2937 vp_p.n2936 13.653
R13459 vp_p.n1505 vp_p.n1504 13.653
R13460 vp_p.n1507 vp_p.n1506 13.653
R13461 vp_p.n16 vp_p.n15 13.653
R13462 vp_p.n18 vp_p.n17 13.653
R13463 vp_p.n8750 vp_p.n8749 13.653
R13464 vp_p.n8752 vp_p.n8751 13.653
R13465 vp_p.n10247 vp_p.n10246 13.653
R13466 vp_p.n10249 vp_p.n10248 13.653
R13467 vp_p.n11680 vp_p.n11679 13.653
R13468 vp_p.n11682 vp_p.n11681 13.653
R13469 vp_p.n13114 vp_p.n13113 13.653
R13470 vp_p.n13116 vp_p.n13115 13.653
R13471 vp_p.n14483 vp_p.n14482 13.653
R13472 vp_p.n14485 vp_p.n14484 13.653
R13473 vp_p.n15916 vp_p.n15915 13.653
R13474 vp_p.n15918 vp_p.n15917 13.653
R13475 vp_p.n17348 vp_p.n17347 13.653
R13476 vp_p.n17350 vp_p.n17349 13.653
R13477 vp_p.n18779 vp_p.n18778 13.653
R13478 vp_p.n18781 vp_p.n18780 13.653
R13479 vp_p.n20209 vp_p.n20208 13.653
R13480 vp_p.n20211 vp_p.n20210 13.653
R13481 vp_p.n21638 vp_p.n21637 13.653
R13482 vp_p.n21640 vp_p.n21639 13.653
R13483 vp_p.n27305 vp_p.n27304 13.653
R13484 vp_p.n25880 vp_p.n25879 13.653
R13485 vp_p.n23063 vp_p.n23062 13.653
R13486 vp_p.n23061 vp_p.n23060 13.653
R13487 vp_p.n23068 vp_p.n23067 13.653
R13488 vp_p.n24442 vp_p.n24441 13.653
R13489 vp_p.n23073 vp_p.n23072 13.653
R13490 vp_p.n24428 vp_p.n24427 13.653
R13491 vp_p.n23078 vp_p.n23077 13.653
R13492 vp_p.n24414 vp_p.n24413 13.653
R13493 vp_p.n23083 vp_p.n23082 13.653
R13494 vp_p.n24400 vp_p.n24399 13.653
R13495 vp_p.n23088 vp_p.n23087 13.653
R13496 vp_p.n24386 vp_p.n24385 13.653
R13497 vp_p.n23093 vp_p.n23092 13.653
R13498 vp_p.n24372 vp_p.n24371 13.653
R13499 vp_p.n23098 vp_p.n23097 13.653
R13500 vp_p.n24358 vp_p.n24357 13.653
R13501 vp_p.n23103 vp_p.n23102 13.653
R13502 vp_p.n24344 vp_p.n24343 13.653
R13503 vp_p.n23108 vp_p.n23107 13.653
R13504 vp_p.n24330 vp_p.n24329 13.653
R13505 vp_p.n23113 vp_p.n23112 13.653
R13506 vp_p.n24316 vp_p.n24315 13.653
R13507 vp_p.n23118 vp_p.n23117 13.653
R13508 vp_p.n24302 vp_p.n24301 13.653
R13509 vp_p.n23123 vp_p.n23122 13.653
R13510 vp_p.n24288 vp_p.n24287 13.653
R13511 vp_p.n23128 vp_p.n23127 13.653
R13512 vp_p.n24274 vp_p.n24273 13.653
R13513 vp_p.n23133 vp_p.n23132 13.653
R13514 vp_p.n24260 vp_p.n24259 13.653
R13515 vp_p.n23138 vp_p.n23137 13.653
R13516 vp_p.n24246 vp_p.n24245 13.653
R13517 vp_p.n23143 vp_p.n23142 13.653
R13518 vp_p.n24232 vp_p.n24231 13.653
R13519 vp_p.n23148 vp_p.n23147 13.653
R13520 vp_p.n24218 vp_p.n24217 13.653
R13521 vp_p.n23153 vp_p.n23152 13.653
R13522 vp_p.n24204 vp_p.n24203 13.653
R13523 vp_p.n23158 vp_p.n23157 13.653
R13524 vp_p.n24190 vp_p.n24189 13.653
R13525 vp_p.n23163 vp_p.n23162 13.653
R13526 vp_p.n24176 vp_p.n24175 13.653
R13527 vp_p.n23168 vp_p.n23167 13.653
R13528 vp_p.n24162 vp_p.n24161 13.653
R13529 vp_p.n23173 vp_p.n23172 13.653
R13530 vp_p.n24148 vp_p.n24147 13.653
R13531 vp_p.n23178 vp_p.n23177 13.653
R13532 vp_p.n24134 vp_p.n24133 13.653
R13533 vp_p.n23183 vp_p.n23182 13.653
R13534 vp_p.n24120 vp_p.n24119 13.653
R13535 vp_p.n23188 vp_p.n23187 13.653
R13536 vp_p.n24106 vp_p.n24105 13.653
R13537 vp_p.n23193 vp_p.n23192 13.653
R13538 vp_p.n24092 vp_p.n24091 13.653
R13539 vp_p.n23198 vp_p.n23197 13.653
R13540 vp_p.n24078 vp_p.n24077 13.653
R13541 vp_p.n23203 vp_p.n23202 13.653
R13542 vp_p.n24064 vp_p.n24063 13.653
R13543 vp_p.n23208 vp_p.n23207 13.653
R13544 vp_p.n24050 vp_p.n24049 13.653
R13545 vp_p.n23213 vp_p.n23212 13.653
R13546 vp_p.n24036 vp_p.n24035 13.653
R13547 vp_p.n23218 vp_p.n23217 13.653
R13548 vp_p.n24022 vp_p.n24021 13.653
R13549 vp_p.n23223 vp_p.n23222 13.653
R13550 vp_p.n24008 vp_p.n24007 13.653
R13551 vp_p.n23228 vp_p.n23227 13.653
R13552 vp_p.n23994 vp_p.n23993 13.653
R13553 vp_p.n23233 vp_p.n23232 13.653
R13554 vp_p.n23980 vp_p.n23979 13.653
R13555 vp_p.n23238 vp_p.n23237 13.653
R13556 vp_p.n23966 vp_p.n23965 13.653
R13557 vp_p.n23243 vp_p.n23242 13.653
R13558 vp_p.n23952 vp_p.n23951 13.653
R13559 vp_p.n23248 vp_p.n23247 13.653
R13560 vp_p.n23938 vp_p.n23937 13.653
R13561 vp_p.n23253 vp_p.n23252 13.653
R13562 vp_p.n23924 vp_p.n23923 13.653
R13563 vp_p.n23258 vp_p.n23257 13.653
R13564 vp_p.n23910 vp_p.n23909 13.653
R13565 vp_p.n23263 vp_p.n23262 13.653
R13566 vp_p.n23896 vp_p.n23895 13.653
R13567 vp_p.n23268 vp_p.n23267 13.653
R13568 vp_p.n23882 vp_p.n23881 13.653
R13569 vp_p.n23273 vp_p.n23272 13.653
R13570 vp_p.n23868 vp_p.n23867 13.653
R13571 vp_p.n23278 vp_p.n23277 13.653
R13572 vp_p.n23854 vp_p.n23853 13.653
R13573 vp_p.n23283 vp_p.n23282 13.653
R13574 vp_p.n23840 vp_p.n23839 13.653
R13575 vp_p.n23288 vp_p.n23287 13.653
R13576 vp_p.n23826 vp_p.n23825 13.653
R13577 vp_p.n23293 vp_p.n23292 13.653
R13578 vp_p.n23812 vp_p.n23811 13.653
R13579 vp_p.n23298 vp_p.n23297 13.653
R13580 vp_p.n23798 vp_p.n23797 13.653
R13581 vp_p.n23303 vp_p.n23302 13.653
R13582 vp_p.n23784 vp_p.n23783 13.653
R13583 vp_p.n23308 vp_p.n23307 13.653
R13584 vp_p.n23770 vp_p.n23769 13.653
R13585 vp_p.n23313 vp_p.n23312 13.653
R13586 vp_p.n23756 vp_p.n23755 13.653
R13587 vp_p.n23318 vp_p.n23317 13.653
R13588 vp_p.n23742 vp_p.n23741 13.653
R13589 vp_p.n23323 vp_p.n23322 13.653
R13590 vp_p.n23728 vp_p.n23727 13.653
R13591 vp_p.n23328 vp_p.n23327 13.653
R13592 vp_p.n23714 vp_p.n23713 13.653
R13593 vp_p.n23333 vp_p.n23332 13.653
R13594 vp_p.n23700 vp_p.n23699 13.653
R13595 vp_p.n23338 vp_p.n23337 13.653
R13596 vp_p.n23686 vp_p.n23685 13.653
R13597 vp_p.n23343 vp_p.n23342 13.653
R13598 vp_p.n23672 vp_p.n23671 13.653
R13599 vp_p.n23348 vp_p.n23347 13.653
R13600 vp_p.n23658 vp_p.n23657 13.653
R13601 vp_p.n23353 vp_p.n23352 13.653
R13602 vp_p.n23644 vp_p.n23643 13.653
R13603 vp_p.n23358 vp_p.n23357 13.653
R13604 vp_p.n23630 vp_p.n23629 13.653
R13605 vp_p.n23363 vp_p.n23362 13.653
R13606 vp_p.n23616 vp_p.n23615 13.653
R13607 vp_p.n23368 vp_p.n23367 13.653
R13608 vp_p.n23602 vp_p.n23601 13.653
R13609 vp_p.n23373 vp_p.n23372 13.653
R13610 vp_p.n23588 vp_p.n23587 13.653
R13611 vp_p.n23378 vp_p.n23377 13.653
R13612 vp_p.n23574 vp_p.n23573 13.653
R13613 vp_p.n23383 vp_p.n23382 13.653
R13614 vp_p.n23560 vp_p.n23559 13.653
R13615 vp_p.n23388 vp_p.n23387 13.653
R13616 vp_p.n23546 vp_p.n23545 13.653
R13617 vp_p.n23393 vp_p.n23392 13.653
R13618 vp_p.n23532 vp_p.n23531 13.653
R13619 vp_p.n23398 vp_p.n23397 13.653
R13620 vp_p.n23518 vp_p.n23517 13.653
R13621 vp_p.n23403 vp_p.n23402 13.653
R13622 vp_p.n23504 vp_p.n23503 13.653
R13623 vp_p.n23408 vp_p.n23407 13.653
R13624 vp_p.n23490 vp_p.n23489 13.653
R13625 vp_p.n23413 vp_p.n23412 13.653
R13626 vp_p.n23476 vp_p.n23475 13.653
R13627 vp_p.n23418 vp_p.n23417 13.653
R13628 vp_p.n23462 vp_p.n23461 13.653
R13629 vp_p.n23423 vp_p.n23422 13.653
R13630 vp_p.n23448 vp_p.n23447 13.653
R13631 vp_p.n25909 vp_p.n25908 13.653
R13632 vp_p.n24483 vp_p.n24482 13.653
R13633 vp_p.n24462 vp_p.n24461 13.653
R13634 vp_p.n24460 vp_p.n24459 13.653
R13635 vp_p.n21633 vp_p.n21632 13.653
R13636 vp_p.n21635 vp_p.n21634 13.653
R13637 vp_p.n20204 vp_p.n20203 13.653
R13638 vp_p.n20206 vp_p.n20205 13.653
R13639 vp_p.n18774 vp_p.n18773 13.653
R13640 vp_p.n18776 vp_p.n18775 13.653
R13641 vp_p.n17343 vp_p.n17342 13.653
R13642 vp_p.n17345 vp_p.n17344 13.653
R13643 vp_p.n15911 vp_p.n15910 13.653
R13644 vp_p.n15913 vp_p.n15912 13.653
R13645 vp_p.n14478 vp_p.n14477 13.653
R13646 vp_p.n14480 vp_p.n14479 13.653
R13647 vp_p.n13109 vp_p.n13108 13.653
R13648 vp_p.n13111 vp_p.n13110 13.653
R13649 vp_p.n11675 vp_p.n11674 13.653
R13650 vp_p.n11677 vp_p.n11676 13.653
R13651 vp_p.n10242 vp_p.n10241 13.653
R13652 vp_p.n10244 vp_p.n10243 13.653
R13653 vp_p.n8745 vp_p.n8744 13.653
R13654 vp_p.n8747 vp_p.n8746 13.653
R13655 vp_p.n11 vp_p.n10 13.653
R13656 vp_p.n13 vp_p.n12 13.653
R13657 vp_p.n1500 vp_p.n1499 13.653
R13658 vp_p.n1502 vp_p.n1501 13.653
R13659 vp_p.n2930 vp_p.n2929 13.653
R13660 vp_p.n2932 vp_p.n2931 13.653
R13661 vp_p.n4359 vp_p.n4358 13.653
R13662 vp_p.n4361 vp_p.n4360 13.653
R13663 vp_p.n5782 vp_p.n5781 13.653
R13664 vp_p.n5784 vp_p.n5783 13.653
R13665 vp_p.n7177 vp_p.n7176 13.653
R13666 vp_p.n5789 vp_p.n5788 13.653
R13667 vp_p.n7163 vp_p.n7162 13.653
R13668 vp_p.n5794 vp_p.n5793 13.653
R13669 vp_p.n7149 vp_p.n7148 13.653
R13670 vp_p.n5799 vp_p.n5798 13.653
R13671 vp_p.n7135 vp_p.n7134 13.653
R13672 vp_p.n5804 vp_p.n5803 13.653
R13673 vp_p.n7121 vp_p.n7120 13.653
R13674 vp_p.n5809 vp_p.n5808 13.653
R13675 vp_p.n7107 vp_p.n7106 13.653
R13676 vp_p.n5814 vp_p.n5813 13.653
R13677 vp_p.n7093 vp_p.n7092 13.653
R13678 vp_p.n5819 vp_p.n5818 13.653
R13679 vp_p.n7079 vp_p.n7078 13.653
R13680 vp_p.n5824 vp_p.n5823 13.653
R13681 vp_p.n7065 vp_p.n7064 13.653
R13682 vp_p.n5829 vp_p.n5828 13.653
R13683 vp_p.n7051 vp_p.n7050 13.653
R13684 vp_p.n5834 vp_p.n5833 13.653
R13685 vp_p.n7037 vp_p.n7036 13.653
R13686 vp_p.n5839 vp_p.n5838 13.653
R13687 vp_p.n7023 vp_p.n7022 13.653
R13688 vp_p.n5844 vp_p.n5843 13.653
R13689 vp_p.n7009 vp_p.n7008 13.653
R13690 vp_p.n5849 vp_p.n5848 13.653
R13691 vp_p.n6995 vp_p.n6994 13.653
R13692 vp_p.n5854 vp_p.n5853 13.653
R13693 vp_p.n6981 vp_p.n6980 13.653
R13694 vp_p.n5859 vp_p.n5858 13.653
R13695 vp_p.n6967 vp_p.n6966 13.653
R13696 vp_p.n5864 vp_p.n5863 13.653
R13697 vp_p.n6953 vp_p.n6952 13.653
R13698 vp_p.n5869 vp_p.n5868 13.653
R13699 vp_p.n6939 vp_p.n6938 13.653
R13700 vp_p.n5874 vp_p.n5873 13.653
R13701 vp_p.n6925 vp_p.n6924 13.653
R13702 vp_p.n5879 vp_p.n5878 13.653
R13703 vp_p.n6911 vp_p.n6910 13.653
R13704 vp_p.n5884 vp_p.n5883 13.653
R13705 vp_p.n6897 vp_p.n6896 13.653
R13706 vp_p.n5889 vp_p.n5888 13.653
R13707 vp_p.n6883 vp_p.n6882 13.653
R13708 vp_p.n5894 vp_p.n5893 13.653
R13709 vp_p.n6869 vp_p.n6868 13.653
R13710 vp_p.n5899 vp_p.n5898 13.653
R13711 vp_p.n6855 vp_p.n6854 13.653
R13712 vp_p.n5904 vp_p.n5903 13.653
R13713 vp_p.n6841 vp_p.n6840 13.653
R13714 vp_p.n5909 vp_p.n5908 13.653
R13715 vp_p.n6827 vp_p.n6826 13.653
R13716 vp_p.n5914 vp_p.n5913 13.653
R13717 vp_p.n6813 vp_p.n6812 13.653
R13718 vp_p.n5919 vp_p.n5918 13.653
R13719 vp_p.n6799 vp_p.n6798 13.653
R13720 vp_p.n5924 vp_p.n5923 13.653
R13721 vp_p.n6785 vp_p.n6784 13.653
R13722 vp_p.n5929 vp_p.n5928 13.653
R13723 vp_p.n6771 vp_p.n6770 13.653
R13724 vp_p.n5934 vp_p.n5933 13.653
R13725 vp_p.n6757 vp_p.n6756 13.653
R13726 vp_p.n5939 vp_p.n5938 13.653
R13727 vp_p.n6743 vp_p.n6742 13.653
R13728 vp_p.n5944 vp_p.n5943 13.653
R13729 vp_p.n6729 vp_p.n6728 13.653
R13730 vp_p.n5949 vp_p.n5948 13.653
R13731 vp_p.n6715 vp_p.n6714 13.653
R13732 vp_p.n5954 vp_p.n5953 13.653
R13733 vp_p.n6701 vp_p.n6700 13.653
R13734 vp_p.n5959 vp_p.n5958 13.653
R13735 vp_p.n6687 vp_p.n6686 13.653
R13736 vp_p.n5964 vp_p.n5963 13.653
R13737 vp_p.n6673 vp_p.n6672 13.653
R13738 vp_p.n5969 vp_p.n5968 13.653
R13739 vp_p.n6659 vp_p.n6658 13.653
R13740 vp_p.n5974 vp_p.n5973 13.653
R13741 vp_p.n6645 vp_p.n6644 13.653
R13742 vp_p.n5979 vp_p.n5978 13.653
R13743 vp_p.n6631 vp_p.n6630 13.653
R13744 vp_p.n5984 vp_p.n5983 13.653
R13745 vp_p.n6617 vp_p.n6616 13.653
R13746 vp_p.n5989 vp_p.n5988 13.653
R13747 vp_p.n6603 vp_p.n6602 13.653
R13748 vp_p.n5994 vp_p.n5993 13.653
R13749 vp_p.n6589 vp_p.n6588 13.653
R13750 vp_p.n5999 vp_p.n5998 13.653
R13751 vp_p.n6575 vp_p.n6574 13.653
R13752 vp_p.n6004 vp_p.n6003 13.653
R13753 vp_p.n6561 vp_p.n6560 13.653
R13754 vp_p.n6009 vp_p.n6008 13.653
R13755 vp_p.n6547 vp_p.n6546 13.653
R13756 vp_p.n6014 vp_p.n6013 13.653
R13757 vp_p.n6533 vp_p.n6532 13.653
R13758 vp_p.n6019 vp_p.n6018 13.653
R13759 vp_p.n6519 vp_p.n6518 13.653
R13760 vp_p.n6024 vp_p.n6023 13.653
R13761 vp_p.n6505 vp_p.n6504 13.653
R13762 vp_p.n6029 vp_p.n6028 13.653
R13763 vp_p.n6491 vp_p.n6490 13.653
R13764 vp_p.n6034 vp_p.n6033 13.653
R13765 vp_p.n6477 vp_p.n6476 13.653
R13766 vp_p.n6039 vp_p.n6038 13.653
R13767 vp_p.n6463 vp_p.n6462 13.653
R13768 vp_p.n6044 vp_p.n6043 13.653
R13769 vp_p.n6449 vp_p.n6448 13.653
R13770 vp_p.n6049 vp_p.n6048 13.653
R13771 vp_p.n6435 vp_p.n6434 13.653
R13772 vp_p.n6054 vp_p.n6053 13.653
R13773 vp_p.n6421 vp_p.n6420 13.653
R13774 vp_p.n6059 vp_p.n6058 13.653
R13775 vp_p.n6407 vp_p.n6406 13.653
R13776 vp_p.n6064 vp_p.n6063 13.653
R13777 vp_p.n6393 vp_p.n6392 13.653
R13778 vp_p.n6069 vp_p.n6068 13.653
R13779 vp_p.n6379 vp_p.n6378 13.653
R13780 vp_p.n6074 vp_p.n6073 13.653
R13781 vp_p.n6365 vp_p.n6364 13.653
R13782 vp_p.n6079 vp_p.n6078 13.653
R13783 vp_p.n6351 vp_p.n6350 13.653
R13784 vp_p.n6084 vp_p.n6083 13.653
R13785 vp_p.n6337 vp_p.n6336 13.653
R13786 vp_p.n6089 vp_p.n6088 13.653
R13787 vp_p.n6323 vp_p.n6322 13.653
R13788 vp_p.n6094 vp_p.n6093 13.653
R13789 vp_p.n6309 vp_p.n6308 13.653
R13790 vp_p.n6099 vp_p.n6098 13.653
R13791 vp_p.n6295 vp_p.n6294 13.653
R13792 vp_p.n6104 vp_p.n6103 13.653
R13793 vp_p.n6281 vp_p.n6280 13.653
R13794 vp_p.n6109 vp_p.n6108 13.653
R13795 vp_p.n6267 vp_p.n6266 13.653
R13796 vp_p.n6114 vp_p.n6113 13.653
R13797 vp_p.n6253 vp_p.n6252 13.653
R13798 vp_p.n6119 vp_p.n6118 13.653
R13799 vp_p.n6239 vp_p.n6238 13.653
R13800 vp_p.n6124 vp_p.n6123 13.653
R13801 vp_p.n6225 vp_p.n6224 13.653
R13802 vp_p.n6129 vp_p.n6128 13.653
R13803 vp_p.n6211 vp_p.n6210 13.653
R13804 vp_p.n6134 vp_p.n6133 13.653
R13805 vp_p.n6197 vp_p.n6196 13.653
R13806 vp_p.n6139 vp_p.n6138 13.653
R13807 vp_p.n6183 vp_p.n6182 13.653
R13808 vp_p.n6144 vp_p.n6143 13.653
R13809 vp_p.n6169 vp_p.n6168 13.653
R13810 vp_p.n8615 vp_p.n8614 13.653
R13811 vp_p.n7191 vp_p.n7190 13.653
R13812 vp_p.n7193 vp_p.n7192 13.653
R13813 vp_p.n4354 vp_p.n4353 13.653
R13814 vp_p.n4356 vp_p.n4355 13.653
R13815 vp_p.n2925 vp_p.n2924 13.653
R13816 vp_p.n2927 vp_p.n2926 13.653
R13817 vp_p.n1495 vp_p.n1494 13.653
R13818 vp_p.n1497 vp_p.n1496 13.653
R13819 vp_p.n6 vp_p.n5 13.653
R13820 vp_p.n8 vp_p.n7 13.653
R13821 vp_p.n8740 vp_p.n8739 13.653
R13822 vp_p.n8742 vp_p.n8741 13.653
R13823 vp_p.n10237 vp_p.n10236 13.653
R13824 vp_p.n10239 vp_p.n10238 13.653
R13825 vp_p.n11670 vp_p.n11669 13.653
R13826 vp_p.n11672 vp_p.n11671 13.653
R13827 vp_p.n13104 vp_p.n13103 13.653
R13828 vp_p.n13106 vp_p.n13105 13.653
R13829 vp_p.n14473 vp_p.n14472 13.653
R13830 vp_p.n14475 vp_p.n14474 13.653
R13831 vp_p.n15906 vp_p.n15905 13.653
R13832 vp_p.n15908 vp_p.n15907 13.653
R13833 vp_p.n17338 vp_p.n17337 13.653
R13834 vp_p.n17340 vp_p.n17339 13.653
R13835 vp_p.n18769 vp_p.n18768 13.653
R13836 vp_p.n18771 vp_p.n18770 13.653
R13837 vp_p.n20199 vp_p.n20198 13.653
R13838 vp_p.n20201 vp_p.n20200 13.653
R13839 vp_p.n21628 vp_p.n21627 13.653
R13840 vp_p.n21630 vp_p.n21629 13.653
R13841 vp_p.n23056 vp_p.n23055 13.653
R13842 vp_p.n23058 vp_p.n23057 13.653
R13843 vp_p.n27319 vp_p.n27318 13.653
R13844 vp_p.n24480 vp_p.n24479 13.653
R13845 vp_p.n24478 vp_p.n24477 13.653
R13846 vp_p.n24485 vp_p.n24484 13.653
R13847 vp_p.n25878 vp_p.n25877 13.653
R13848 vp_p.n24490 vp_p.n24489 13.653
R13849 vp_p.n25864 vp_p.n25863 13.653
R13850 vp_p.n24495 vp_p.n24494 13.653
R13851 vp_p.n25850 vp_p.n25849 13.653
R13852 vp_p.n24500 vp_p.n24499 13.653
R13853 vp_p.n25836 vp_p.n25835 13.653
R13854 vp_p.n24505 vp_p.n24504 13.653
R13855 vp_p.n25822 vp_p.n25821 13.653
R13856 vp_p.n24510 vp_p.n24509 13.653
R13857 vp_p.n25808 vp_p.n25807 13.653
R13858 vp_p.n24515 vp_p.n24514 13.653
R13859 vp_p.n25794 vp_p.n25793 13.653
R13860 vp_p.n24520 vp_p.n24519 13.653
R13861 vp_p.n25780 vp_p.n25779 13.653
R13862 vp_p.n24525 vp_p.n24524 13.653
R13863 vp_p.n25766 vp_p.n25765 13.653
R13864 vp_p.n24530 vp_p.n24529 13.653
R13865 vp_p.n25752 vp_p.n25751 13.653
R13866 vp_p.n24535 vp_p.n24534 13.653
R13867 vp_p.n25738 vp_p.n25737 13.653
R13868 vp_p.n24540 vp_p.n24539 13.653
R13869 vp_p.n25724 vp_p.n25723 13.653
R13870 vp_p.n24545 vp_p.n24544 13.653
R13871 vp_p.n25710 vp_p.n25709 13.653
R13872 vp_p.n24550 vp_p.n24549 13.653
R13873 vp_p.n25696 vp_p.n25695 13.653
R13874 vp_p.n24555 vp_p.n24554 13.653
R13875 vp_p.n25682 vp_p.n25681 13.653
R13876 vp_p.n24560 vp_p.n24559 13.653
R13877 vp_p.n25668 vp_p.n25667 13.653
R13878 vp_p.n24565 vp_p.n24564 13.653
R13879 vp_p.n25654 vp_p.n25653 13.653
R13880 vp_p.n24570 vp_p.n24569 13.653
R13881 vp_p.n25640 vp_p.n25639 13.653
R13882 vp_p.n24575 vp_p.n24574 13.653
R13883 vp_p.n25626 vp_p.n25625 13.653
R13884 vp_p.n24580 vp_p.n24579 13.653
R13885 vp_p.n25612 vp_p.n25611 13.653
R13886 vp_p.n24585 vp_p.n24584 13.653
R13887 vp_p.n25598 vp_p.n25597 13.653
R13888 vp_p.n24590 vp_p.n24589 13.653
R13889 vp_p.n25584 vp_p.n25583 13.653
R13890 vp_p.n24595 vp_p.n24594 13.653
R13891 vp_p.n25570 vp_p.n25569 13.653
R13892 vp_p.n24600 vp_p.n24599 13.653
R13893 vp_p.n25556 vp_p.n25555 13.653
R13894 vp_p.n24605 vp_p.n24604 13.653
R13895 vp_p.n25542 vp_p.n25541 13.653
R13896 vp_p.n24610 vp_p.n24609 13.653
R13897 vp_p.n25528 vp_p.n25527 13.653
R13898 vp_p.n24615 vp_p.n24614 13.653
R13899 vp_p.n25514 vp_p.n25513 13.653
R13900 vp_p.n24620 vp_p.n24619 13.653
R13901 vp_p.n25500 vp_p.n25499 13.653
R13902 vp_p.n24625 vp_p.n24624 13.653
R13903 vp_p.n25486 vp_p.n25485 13.653
R13904 vp_p.n24630 vp_p.n24629 13.653
R13905 vp_p.n25472 vp_p.n25471 13.653
R13906 vp_p.n24635 vp_p.n24634 13.653
R13907 vp_p.n25458 vp_p.n25457 13.653
R13908 vp_p.n24640 vp_p.n24639 13.653
R13909 vp_p.n25444 vp_p.n25443 13.653
R13910 vp_p.n24645 vp_p.n24644 13.653
R13911 vp_p.n25430 vp_p.n25429 13.653
R13912 vp_p.n24650 vp_p.n24649 13.653
R13913 vp_p.n25416 vp_p.n25415 13.653
R13914 vp_p.n24655 vp_p.n24654 13.653
R13915 vp_p.n25402 vp_p.n25401 13.653
R13916 vp_p.n24660 vp_p.n24659 13.653
R13917 vp_p.n25388 vp_p.n25387 13.653
R13918 vp_p.n24665 vp_p.n24664 13.653
R13919 vp_p.n25374 vp_p.n25373 13.653
R13920 vp_p.n24670 vp_p.n24669 13.653
R13921 vp_p.n25360 vp_p.n25359 13.653
R13922 vp_p.n24675 vp_p.n24674 13.653
R13923 vp_p.n25346 vp_p.n25345 13.653
R13924 vp_p.n24680 vp_p.n24679 13.653
R13925 vp_p.n25332 vp_p.n25331 13.653
R13926 vp_p.n24685 vp_p.n24684 13.653
R13927 vp_p.n25318 vp_p.n25317 13.653
R13928 vp_p.n24690 vp_p.n24689 13.653
R13929 vp_p.n25304 vp_p.n25303 13.653
R13930 vp_p.n24695 vp_p.n24694 13.653
R13931 vp_p.n25290 vp_p.n25289 13.653
R13932 vp_p.n24700 vp_p.n24699 13.653
R13933 vp_p.n25276 vp_p.n25275 13.653
R13934 vp_p.n24705 vp_p.n24704 13.653
R13935 vp_p.n25262 vp_p.n25261 13.653
R13936 vp_p.n24710 vp_p.n24709 13.653
R13937 vp_p.n25248 vp_p.n25247 13.653
R13938 vp_p.n24715 vp_p.n24714 13.653
R13939 vp_p.n25234 vp_p.n25233 13.653
R13940 vp_p.n24720 vp_p.n24719 13.653
R13941 vp_p.n25220 vp_p.n25219 13.653
R13942 vp_p.n24725 vp_p.n24724 13.653
R13943 vp_p.n25206 vp_p.n25205 13.653
R13944 vp_p.n24730 vp_p.n24729 13.653
R13945 vp_p.n25192 vp_p.n25191 13.653
R13946 vp_p.n24735 vp_p.n24734 13.653
R13947 vp_p.n25178 vp_p.n25177 13.653
R13948 vp_p.n24740 vp_p.n24739 13.653
R13949 vp_p.n25164 vp_p.n25163 13.653
R13950 vp_p.n24745 vp_p.n24744 13.653
R13951 vp_p.n25150 vp_p.n25149 13.653
R13952 vp_p.n24750 vp_p.n24749 13.653
R13953 vp_p.n25136 vp_p.n25135 13.653
R13954 vp_p.n24755 vp_p.n24754 13.653
R13955 vp_p.n25122 vp_p.n25121 13.653
R13956 vp_p.n24760 vp_p.n24759 13.653
R13957 vp_p.n25108 vp_p.n25107 13.653
R13958 vp_p.n24765 vp_p.n24764 13.653
R13959 vp_p.n25094 vp_p.n25093 13.653
R13960 vp_p.n24770 vp_p.n24769 13.653
R13961 vp_p.n25080 vp_p.n25079 13.653
R13962 vp_p.n24775 vp_p.n24774 13.653
R13963 vp_p.n25066 vp_p.n25065 13.653
R13964 vp_p.n24780 vp_p.n24779 13.653
R13965 vp_p.n25052 vp_p.n25051 13.653
R13966 vp_p.n24785 vp_p.n24784 13.653
R13967 vp_p.n25038 vp_p.n25037 13.653
R13968 vp_p.n24790 vp_p.n24789 13.653
R13969 vp_p.n25024 vp_p.n25023 13.653
R13970 vp_p.n24795 vp_p.n24794 13.653
R13971 vp_p.n25010 vp_p.n25009 13.653
R13972 vp_p.n24800 vp_p.n24799 13.653
R13973 vp_p.n24996 vp_p.n24995 13.653
R13974 vp_p.n24805 vp_p.n24804 13.653
R13975 vp_p.n24982 vp_p.n24981 13.653
R13976 vp_p.n24810 vp_p.n24809 13.653
R13977 vp_p.n24968 vp_p.n24967 13.653
R13978 vp_p.n24815 vp_p.n24814 13.653
R13979 vp_p.n24954 vp_p.n24953 13.653
R13980 vp_p.n24820 vp_p.n24819 13.653
R13981 vp_p.n24940 vp_p.n24939 13.653
R13982 vp_p.n24825 vp_p.n24824 13.653
R13983 vp_p.n24926 vp_p.n24925 13.653
R13984 vp_p.n24830 vp_p.n24829 13.653
R13985 vp_p.n24912 vp_p.n24911 13.653
R13986 vp_p.n24835 vp_p.n24834 13.653
R13987 vp_p.n24898 vp_p.n24897 13.653
R13988 vp_p.n24840 vp_p.n24839 13.653
R13989 vp_p.n24884 vp_p.n24883 13.653
R13990 vp_p.n24845 vp_p.n24844 13.653
R13991 vp_p.n24870 vp_p.n24869 13.653
R13992 vp_p.n25904 vp_p.n25903 13.653
R13993 vp_p.n25898 vp_p.n25897 13.653
R13994 vp_p.n25896 vp_p.n25895 13.653
R13995 vp_p.n23051 vp_p.n23050 13.653
R13996 vp_p.n23053 vp_p.n23052 13.653
R13997 vp_p.n21623 vp_p.n21622 13.653
R13998 vp_p.n21625 vp_p.n21624 13.653
R13999 vp_p.n20194 vp_p.n20193 13.653
R14000 vp_p.n20196 vp_p.n20195 13.653
R14001 vp_p.n18764 vp_p.n18763 13.653
R14002 vp_p.n18766 vp_p.n18765 13.653
R14003 vp_p.n17333 vp_p.n17332 13.653
R14004 vp_p.n17335 vp_p.n17334 13.653
R14005 vp_p.n15901 vp_p.n15900 13.653
R14006 vp_p.n15903 vp_p.n15902 13.653
R14007 vp_p.n14468 vp_p.n14467 13.653
R14008 vp_p.n14470 vp_p.n14469 13.653
R14009 vp_p.n13099 vp_p.n13098 13.653
R14010 vp_p.n13101 vp_p.n13100 13.653
R14011 vp_p.n11665 vp_p.n11664 13.653
R14012 vp_p.n11667 vp_p.n11666 13.653
R14013 vp_p.n10232 vp_p.n10231 13.653
R14014 vp_p.n10234 vp_p.n10233 13.653
R14015 vp_p.n8735 vp_p.n8734 13.653
R14016 vp_p.n8737 vp_p.n8736 13.653
R14017 vp_p.n1 vp_p.n0 13.653
R14018 vp_p.n3 vp_p.n2 13.653
R14019 vp_p.n1490 vp_p.n1489 13.653
R14020 vp_p.n1492 vp_p.n1491 13.653
R14021 vp_p.n2920 vp_p.n2919 13.653
R14022 vp_p.n2922 vp_p.n2921 13.653
R14023 vp_p.n4349 vp_p.n4348 13.653
R14024 vp_p.n4351 vp_p.n4350 13.653
R14025 vp_p.n5777 vp_p.n5776 13.653
R14026 vp_p.n5779 vp_p.n5778 13.653
R14027 vp_p.n8623 vp_p.n8622 13.653
R14028 vp_p.n7591 vp_p.n7590 13.653
R14029 vp_p.n7566 vp_p.n7565 13.653
R14030 vp_p.n7605 vp_p.n7604 13.653
R14031 vp_p.n7561 vp_p.n7560 13.653
R14032 vp_p.n7619 vp_p.n7618 13.653
R14033 vp_p.n7556 vp_p.n7555 13.653
R14034 vp_p.n7633 vp_p.n7632 13.653
R14035 vp_p.n7551 vp_p.n7550 13.653
R14036 vp_p.n7647 vp_p.n7646 13.653
R14037 vp_p.n7546 vp_p.n7545 13.653
R14038 vp_p.n7661 vp_p.n7660 13.653
R14039 vp_p.n7541 vp_p.n7540 13.653
R14040 vp_p.n7675 vp_p.n7674 13.653
R14041 vp_p.n7536 vp_p.n7535 13.653
R14042 vp_p.n7689 vp_p.n7688 13.653
R14043 vp_p.n7531 vp_p.n7530 13.653
R14044 vp_p.n7703 vp_p.n7702 13.653
R14045 vp_p.n7526 vp_p.n7525 13.653
R14046 vp_p.n7717 vp_p.n7716 13.653
R14047 vp_p.n7521 vp_p.n7520 13.653
R14048 vp_p.n7731 vp_p.n7730 13.653
R14049 vp_p.n7516 vp_p.n7515 13.653
R14050 vp_p.n7745 vp_p.n7744 13.653
R14051 vp_p.n7511 vp_p.n7510 13.653
R14052 vp_p.n7759 vp_p.n7758 13.653
R14053 vp_p.n7506 vp_p.n7505 13.653
R14054 vp_p.n7773 vp_p.n7772 13.653
R14055 vp_p.n7501 vp_p.n7500 13.653
R14056 vp_p.n7787 vp_p.n7786 13.653
R14057 vp_p.n7496 vp_p.n7495 13.653
R14058 vp_p.n7801 vp_p.n7800 13.653
R14059 vp_p.n7491 vp_p.n7490 13.653
R14060 vp_p.n7815 vp_p.n7814 13.653
R14061 vp_p.n7486 vp_p.n7485 13.653
R14062 vp_p.n7829 vp_p.n7828 13.653
R14063 vp_p.n7481 vp_p.n7480 13.653
R14064 vp_p.n7843 vp_p.n7842 13.653
R14065 vp_p.n7476 vp_p.n7475 13.653
R14066 vp_p.n7857 vp_p.n7856 13.653
R14067 vp_p.n7471 vp_p.n7470 13.653
R14068 vp_p.n7871 vp_p.n7870 13.653
R14069 vp_p.n7466 vp_p.n7465 13.653
R14070 vp_p.n7885 vp_p.n7884 13.653
R14071 vp_p.n7461 vp_p.n7460 13.653
R14072 vp_p.n7899 vp_p.n7898 13.653
R14073 vp_p.n7456 vp_p.n7455 13.653
R14074 vp_p.n7913 vp_p.n7912 13.653
R14075 vp_p.n7451 vp_p.n7450 13.653
R14076 vp_p.n7927 vp_p.n7926 13.653
R14077 vp_p.n7446 vp_p.n7445 13.653
R14078 vp_p.n7941 vp_p.n7940 13.653
R14079 vp_p.n7441 vp_p.n7440 13.653
R14080 vp_p.n7955 vp_p.n7954 13.653
R14081 vp_p.n7436 vp_p.n7435 13.653
R14082 vp_p.n7969 vp_p.n7968 13.653
R14083 vp_p.n7431 vp_p.n7430 13.653
R14084 vp_p.n7983 vp_p.n7982 13.653
R14085 vp_p.n7426 vp_p.n7425 13.653
R14086 vp_p.n7997 vp_p.n7996 13.653
R14087 vp_p.n7421 vp_p.n7420 13.653
R14088 vp_p.n8011 vp_p.n8010 13.653
R14089 vp_p.n7416 vp_p.n7415 13.653
R14090 vp_p.n8025 vp_p.n8024 13.653
R14091 vp_p.n7411 vp_p.n7410 13.653
R14092 vp_p.n8039 vp_p.n8038 13.653
R14093 vp_p.n7406 vp_p.n7405 13.653
R14094 vp_p.n8053 vp_p.n8052 13.653
R14095 vp_p.n7401 vp_p.n7400 13.653
R14096 vp_p.n8067 vp_p.n8066 13.653
R14097 vp_p.n7396 vp_p.n7395 13.653
R14098 vp_p.n8081 vp_p.n8080 13.653
R14099 vp_p.n7391 vp_p.n7390 13.653
R14100 vp_p.n8095 vp_p.n8094 13.653
R14101 vp_p.n7386 vp_p.n7385 13.653
R14102 vp_p.n8109 vp_p.n8108 13.653
R14103 vp_p.n7381 vp_p.n7380 13.653
R14104 vp_p.n8123 vp_p.n8122 13.653
R14105 vp_p.n7376 vp_p.n7375 13.653
R14106 vp_p.n8137 vp_p.n8136 13.653
R14107 vp_p.n7371 vp_p.n7370 13.653
R14108 vp_p.n8151 vp_p.n8150 13.653
R14109 vp_p.n7366 vp_p.n7365 13.653
R14110 vp_p.n8165 vp_p.n8164 13.653
R14111 vp_p.n7361 vp_p.n7360 13.653
R14112 vp_p.n8179 vp_p.n8178 13.653
R14113 vp_p.n7356 vp_p.n7355 13.653
R14114 vp_p.n8193 vp_p.n8192 13.653
R14115 vp_p.n7351 vp_p.n7350 13.653
R14116 vp_p.n8207 vp_p.n8206 13.653
R14117 vp_p.n7346 vp_p.n7345 13.653
R14118 vp_p.n8221 vp_p.n8220 13.653
R14119 vp_p.n7341 vp_p.n7340 13.653
R14120 vp_p.n8235 vp_p.n8234 13.653
R14121 vp_p.n7336 vp_p.n7335 13.653
R14122 vp_p.n8249 vp_p.n8248 13.653
R14123 vp_p.n7331 vp_p.n7330 13.653
R14124 vp_p.n8263 vp_p.n8262 13.653
R14125 vp_p.n7326 vp_p.n7325 13.653
R14126 vp_p.n8277 vp_p.n8276 13.653
R14127 vp_p.n7321 vp_p.n7320 13.653
R14128 vp_p.n8291 vp_p.n8290 13.653
R14129 vp_p.n7316 vp_p.n7315 13.653
R14130 vp_p.n8305 vp_p.n8304 13.653
R14131 vp_p.n7311 vp_p.n7310 13.653
R14132 vp_p.n8319 vp_p.n8318 13.653
R14133 vp_p.n7306 vp_p.n7305 13.653
R14134 vp_p.n8333 vp_p.n8332 13.653
R14135 vp_p.n7301 vp_p.n7300 13.653
R14136 vp_p.n8347 vp_p.n8346 13.653
R14137 vp_p.n7296 vp_p.n7295 13.653
R14138 vp_p.n8361 vp_p.n8360 13.653
R14139 vp_p.n7291 vp_p.n7290 13.653
R14140 vp_p.n8375 vp_p.n8374 13.653
R14141 vp_p.n7286 vp_p.n7285 13.653
R14142 vp_p.n8389 vp_p.n8388 13.653
R14143 vp_p.n7281 vp_p.n7280 13.653
R14144 vp_p.n8403 vp_p.n8402 13.653
R14145 vp_p.n7276 vp_p.n7275 13.653
R14146 vp_p.n8417 vp_p.n8416 13.653
R14147 vp_p.n7271 vp_p.n7270 13.653
R14148 vp_p.n8431 vp_p.n8430 13.653
R14149 vp_p.n7266 vp_p.n7265 13.653
R14150 vp_p.n8445 vp_p.n8444 13.653
R14151 vp_p.n7261 vp_p.n7260 13.653
R14152 vp_p.n8459 vp_p.n8458 13.653
R14153 vp_p.n7256 vp_p.n7255 13.653
R14154 vp_p.n8473 vp_p.n8472 13.653
R14155 vp_p.n7251 vp_p.n7250 13.653
R14156 vp_p.n8487 vp_p.n8486 13.653
R14157 vp_p.n7246 vp_p.n7245 13.653
R14158 vp_p.n8501 vp_p.n8500 13.653
R14159 vp_p.n7241 vp_p.n7240 13.653
R14160 vp_p.n8515 vp_p.n8514 13.653
R14161 vp_p.n7236 vp_p.n7235 13.653
R14162 vp_p.n8529 vp_p.n8528 13.653
R14163 vp_p.n7231 vp_p.n7230 13.653
R14164 vp_p.n8543 vp_p.n8542 13.653
R14165 vp_p.n7226 vp_p.n7225 13.653
R14166 vp_p.n8557 vp_p.n8556 13.653
R14167 vp_p.n7221 vp_p.n7220 13.653
R14168 vp_p.n8571 vp_p.n8570 13.653
R14169 vp_p.n7216 vp_p.n7215 13.653
R14170 vp_p.n8585 vp_p.n8584 13.653
R14171 vp_p.n7211 vp_p.n7210 13.653
R14172 vp_p.n8599 vp_p.n8598 13.653
R14173 vp_p.n7206 vp_p.n7205 13.653
R14174 vp_p.n8613 vp_p.n8612 13.653
R14175 vp_p.n8625 vp_p.n8624 13.653
R14176 vp_p.n7583 vp_p.n7582 13.653
R14177 vp_p.n7581 vp_p.n7580 13.653
R14178 vp_p.n6147 vp_p.n6146 13.653
R14179 vp_p.n6149 vp_p.n6148 13.653
R14180 vp_p.n4724 vp_p.n4723 13.653
R14181 vp_p.n4726 vp_p.n4725 13.653
R14182 vp_p.n3300 vp_p.n3299 13.653
R14183 vp_p.n3302 vp_p.n3301 13.653
R14184 vp_p.n1875 vp_p.n1874 13.653
R14185 vp_p.n1877 vp_p.n1876 13.653
R14186 vp_p.n391 vp_p.n390 13.653
R14187 vp_p.n393 vp_p.n392 13.653
R14188 vp_p.n9130 vp_p.n9129 13.653
R14189 vp_p.n9132 vp_p.n9131 13.653
R14190 vp_p.n10632 vp_p.n10631 13.653
R14191 vp_p.n10634 vp_p.n10633 13.653
R14192 vp_p.n12070 vp_p.n12069 13.653
R14193 vp_p.n12072 vp_p.n12071 13.653
R14194 vp_p.n13834 vp_p.n13833 13.653
R14195 vp_p.n13836 vp_p.n13835 13.653
R14196 vp_p.n14873 vp_p.n14872 13.653
R14197 vp_p.n14875 vp_p.n14874 13.653
R14198 vp_p.n16301 vp_p.n16300 13.653
R14199 vp_p.n16303 vp_p.n16302 13.653
R14200 vp_p.n17728 vp_p.n17727 13.653
R14201 vp_p.n17730 vp_p.n17729 13.653
R14202 vp_p.n19154 vp_p.n19153 13.653
R14203 vp_p.n19156 vp_p.n19155 13.653
R14204 vp_p.n20579 vp_p.n20578 13.653
R14205 vp_p.n20581 vp_p.n20580 13.653
R14206 vp_p.n22003 vp_p.n22002 13.653
R14207 vp_p.n22005 vp_p.n22004 13.653
R14208 vp_p.n23426 vp_p.n23425 13.653
R14209 vp_p.n23428 vp_p.n23427 13.653
R14210 vp_p.n24848 vp_p.n24847 13.653
R14211 vp_p.n24850 vp_p.n24849 13.653
R14212 vp_p.n26274 vp_p.n26273 13.653
R14213 vp_p.n26276 vp_p.n26275 13.653
R14214 vp_p.n26295 vp_p.n26294 13.653
R14215 vp_p.n26271 vp_p.n26270 13.653
R14216 vp_p.n26309 vp_p.n26308 13.653
R14217 vp_p.n26266 vp_p.n26265 13.653
R14218 vp_p.n26323 vp_p.n26322 13.653
R14219 vp_p.n26261 vp_p.n26260 13.653
R14220 vp_p.n26337 vp_p.n26336 13.653
R14221 vp_p.n26256 vp_p.n26255 13.653
R14222 vp_p.n26351 vp_p.n26350 13.653
R14223 vp_p.n26251 vp_p.n26250 13.653
R14224 vp_p.n26365 vp_p.n26364 13.653
R14225 vp_p.n26246 vp_p.n26245 13.653
R14226 vp_p.n26379 vp_p.n26378 13.653
R14227 vp_p.n26241 vp_p.n26240 13.653
R14228 vp_p.n26393 vp_p.n26392 13.653
R14229 vp_p.n26236 vp_p.n26235 13.653
R14230 vp_p.n26407 vp_p.n26406 13.653
R14231 vp_p.n26231 vp_p.n26230 13.653
R14232 vp_p.n26421 vp_p.n26420 13.653
R14233 vp_p.n26226 vp_p.n26225 13.653
R14234 vp_p.n26435 vp_p.n26434 13.653
R14235 vp_p.n26221 vp_p.n26220 13.653
R14236 vp_p.n26449 vp_p.n26448 13.653
R14237 vp_p.n26216 vp_p.n26215 13.653
R14238 vp_p.n26463 vp_p.n26462 13.653
R14239 vp_p.n26211 vp_p.n26210 13.653
R14240 vp_p.n26477 vp_p.n26476 13.653
R14241 vp_p.n26206 vp_p.n26205 13.653
R14242 vp_p.n26491 vp_p.n26490 13.653
R14243 vp_p.n26201 vp_p.n26200 13.653
R14244 vp_p.n26505 vp_p.n26504 13.653
R14245 vp_p.n26196 vp_p.n26195 13.653
R14246 vp_p.n26519 vp_p.n26518 13.653
R14247 vp_p.n26191 vp_p.n26190 13.653
R14248 vp_p.n26533 vp_p.n26532 13.653
R14249 vp_p.n26186 vp_p.n26185 13.653
R14250 vp_p.n26547 vp_p.n26546 13.653
R14251 vp_p.n26181 vp_p.n26180 13.653
R14252 vp_p.n26561 vp_p.n26560 13.653
R14253 vp_p.n26176 vp_p.n26175 13.653
R14254 vp_p.n26575 vp_p.n26574 13.653
R14255 vp_p.n26171 vp_p.n26170 13.653
R14256 vp_p.n26589 vp_p.n26588 13.653
R14257 vp_p.n26166 vp_p.n26165 13.653
R14258 vp_p.n26603 vp_p.n26602 13.653
R14259 vp_p.n26161 vp_p.n26160 13.653
R14260 vp_p.n26617 vp_p.n26616 13.653
R14261 vp_p.n26156 vp_p.n26155 13.653
R14262 vp_p.n26631 vp_p.n26630 13.653
R14263 vp_p.n26151 vp_p.n26150 13.653
R14264 vp_p.n26645 vp_p.n26644 13.653
R14265 vp_p.n26146 vp_p.n26145 13.653
R14266 vp_p.n26659 vp_p.n26658 13.653
R14267 vp_p.n26141 vp_p.n26140 13.653
R14268 vp_p.n26673 vp_p.n26672 13.653
R14269 vp_p.n26136 vp_p.n26135 13.653
R14270 vp_p.n26687 vp_p.n26686 13.653
R14271 vp_p.n26131 vp_p.n26130 13.653
R14272 vp_p.n26701 vp_p.n26700 13.653
R14273 vp_p.n26126 vp_p.n26125 13.653
R14274 vp_p.n26715 vp_p.n26714 13.653
R14275 vp_p.n26121 vp_p.n26120 13.653
R14276 vp_p.n26729 vp_p.n26728 13.653
R14277 vp_p.n26116 vp_p.n26115 13.653
R14278 vp_p.n26743 vp_p.n26742 13.653
R14279 vp_p.n26111 vp_p.n26110 13.653
R14280 vp_p.n26757 vp_p.n26756 13.653
R14281 vp_p.n26106 vp_p.n26105 13.653
R14282 vp_p.n26771 vp_p.n26770 13.653
R14283 vp_p.n26101 vp_p.n26100 13.653
R14284 vp_p.n26785 vp_p.n26784 13.653
R14285 vp_p.n26096 vp_p.n26095 13.653
R14286 vp_p.n26799 vp_p.n26798 13.653
R14287 vp_p.n26091 vp_p.n26090 13.653
R14288 vp_p.n26813 vp_p.n26812 13.653
R14289 vp_p.n26086 vp_p.n26085 13.653
R14290 vp_p.n26827 vp_p.n26826 13.653
R14291 vp_p.n26081 vp_p.n26080 13.653
R14292 vp_p.n26841 vp_p.n26840 13.653
R14293 vp_p.n26076 vp_p.n26075 13.653
R14294 vp_p.n26855 vp_p.n26854 13.653
R14295 vp_p.n26071 vp_p.n26070 13.653
R14296 vp_p.n26869 vp_p.n26868 13.653
R14297 vp_p.n26066 vp_p.n26065 13.653
R14298 vp_p.n26883 vp_p.n26882 13.653
R14299 vp_p.n26061 vp_p.n26060 13.653
R14300 vp_p.n26897 vp_p.n26896 13.653
R14301 vp_p.n26056 vp_p.n26055 13.653
R14302 vp_p.n26911 vp_p.n26910 13.653
R14303 vp_p.n26051 vp_p.n26050 13.653
R14304 vp_p.n26925 vp_p.n26924 13.653
R14305 vp_p.n26046 vp_p.n26045 13.653
R14306 vp_p.n26939 vp_p.n26938 13.653
R14307 vp_p.n26041 vp_p.n26040 13.653
R14308 vp_p.n26953 vp_p.n26952 13.653
R14309 vp_p.n26036 vp_p.n26035 13.653
R14310 vp_p.n26967 vp_p.n26966 13.653
R14311 vp_p.n26031 vp_p.n26030 13.653
R14312 vp_p.n26981 vp_p.n26980 13.653
R14313 vp_p.n26026 vp_p.n26025 13.653
R14314 vp_p.n26995 vp_p.n26994 13.653
R14315 vp_p.n26021 vp_p.n26020 13.653
R14316 vp_p.n27009 vp_p.n27008 13.653
R14317 vp_p.n26016 vp_p.n26015 13.653
R14318 vp_p.n27023 vp_p.n27022 13.653
R14319 vp_p.n26011 vp_p.n26010 13.653
R14320 vp_p.n27037 vp_p.n27036 13.653
R14321 vp_p.n26006 vp_p.n26005 13.653
R14322 vp_p.n27051 vp_p.n27050 13.653
R14323 vp_p.n26001 vp_p.n26000 13.653
R14324 vp_p.n27065 vp_p.n27064 13.653
R14325 vp_p.n25996 vp_p.n25995 13.653
R14326 vp_p.n27079 vp_p.n27078 13.653
R14327 vp_p.n25991 vp_p.n25990 13.653
R14328 vp_p.n27093 vp_p.n27092 13.653
R14329 vp_p.n25986 vp_p.n25985 13.653
R14330 vp_p.n27107 vp_p.n27106 13.653
R14331 vp_p.n25981 vp_p.n25980 13.653
R14332 vp_p.n27121 vp_p.n27120 13.653
R14333 vp_p.n25976 vp_p.n25975 13.653
R14334 vp_p.n27135 vp_p.n27134 13.653
R14335 vp_p.n25971 vp_p.n25970 13.653
R14336 vp_p.n27149 vp_p.n27148 13.653
R14337 vp_p.n25966 vp_p.n25965 13.653
R14338 vp_p.n27163 vp_p.n27162 13.653
R14339 vp_p.n25961 vp_p.n25960 13.653
R14340 vp_p.n27177 vp_p.n27176 13.653
R14341 vp_p.n25956 vp_p.n25955 13.653
R14342 vp_p.n27191 vp_p.n27190 13.653
R14343 vp_p.n25951 vp_p.n25950 13.653
R14344 vp_p.n27205 vp_p.n27204 13.653
R14345 vp_p.n25946 vp_p.n25945 13.653
R14346 vp_p.n27219 vp_p.n27218 13.653
R14347 vp_p.n25941 vp_p.n25940 13.653
R14348 vp_p.n27233 vp_p.n27232 13.653
R14349 vp_p.n25936 vp_p.n25935 13.653
R14350 vp_p.n27247 vp_p.n27246 13.653
R14351 vp_p.n25931 vp_p.n25930 13.653
R14352 vp_p.n27261 vp_p.n27260 13.653
R14353 vp_p.n25926 vp_p.n25925 13.653
R14354 vp_p.n27275 vp_p.n27274 13.653
R14355 vp_p.n25921 vp_p.n25920 13.653
R14356 vp_p.n27289 vp_p.n27288 13.653
R14357 vp_p.n25916 vp_p.n25915 13.653
R14358 vp_p.n27303 vp_p.n27302 13.653
R14359 vp_p.n25911 vp_p.n25910 13.653
R14360 vp_p.n27317 vp_p.n27316 13.653
R14361 vp_p.n25906 vp_p.n25905 13.653
R14362 vp_p.n26283 vp_p.n26282 13.653
R14363 vp_p.n26281 vp_p.n26280 13.653
R14364 vp_p.n24853 vp_p.n24852 13.653
R14365 vp_p.n24855 vp_p.n24854 13.653
R14366 vp_p.n23431 vp_p.n23430 13.653
R14367 vp_p.n23433 vp_p.n23432 13.653
R14368 vp_p.n22008 vp_p.n22007 13.653
R14369 vp_p.n22010 vp_p.n22009 13.653
R14370 vp_p.n20584 vp_p.n20583 13.653
R14371 vp_p.n20586 vp_p.n20585 13.653
R14372 vp_p.n19159 vp_p.n19158 13.653
R14373 vp_p.n19161 vp_p.n19160 13.653
R14374 vp_p.n17733 vp_p.n17732 13.653
R14375 vp_p.n17735 vp_p.n17734 13.653
R14376 vp_p.n16306 vp_p.n16305 13.653
R14377 vp_p.n16308 vp_p.n16307 13.653
R14378 vp_p.n14878 vp_p.n14877 13.653
R14379 vp_p.n14880 vp_p.n14879 13.653
R14380 vp_p.n13839 vp_p.n13838 13.653
R14381 vp_p.n13841 vp_p.n13840 13.653
R14382 vp_p.n12075 vp_p.n12074 13.653
R14383 vp_p.n12077 vp_p.n12076 13.653
R14384 vp_p.n10637 vp_p.n10636 13.653
R14385 vp_p.n10639 vp_p.n10638 13.653
R14386 vp_p.n9135 vp_p.n9134 13.653
R14387 vp_p.n9137 vp_p.n9136 13.653
R14388 vp_p.n396 vp_p.n395 13.653
R14389 vp_p.n398 vp_p.n397 13.653
R14390 vp_p.n1880 vp_p.n1879 13.653
R14391 vp_p.n1882 vp_p.n1881 13.653
R14392 vp_p.n3305 vp_p.n3304 13.653
R14393 vp_p.n3307 vp_p.n3306 13.653
R14394 vp_p.n4729 vp_p.n4728 13.653
R14395 vp_p.n4731 vp_p.n4730 13.653
R14396 vp_p.n6152 vp_p.n6151 13.653
R14397 vp_p.n6154 vp_p.n6153 13.653
R14398 vp_p.n7569 vp_p.n7568 13.653
R14399 vp_p.n7571 vp_p.n7570 13.653
R14400 vp_p.n452 vp_p.n451 1.165
R14401 vp_p.n9191 vp_p.n9190 1.165
R14402 vp_p.n451 vp_p.n450 1.043
R14403 vp_p.n450 vp_p.n449 1.043
R14404 vp_p.n449 vp_p.n448 1.043
R14405 vp_p.n448 vp_p.n447 1.043
R14406 vp_p.n447 vp_p.n446 1.043
R14407 vp_p.n446 vp_p.n445 1.043
R14408 vp_p.n445 vp_p.n444 1.043
R14409 vp_p.n444 vp_p.n443 1.043
R14410 vp_p.n443 vp_p.n442 1.043
R14411 vp_p.n442 vp_p.n441 1.043
R14412 vp_p.n441 vp_p.n440 1.043
R14413 vp_p.n440 vp_p.n439 1.043
R14414 vp_p.n439 vp_p.n438 1.043
R14415 vp_p.n438 vp_p.n437 1.043
R14416 vp_p.n437 vp_p.n436 1.043
R14417 vp_p.n436 vp_p.n435 1.043
R14418 vp_p.n435 vp_p.n434 1.043
R14419 vp_p.n434 vp_p.n433 1.043
R14420 vp_p.n433 vp_p.n432 1.043
R14421 vp_p.n432 vp_p.n431 1.043
R14422 vp_p.n431 vp_p.n430 1.043
R14423 vp_p.n430 vp_p.n429 1.043
R14424 vp_p.n429 vp_p.n428 1.043
R14425 vp_p.n428 vp_p.n427 1.043
R14426 vp_p.n427 vp_p.n426 1.043
R14427 vp_p.n426 vp_p.n425 1.043
R14428 vp_p.n425 vp_p.n424 1.043
R14429 vp_p.n424 vp_p.n423 1.043
R14430 vp_p.n423 vp_p.n422 1.043
R14431 vp_p.n422 vp_p.n421 1.043
R14432 vp_p.n421 vp_p.n420 1.043
R14433 vp_p.n420 vp_p.n419 1.043
R14434 vp_p.n419 vp_p.n418 1.043
R14435 vp_p.n418 vp_p.n417 1.043
R14436 vp_p.n417 vp_p.n416 1.043
R14437 vp_p.n416 vp_p.n415 1.043
R14438 vp_p.n415 vp_p.n414 1.043
R14439 vp_p.n414 vp_p.n413 1.043
R14440 vp_p.n413 vp_p.n412 1.043
R14441 vp_p.n412 vp_p.n411 1.043
R14442 vp_p.n411 vp_p.n410 1.043
R14443 vp_p.n410 vp_p.n409 1.043
R14444 vp_p.n409 vp_p.n408 1.043
R14445 vp_p.n408 vp_p.n407 1.043
R14446 vp_p.n407 vp_p.n406 1.043
R14447 vp_p.n406 vp_p.n405 1.043
R14448 vp_p.n405 vp_p.n404 1.043
R14449 vp_p.n404 vp_p.n403 1.043
R14450 vp_p.n403 vp_p.n402 1.043
R14451 vp_p.n402 vp_p.n401 1.043
R14452 vp_p.n401 vp_p.n400 1.043
R14453 vp_p.n8631 vp_p.n8630 1.043
R14454 vp_p.n8632 vp_p.n8631 1.043
R14455 vp_p.n8633 vp_p.n8632 1.043
R14456 vp_p.n8634 vp_p.n8633 1.043
R14457 vp_p.n8635 vp_p.n8634 1.043
R14458 vp_p.n8636 vp_p.n8635 1.043
R14459 vp_p.n8637 vp_p.n8636 1.043
R14460 vp_p.n8638 vp_p.n8637 1.043
R14461 vp_p.n8639 vp_p.n8638 1.043
R14462 vp_p.n8640 vp_p.n8639 1.043
R14463 vp_p.n8641 vp_p.n8640 1.043
R14464 vp_p.n8642 vp_p.n8641 1.043
R14465 vp_p.n8643 vp_p.n8642 1.043
R14466 vp_p.n8644 vp_p.n8643 1.043
R14467 vp_p.n8645 vp_p.n8644 1.043
R14468 vp_p.n8646 vp_p.n8645 1.043
R14469 vp_p.n8647 vp_p.n8646 1.043
R14470 vp_p.n8648 vp_p.n8647 1.043
R14471 vp_p.n8649 vp_p.n8648 1.043
R14472 vp_p.n8650 vp_p.n8649 1.043
R14473 vp_p.n8651 vp_p.n8650 1.043
R14474 vp_p.n8652 vp_p.n8651 1.043
R14475 vp_p.n8653 vp_p.n8652 1.043
R14476 vp_p.n8654 vp_p.n8653 1.043
R14477 vp_p.n8655 vp_p.n8654 1.043
R14478 vp_p.n8656 vp_p.n8655 1.043
R14479 vp_p.n8657 vp_p.n8656 1.043
R14480 vp_p.n8658 vp_p.n8657 1.043
R14481 vp_p.n8659 vp_p.n8658 1.043
R14482 vp_p.n8660 vp_p.n8659 1.043
R14483 vp_p.n8661 vp_p.n8660 1.043
R14484 vp_p.n8662 vp_p.n8661 1.043
R14485 vp_p.n8663 vp_p.n8662 1.043
R14486 vp_p.n8664 vp_p.n8663 1.043
R14487 vp_p.n8665 vp_p.n8664 1.043
R14488 vp_p.n8666 vp_p.n8665 1.043
R14489 vp_p.n8667 vp_p.n8666 1.043
R14490 vp_p.n8668 vp_p.n8667 1.043
R14491 vp_p.n8669 vp_p.n8668 1.043
R14492 vp_p.n8670 vp_p.n8669 1.043
R14493 vp_p.n8671 vp_p.n8670 1.043
R14494 vp_p.n8672 vp_p.n8671 1.043
R14495 vp_p.n8673 vp_p.n8672 1.043
R14496 vp_p.n8674 vp_p.n8673 1.043
R14497 vp_p.n8675 vp_p.n8674 1.043
R14498 vp_p.n8676 vp_p.n8675 1.043
R14499 vp_p.n8677 vp_p.n8676 1.043
R14500 vp_p.n8678 vp_p.n8677 1.043
R14501 vp_p.n8679 vp_p.n8678 1.043
R14502 vp_p.n8680 vp_p.n8679 1.043
R14503 vp_p.n8681 vp_p.n8680 1.043
R14504 vp_p.n8682 vp_p.n8681 1.043
R14505 vp_p.n8683 vp_p.n8682 1.043
R14506 vp_p.n8684 vp_p.n8683 1.043
R14507 vp_p.n8685 vp_p.n8684 1.043
R14508 vp_p.n8686 vp_p.n8685 1.043
R14509 vp_p.n8687 vp_p.n8686 1.043
R14510 vp_p.n8688 vp_p.n8687 1.043
R14511 vp_p.n8689 vp_p.n8688 1.043
R14512 vp_p.n8690 vp_p.n8689 1.043
R14513 vp_p.n8691 vp_p.n8690 1.043
R14514 vp_p.n8692 vp_p.n8691 1.043
R14515 vp_p.n8693 vp_p.n8692 1.043
R14516 vp_p.n8694 vp_p.n8693 1.043
R14517 vp_p.n8695 vp_p.n8694 1.043
R14518 vp_p.n8696 vp_p.n8695 1.043
R14519 vp_p.n8697 vp_p.n8696 1.043
R14520 vp_p.n8698 vp_p.n8697 1.043
R14521 vp_p.n8699 vp_p.n8698 1.043
R14522 vp_p.n8700 vp_p.n8699 1.043
R14523 vp_p.n8701 vp_p.n8700 1.043
R14524 vp_p.n8702 vp_p.n8701 1.043
R14525 vp_p.n8703 vp_p.n8702 1.043
R14526 vp_p.n8704 vp_p.n8703 1.043
R14527 vp_p.n8705 vp_p.n8704 1.043
R14528 vp_p.n8706 vp_p.n8705 1.043
R14529 vp_p.n8707 vp_p.n8706 1.043
R14530 vp_p.n8708 vp_p.n8707 1.043
R14531 vp_p.n8709 vp_p.n8708 1.043
R14532 vp_p.n8710 vp_p.n8709 1.043
R14533 vp_p.n8711 vp_p.n8710 1.043
R14534 vp_p.n8712 vp_p.n8711 1.043
R14535 vp_p.n8713 vp_p.n8712 1.043
R14536 vp_p.n8714 vp_p.n8713 1.043
R14537 vp_p.n8715 vp_p.n8714 1.043
R14538 vp_p.n8716 vp_p.n8715 1.043
R14539 vp_p.n8717 vp_p.n8716 1.043
R14540 vp_p.n8718 vp_p.n8717 1.043
R14541 vp_p.n8719 vp_p.n8718 1.043
R14542 vp_p.n8720 vp_p.n8719 1.043
R14543 vp_p.n8721 vp_p.n8720 1.043
R14544 vp_p.n8722 vp_p.n8721 1.043
R14545 vp_p.n8723 vp_p.n8722 1.043
R14546 vp_p.n8724 vp_p.n8723 1.043
R14547 vp_p.n8725 vp_p.n8724 1.043
R14548 vp_p.n8726 vp_p.n8725 1.043
R14549 vp_p.n8727 vp_p.n8726 1.043
R14550 vp_p.n9190 vp_p.n9189 1.043
R14551 vp_p.n9189 vp_p.n9188 1.043
R14552 vp_p.n9188 vp_p.n9187 1.043
R14553 vp_p.n9187 vp_p.n9186 1.043
R14554 vp_p.n9186 vp_p.n9185 1.043
R14555 vp_p.n9185 vp_p.n9184 1.043
R14556 vp_p.n9184 vp_p.n9183 1.043
R14557 vp_p.n9183 vp_p.n9182 1.043
R14558 vp_p.n9182 vp_p.n9181 1.043
R14559 vp_p.n9181 vp_p.n9180 1.043
R14560 vp_p.n9180 vp_p.n9179 1.043
R14561 vp_p.n9179 vp_p.n9178 1.043
R14562 vp_p.n9178 vp_p.n9177 1.043
R14563 vp_p.n9177 vp_p.n9176 1.043
R14564 vp_p.n9176 vp_p.n9175 1.043
R14565 vp_p.n9175 vp_p.n9174 1.043
R14566 vp_p.n9174 vp_p.n9173 1.043
R14567 vp_p.n9173 vp_p.n9172 1.043
R14568 vp_p.n9172 vp_p.n9171 1.043
R14569 vp_p.n9171 vp_p.n9170 1.043
R14570 vp_p.n9170 vp_p.n9169 1.043
R14571 vp_p.n9169 vp_p.n9168 1.043
R14572 vp_p.n9168 vp_p.n9167 1.043
R14573 vp_p.n9167 vp_p.n9166 1.043
R14574 vp_p.n9166 vp_p.n9165 1.043
R14575 vp_p.n9165 vp_p.n9164 1.043
R14576 vp_p.n9164 vp_p.n9163 1.043
R14577 vp_p.n9163 vp_p.n9162 1.043
R14578 vp_p.n9162 vp_p.n9161 1.043
R14579 vp_p.n9161 vp_p.n9160 1.043
R14580 vp_p.n9160 vp_p.n9159 1.043
R14581 vp_p.n9159 vp_p.n9158 1.043
R14582 vp_p.n9158 vp_p.n9157 1.043
R14583 vp_p.n9157 vp_p.n9156 1.043
R14584 vp_p.n9156 vp_p.n9155 1.043
R14585 vp_p.n9155 vp_p.n9154 1.043
R14586 vp_p.n9154 vp_p.n9153 1.043
R14587 vp_p.n9153 vp_p.n9152 1.043
R14588 vp_p.n9152 vp_p.n9151 1.043
R14589 vp_p.n9151 vp_p.n9150 1.043
R14590 vp_p.n9150 vp_p.n9149 1.043
R14591 vp_p.n9149 vp_p.n9148 1.043
R14592 vp_p.n9148 vp_p.n9147 1.043
R14593 vp_p.n9147 vp_p.n9146 1.043
R14594 vp_p.n9146 vp_p.n9145 1.043
R14595 vp_p.n9145 vp_p.n9144 1.043
R14596 vp_p.n9144 vp_p.n9143 1.043
R14597 vp_p.n9143 vp_p.n9142 1.043
R14598 vp_p.n9142 vp_p.n9141 1.043
R14599 vp_p.n9141 vp_p.n9140 1.043
R14600 vp_p.n9140 vp_p.n9139 1.043
R14601 vp_p.n27329 vp_p.n27328 1.043
R14602 vp_p.n27330 vp_p.n27329 1.043
R14603 vp_p.n27331 vp_p.n27330 1.043
R14604 vp_p.n27332 vp_p.n27331 1.043
R14605 vp_p.n27333 vp_p.n27332 1.043
R14606 vp_p.n27334 vp_p.n27333 1.043
R14607 vp_p.n27335 vp_p.n27334 1.043
R14608 vp_p.n27336 vp_p.n27335 1.043
R14609 vp_p.n27337 vp_p.n27336 1.043
R14610 vp_p.n27338 vp_p.n27337 1.043
R14611 vp_p.n27339 vp_p.n27338 1.043
R14612 vp_p.n27340 vp_p.n27339 1.043
R14613 vp_p.n27341 vp_p.n27340 1.043
R14614 vp_p.n27342 vp_p.n27341 1.043
R14615 vp_p.n27343 vp_p.n27342 1.043
R14616 vp_p.n27344 vp_p.n27343 1.043
R14617 vp_p.n27345 vp_p.n27344 1.043
R14618 vp_p.n27346 vp_p.n27345 1.043
R14619 vp_p.n27347 vp_p.n27346 1.043
R14620 vp_p.n27348 vp_p.n27347 1.043
R14621 vp_p.n27349 vp_p.n27348 1.043
R14622 vp_p.n27350 vp_p.n27349 1.043
R14623 vp_p.n27351 vp_p.n27350 1.043
R14624 vp_p.n27352 vp_p.n27351 1.043
R14625 vp_p.n27353 vp_p.n27352 1.043
R14626 vp_p.n27354 vp_p.n27353 1.043
R14627 vp_p.n27355 vp_p.n27354 1.043
R14628 vp_p.n27356 vp_p.n27355 1.043
R14629 vp_p.n27357 vp_p.n27356 1.043
R14630 vp_p.n27358 vp_p.n27357 1.043
R14631 vp_p.n27359 vp_p.n27358 1.043
R14632 vp_p.n27360 vp_p.n27359 1.043
R14633 vp_p.n27361 vp_p.n27360 1.043
R14634 vp_p.n27362 vp_p.n27361 1.043
R14635 vp_p.n27363 vp_p.n27362 1.043
R14636 vp_p.n27364 vp_p.n27363 1.043
R14637 vp_p.n27365 vp_p.n27364 1.043
R14638 vp_p.n27366 vp_p.n27365 1.043
R14639 vp_p.n27367 vp_p.n27366 1.043
R14640 vp_p.n27368 vp_p.n27367 1.043
R14641 vp_p.n27369 vp_p.n27368 1.043
R14642 vp_p.n27370 vp_p.n27369 1.043
R14643 vp_p.n27371 vp_p.n27370 1.043
R14644 vp_p.n27372 vp_p.n27371 1.043
R14645 vp_p.n27373 vp_p.n27372 1.043
R14646 vp_p.n27374 vp_p.n27373 1.043
R14647 vp_p.n27375 vp_p.n27374 1.043
R14648 vp_p.n27376 vp_p.n27375 1.043
R14649 vp_p.n27377 vp_p.n27376 1.043
R14650 vp_p.n27378 vp_p.n27377 1.043
R14651 vp_p.n27379 vp_p.n27378 1.043
R14652 vp_p.n27380 vp_p.n27379 1.043
R14653 vp_p.n27381 vp_p.n27380 1.043
R14654 vp_p.n27382 vp_p.n27381 1.043
R14655 vp_p.n27383 vp_p.n27382 1.043
R14656 vp_p.n27384 vp_p.n27383 1.043
R14657 vp_p.n27385 vp_p.n27384 1.043
R14658 vp_p.n27386 vp_p.n27385 1.043
R14659 vp_p.n27387 vp_p.n27386 1.043
R14660 vp_p.n27388 vp_p.n27387 1.043
R14661 vp_p.n27389 vp_p.n27388 1.043
R14662 vp_p.n27390 vp_p.n27389 1.043
R14663 vp_p.n27391 vp_p.n27390 1.043
R14664 vp_p.n27392 vp_p.n27391 1.043
R14665 vp_p.n27393 vp_p.n27392 1.043
R14666 vp_p.n27394 vp_p.n27393 1.043
R14667 vp_p.n27395 vp_p.n27394 1.043
R14668 vp_p.n27396 vp_p.n27395 1.043
R14669 vp_p.n27397 vp_p.n27396 1.043
R14670 vp_p.n27398 vp_p.n27397 1.043
R14671 vp_p.n27399 vp_p.n27398 1.043
R14672 vp_p.n27400 vp_p.n27399 1.043
R14673 vp_p.n27401 vp_p.n27400 1.043
R14674 vp_p.n27402 vp_p.n27401 1.043
R14675 vp_p.n27403 vp_p.n27402 1.043
R14676 vp_p.n27404 vp_p.n27403 1.043
R14677 vp_p.n27405 vp_p.n27404 1.043
R14678 vp_p.n27406 vp_p.n27405 1.043
R14679 vp_p.n27407 vp_p.n27406 1.043
R14680 vp_p.n27408 vp_p.n27407 1.043
R14681 vp_p.n27409 vp_p.n27408 1.043
R14682 vp_p.n27410 vp_p.n27409 1.043
R14683 vp_p.n27411 vp_p.n27410 1.043
R14684 vp_p.n27412 vp_p.n27411 1.043
R14685 vp_p.n27413 vp_p.n27412 1.043
R14686 vp_p.n27414 vp_p.n27413 1.043
R14687 vp_p.n27415 vp_p.n27414 1.043
R14688 vp_p.n27416 vp_p.n27415 1.043
R14689 vp_p.n27417 vp_p.n27416 1.043
R14690 vp_p.n27418 vp_p.n27417 1.043
R14691 vp_p.n27419 vp_p.n27418 1.043
R14692 vp_p.n27420 vp_p.n27419 1.043
R14693 vp_p.n27421 vp_p.n27420 1.043
R14694 vp_p.n27422 vp_p.n27421 1.043
R14695 vp_p.n27423 vp_p.n27422 1.043
R14696 vp_p.n27424 vp_p.n27423 1.043
R14697 vp_p.n27425 vp_p.n27424 1.043
R14698 vp_p.n8728 vp_p.n8727 0.979
R14699 vp_p.n27426 vp_p.n27425 0.979
R14700 vp_p.n13848 vp_p.n13847 0.296
R14701 vp_p.n13853 vp_p.n13852 0.296
R14702 vp_p.n13857 vp_p.n13856 0.296
R14703 vp_p.n13861 vp_p.n13860 0.296
R14704 vp_p.n13865 vp_p.n13864 0.296
R14705 vp_p.n13869 vp_p.n13868 0.296
R14706 vp_p.n13873 vp_p.n13872 0.296
R14707 vp_p.n13877 vp_p.n13876 0.296
R14708 vp_p.n13881 vp_p.n13880 0.296
R14709 vp_p.n13885 vp_p.n13884 0.296
R14710 vp_p.n13889 vp_p.n13888 0.296
R14711 vp_p.n13893 vp_p.n13892 0.296
R14712 vp_p.n13897 vp_p.n13896 0.296
R14713 vp_p.n13901 vp_p.n13900 0.296
R14714 vp_p.n13905 vp_p.n13904 0.296
R14715 vp_p.n13909 vp_p.n13908 0.296
R14716 vp_p.n13913 vp_p.n13912 0.296
R14717 vp_p.n13917 vp_p.n13916 0.296
R14718 vp_p.n13921 vp_p.n13920 0.296
R14719 vp_p.n13925 vp_p.n13924 0.296
R14720 vp_p.n13929 vp_p.n13928 0.296
R14721 vp_p.n13933 vp_p.n13932 0.296
R14722 vp_p.n13937 vp_p.n13936 0.296
R14723 vp_p.n13941 vp_p.n13940 0.296
R14724 vp_p.n13945 vp_p.n13944 0.296
R14725 vp_p.n13949 vp_p.n13948 0.296
R14726 vp_p.n13953 vp_p.n13952 0.296
R14727 vp_p.n13957 vp_p.n13956 0.296
R14728 vp_p.n13961 vp_p.n13960 0.296
R14729 vp_p.n13965 vp_p.n13964 0.296
R14730 vp_p.n13969 vp_p.n13968 0.296
R14731 vp_p.n13973 vp_p.n13972 0.296
R14732 vp_p.n13977 vp_p.n13976 0.296
R14733 vp_p.n13981 vp_p.n13980 0.296
R14734 vp_p.n13985 vp_p.n13984 0.296
R14735 vp_p.n13989 vp_p.n13988 0.296
R14736 vp_p.n13993 vp_p.n13992 0.296
R14737 vp_p.n13997 vp_p.n13996 0.296
R14738 vp_p.n14001 vp_p.n14000 0.296
R14739 vp_p.n14005 vp_p.n14004 0.296
R14740 vp_p.n14009 vp_p.n14008 0.296
R14741 vp_p.n14013 vp_p.n14012 0.296
R14742 vp_p.n14017 vp_p.n14016 0.296
R14743 vp_p.n14021 vp_p.n14020 0.296
R14744 vp_p.n14025 vp_p.n14024 0.296
R14745 vp_p.n14029 vp_p.n14028 0.296
R14746 vp_p.n14033 vp_p.n14032 0.296
R14747 vp_p.n14037 vp_p.n14036 0.296
R14748 vp_p.n14041 vp_p.n14040 0.296
R14749 vp_p.n14045 vp_p.n14044 0.296
R14750 vp_p.n14049 vp_p.n14048 0.296
R14751 vp_p.n14053 vp_p.n14052 0.296
R14752 vp_p.n14057 vp_p.n14056 0.296
R14753 vp_p.n14061 vp_p.n14060 0.296
R14754 vp_p.n14065 vp_p.n14064 0.296
R14755 vp_p.n14069 vp_p.n14068 0.296
R14756 vp_p.n14073 vp_p.n14072 0.296
R14757 vp_p.n14077 vp_p.n14076 0.296
R14758 vp_p.n14081 vp_p.n14080 0.296
R14759 vp_p.n14085 vp_p.n14084 0.296
R14760 vp_p.n14089 vp_p.n14088 0.296
R14761 vp_p.n14093 vp_p.n14092 0.296
R14762 vp_p.n14097 vp_p.n14096 0.296
R14763 vp_p.n14101 vp_p.n14100 0.296
R14764 vp_p.n14105 vp_p.n14104 0.296
R14765 vp_p.n14109 vp_p.n14108 0.296
R14766 vp_p.n14113 vp_p.n14112 0.296
R14767 vp_p.n14117 vp_p.n14116 0.296
R14768 vp_p.n14121 vp_p.n14120 0.296
R14769 vp_p.n14125 vp_p.n14124 0.296
R14770 vp_p.n14129 vp_p.n14128 0.296
R14771 vp_p.n14133 vp_p.n14132 0.296
R14772 vp_p.n14137 vp_p.n14136 0.296
R14773 vp_p.n14141 vp_p.n14140 0.296
R14774 vp_p.n14145 vp_p.n14144 0.296
R14775 vp_p.n14149 vp_p.n14148 0.296
R14776 vp_p.n14153 vp_p.n14152 0.296
R14777 vp_p.n14157 vp_p.n14156 0.296
R14778 vp_p.n14161 vp_p.n14160 0.296
R14779 vp_p.n14165 vp_p.n14164 0.296
R14780 vp_p.n14169 vp_p.n14168 0.296
R14781 vp_p.n14173 vp_p.n14172 0.296
R14782 vp_p.n14177 vp_p.n14176 0.296
R14783 vp_p.n14181 vp_p.n14180 0.296
R14784 vp_p.n14185 vp_p.n14184 0.296
R14785 vp_p.n14189 vp_p.n14188 0.296
R14786 vp_p.n14193 vp_p.n14192 0.296
R14787 vp_p.n14197 vp_p.n14196 0.296
R14788 vp_p.n14201 vp_p.n14200 0.296
R14789 vp_p.n14205 vp_p.n14204 0.296
R14790 vp_p.n14209 vp_p.n14208 0.296
R14791 vp_p.n14213 vp_p.n14212 0.296
R14792 vp_p.n14217 vp_p.n14216 0.296
R14793 vp_p.n14221 vp_p.n14220 0.296
R14794 vp_p.n14225 vp_p.n14224 0.296
R14795 vp_p.n14229 vp_p.n14228 0.296
R14796 vp_p.n14233 vp_p.n14232 0.296
R14797 vp_p.n14237 vp_p.n14236 0.296
R14798 vp_p.n14241 vp_p.n14240 0.296
R14799 vp_p.n14245 vp_p.n14244 0.296
R14800 vp_p.n14249 vp_p.n14248 0.296
R14801 vp_p.n14253 vp_p.n14252 0.296
R14802 vp_p.n14257 vp_p.n14256 0.296
R14803 vp_p.n14261 vp_p.n14260 0.296
R14804 vp_p.n14265 vp_p.n14264 0.296
R14805 vp_p.n14269 vp_p.n14268 0.296
R14806 vp_p.n14273 vp_p.n14272 0.296
R14807 vp_p.n14277 vp_p.n14276 0.296
R14808 vp_p.n14281 vp_p.n14280 0.296
R14809 vp_p.n14285 vp_p.n14284 0.296
R14810 vp_p.n14289 vp_p.n14288 0.296
R14811 vp_p.n14293 vp_p.n14292 0.296
R14812 vp_p.n14297 vp_p.n14296 0.296
R14813 vp_p.n14301 vp_p.n14300 0.296
R14814 vp_p.n14305 vp_p.n14304 0.296
R14815 vp_p.n14309 vp_p.n14308 0.296
R14816 vp_p.n14313 vp_p.n14312 0.296
R14817 vp_p.n14317 vp_p.n14316 0.296
R14818 vp_p.n14321 vp_p.n14320 0.296
R14819 vp_p.n14325 vp_p.n14324 0.296
R14820 vp_p.n14329 vp_p.n14328 0.296
R14821 vp_p.n14333 vp_p.n14332 0.296
R14822 vp_p.n14337 vp_p.n14336 0.296
R14823 vp_p.n14341 vp_p.n14340 0.296
R14824 vp_p.n14345 vp_p.n14344 0.296
R14825 vp_p.n14349 vp_p.n14348 0.296
R14826 vp_p.n14353 vp_p.n14352 0.296
R14827 vp_p.n14357 vp_p.n14356 0.296
R14828 vp_p.n14361 vp_p.n14360 0.296
R14829 vp_p.n14365 vp_p.n14364 0.296
R14830 vp_p.n14369 vp_p.n14368 0.296
R14831 vp_p.n14373 vp_p.n14372 0.296
R14832 vp_p.n14377 vp_p.n14376 0.296
R14833 vp_p.n14387 vp_p.n14386 0.296
R14834 vp_p.n14392 vp_p.n14391 0.296
R14835 vp_p.n14397 vp_p.n14396 0.296
R14836 vp_p.n14402 vp_p.n14401 0.296
R14837 vp_p.n14407 vp_p.n14406 0.296
R14838 vp_p.n14412 vp_p.n14411 0.296
R14839 vp_p.n14417 vp_p.n14416 0.296
R14840 vp_p.n14422 vp_p.n14421 0.296
R14841 vp_p.n14427 vp_p.n14426 0.296
R14842 vp_p.n14432 vp_p.n14431 0.296
R14843 vp_p.n14437 vp_p.n14436 0.296
R14844 vp_p.n14442 vp_p.n14441 0.296
R14845 vp_p.n14447 vp_p.n14446 0.296
R14846 vp_p.n14452 vp_p.n14451 0.296
R14847 vp_p.n14457 vp_p.n14456 0.296
R14848 vp_p.n14462 vp_p.n14461 0.296
R14849 vp_p.n12084 vp_p.n12083 0.296
R14850 vp_p.n12089 vp_p.n12088 0.296
R14851 vp_p.n12099 vp_p.n12098 0.296
R14852 vp_p.n12103 vp_p.n12102 0.296
R14853 vp_p.n12113 vp_p.n12112 0.296
R14854 vp_p.n12117 vp_p.n12116 0.296
R14855 vp_p.n12127 vp_p.n12126 0.296
R14856 vp_p.n12131 vp_p.n12130 0.296
R14857 vp_p.n12141 vp_p.n12140 0.296
R14858 vp_p.n12145 vp_p.n12144 0.296
R14859 vp_p.n12155 vp_p.n12154 0.296
R14860 vp_p.n12159 vp_p.n12158 0.296
R14861 vp_p.n12169 vp_p.n12168 0.296
R14862 vp_p.n12173 vp_p.n12172 0.296
R14863 vp_p.n12183 vp_p.n12182 0.296
R14864 vp_p.n12187 vp_p.n12186 0.296
R14865 vp_p.n12197 vp_p.n12196 0.296
R14866 vp_p.n12201 vp_p.n12200 0.296
R14867 vp_p.n12211 vp_p.n12210 0.296
R14868 vp_p.n12215 vp_p.n12214 0.296
R14869 vp_p.n12225 vp_p.n12224 0.296
R14870 vp_p.n12229 vp_p.n12228 0.296
R14871 vp_p.n12239 vp_p.n12238 0.296
R14872 vp_p.n12243 vp_p.n12242 0.296
R14873 vp_p.n12253 vp_p.n12252 0.296
R14874 vp_p.n12257 vp_p.n12256 0.296
R14875 vp_p.n12267 vp_p.n12266 0.296
R14876 vp_p.n12271 vp_p.n12270 0.296
R14877 vp_p.n12281 vp_p.n12280 0.296
R14878 vp_p.n12285 vp_p.n12284 0.296
R14879 vp_p.n12295 vp_p.n12294 0.296
R14880 vp_p.n12299 vp_p.n12298 0.296
R14881 vp_p.n12309 vp_p.n12308 0.296
R14882 vp_p.n12313 vp_p.n12312 0.296
R14883 vp_p.n12323 vp_p.n12322 0.296
R14884 vp_p.n12327 vp_p.n12326 0.296
R14885 vp_p.n12337 vp_p.n12336 0.296
R14886 vp_p.n12341 vp_p.n12340 0.296
R14887 vp_p.n12351 vp_p.n12350 0.296
R14888 vp_p.n12355 vp_p.n12354 0.296
R14889 vp_p.n12365 vp_p.n12364 0.296
R14890 vp_p.n12369 vp_p.n12368 0.296
R14891 vp_p.n12379 vp_p.n12378 0.296
R14892 vp_p.n12383 vp_p.n12382 0.296
R14893 vp_p.n12393 vp_p.n12392 0.296
R14894 vp_p.n12397 vp_p.n12396 0.296
R14895 vp_p.n12407 vp_p.n12406 0.296
R14896 vp_p.n12411 vp_p.n12410 0.296
R14897 vp_p.n12421 vp_p.n12420 0.296
R14898 vp_p.n12425 vp_p.n12424 0.296
R14899 vp_p.n12435 vp_p.n12434 0.296
R14900 vp_p.n12439 vp_p.n12438 0.296
R14901 vp_p.n12449 vp_p.n12448 0.296
R14902 vp_p.n12453 vp_p.n12452 0.296
R14903 vp_p.n12463 vp_p.n12462 0.296
R14904 vp_p.n12467 vp_p.n12466 0.296
R14905 vp_p.n12477 vp_p.n12476 0.296
R14906 vp_p.n12481 vp_p.n12480 0.296
R14907 vp_p.n12491 vp_p.n12490 0.296
R14908 vp_p.n12495 vp_p.n12494 0.296
R14909 vp_p.n12505 vp_p.n12504 0.296
R14910 vp_p.n12509 vp_p.n12508 0.296
R14911 vp_p.n12519 vp_p.n12518 0.296
R14912 vp_p.n12523 vp_p.n12522 0.296
R14913 vp_p.n12533 vp_p.n12532 0.296
R14914 vp_p.n12537 vp_p.n12536 0.296
R14915 vp_p.n12547 vp_p.n12546 0.296
R14916 vp_p.n12551 vp_p.n12550 0.296
R14917 vp_p.n12561 vp_p.n12560 0.296
R14918 vp_p.n12565 vp_p.n12564 0.296
R14919 vp_p.n12575 vp_p.n12574 0.296
R14920 vp_p.n12579 vp_p.n12578 0.296
R14921 vp_p.n12589 vp_p.n12588 0.296
R14922 vp_p.n12593 vp_p.n12592 0.296
R14923 vp_p.n12603 vp_p.n12602 0.296
R14924 vp_p.n12607 vp_p.n12606 0.296
R14925 vp_p.n12617 vp_p.n12616 0.296
R14926 vp_p.n12621 vp_p.n12620 0.296
R14927 vp_p.n12631 vp_p.n12630 0.296
R14928 vp_p.n12635 vp_p.n12634 0.296
R14929 vp_p.n12645 vp_p.n12644 0.296
R14930 vp_p.n12649 vp_p.n12648 0.296
R14931 vp_p.n12659 vp_p.n12658 0.296
R14932 vp_p.n12663 vp_p.n12662 0.296
R14933 vp_p.n12673 vp_p.n12672 0.296
R14934 vp_p.n12677 vp_p.n12676 0.296
R14935 vp_p.n12687 vp_p.n12686 0.296
R14936 vp_p.n12691 vp_p.n12690 0.296
R14937 vp_p.n12701 vp_p.n12700 0.296
R14938 vp_p.n12705 vp_p.n12704 0.296
R14939 vp_p.n12715 vp_p.n12714 0.296
R14940 vp_p.n12719 vp_p.n12718 0.296
R14941 vp_p.n12729 vp_p.n12728 0.296
R14942 vp_p.n12733 vp_p.n12732 0.296
R14943 vp_p.n12743 vp_p.n12742 0.296
R14944 vp_p.n12747 vp_p.n12746 0.296
R14945 vp_p.n12757 vp_p.n12756 0.296
R14946 vp_p.n12761 vp_p.n12760 0.296
R14947 vp_p.n12771 vp_p.n12770 0.296
R14948 vp_p.n12775 vp_p.n12774 0.296
R14949 vp_p.n12785 vp_p.n12784 0.296
R14950 vp_p.n12789 vp_p.n12788 0.296
R14951 vp_p.n12799 vp_p.n12798 0.296
R14952 vp_p.n12803 vp_p.n12802 0.296
R14953 vp_p.n12813 vp_p.n12812 0.296
R14954 vp_p.n12817 vp_p.n12816 0.296
R14955 vp_p.n12827 vp_p.n12826 0.296
R14956 vp_p.n12831 vp_p.n12830 0.296
R14957 vp_p.n12841 vp_p.n12840 0.296
R14958 vp_p.n12845 vp_p.n12844 0.296
R14959 vp_p.n12855 vp_p.n12854 0.296
R14960 vp_p.n12859 vp_p.n12858 0.296
R14961 vp_p.n12869 vp_p.n12868 0.296
R14962 vp_p.n12873 vp_p.n12872 0.296
R14963 vp_p.n12883 vp_p.n12882 0.296
R14964 vp_p.n12887 vp_p.n12886 0.296
R14965 vp_p.n12897 vp_p.n12896 0.296
R14966 vp_p.n12901 vp_p.n12900 0.296
R14967 vp_p.n12911 vp_p.n12910 0.296
R14968 vp_p.n12915 vp_p.n12914 0.296
R14969 vp_p.n12925 vp_p.n12924 0.296
R14970 vp_p.n12929 vp_p.n12928 0.296
R14971 vp_p.n12939 vp_p.n12938 0.296
R14972 vp_p.n12943 vp_p.n12942 0.296
R14973 vp_p.n12953 vp_p.n12952 0.296
R14974 vp_p.n12957 vp_p.n12956 0.296
R14975 vp_p.n12967 vp_p.n12966 0.296
R14976 vp_p.n12971 vp_p.n12970 0.296
R14977 vp_p.n12981 vp_p.n12980 0.296
R14978 vp_p.n12985 vp_p.n12984 0.296
R14979 vp_p.n12995 vp_p.n12994 0.296
R14980 vp_p.n12999 vp_p.n12998 0.296
R14981 vp_p.n13009 vp_p.n13008 0.296
R14982 vp_p.n13013 vp_p.n13012 0.296
R14983 vp_p.n13023 vp_p.n13022 0.296
R14984 vp_p.n13028 vp_p.n13027 0.296
R14985 vp_p.n13033 vp_p.n13032 0.296
R14986 vp_p.n13038 vp_p.n13037 0.296
R14987 vp_p.n13043 vp_p.n13042 0.296
R14988 vp_p.n13048 vp_p.n13047 0.296
R14989 vp_p.n13053 vp_p.n13052 0.296
R14990 vp_p.n13058 vp_p.n13057 0.296
R14991 vp_p.n13063 vp_p.n13062 0.296
R14992 vp_p.n13068 vp_p.n13067 0.296
R14993 vp_p.n13073 vp_p.n13072 0.296
R14994 vp_p.n13078 vp_p.n13077 0.296
R14995 vp_p.n13083 vp_p.n13082 0.296
R14996 vp_p.n13088 vp_p.n13087 0.296
R14997 vp_p.n13093 vp_p.n13092 0.296
R14998 vp_p.n14887 vp_p.n14886 0.296
R14999 vp_p.n14892 vp_p.n14891 0.296
R15000 vp_p.n14902 vp_p.n14901 0.296
R15001 vp_p.n14906 vp_p.n14905 0.296
R15002 vp_p.n14916 vp_p.n14915 0.296
R15003 vp_p.n14920 vp_p.n14919 0.296
R15004 vp_p.n14930 vp_p.n14929 0.296
R15005 vp_p.n14934 vp_p.n14933 0.296
R15006 vp_p.n14944 vp_p.n14943 0.296
R15007 vp_p.n14948 vp_p.n14947 0.296
R15008 vp_p.n14958 vp_p.n14957 0.296
R15009 vp_p.n14962 vp_p.n14961 0.296
R15010 vp_p.n14972 vp_p.n14971 0.296
R15011 vp_p.n14976 vp_p.n14975 0.296
R15012 vp_p.n14986 vp_p.n14985 0.296
R15013 vp_p.n14990 vp_p.n14989 0.296
R15014 vp_p.n15000 vp_p.n14999 0.296
R15015 vp_p.n15004 vp_p.n15003 0.296
R15016 vp_p.n15014 vp_p.n15013 0.296
R15017 vp_p.n15018 vp_p.n15017 0.296
R15018 vp_p.n15028 vp_p.n15027 0.296
R15019 vp_p.n15032 vp_p.n15031 0.296
R15020 vp_p.n15042 vp_p.n15041 0.296
R15021 vp_p.n15046 vp_p.n15045 0.296
R15022 vp_p.n15056 vp_p.n15055 0.296
R15023 vp_p.n15060 vp_p.n15059 0.296
R15024 vp_p.n15070 vp_p.n15069 0.296
R15025 vp_p.n15074 vp_p.n15073 0.296
R15026 vp_p.n15084 vp_p.n15083 0.296
R15027 vp_p.n15088 vp_p.n15087 0.296
R15028 vp_p.n15098 vp_p.n15097 0.296
R15029 vp_p.n15102 vp_p.n15101 0.296
R15030 vp_p.n15112 vp_p.n15111 0.296
R15031 vp_p.n15116 vp_p.n15115 0.296
R15032 vp_p.n15126 vp_p.n15125 0.296
R15033 vp_p.n15130 vp_p.n15129 0.296
R15034 vp_p.n15140 vp_p.n15139 0.296
R15035 vp_p.n15144 vp_p.n15143 0.296
R15036 vp_p.n15154 vp_p.n15153 0.296
R15037 vp_p.n15158 vp_p.n15157 0.296
R15038 vp_p.n15168 vp_p.n15167 0.296
R15039 vp_p.n15172 vp_p.n15171 0.296
R15040 vp_p.n15182 vp_p.n15181 0.296
R15041 vp_p.n15186 vp_p.n15185 0.296
R15042 vp_p.n15196 vp_p.n15195 0.296
R15043 vp_p.n15200 vp_p.n15199 0.296
R15044 vp_p.n15210 vp_p.n15209 0.296
R15045 vp_p.n15214 vp_p.n15213 0.296
R15046 vp_p.n15224 vp_p.n15223 0.296
R15047 vp_p.n15228 vp_p.n15227 0.296
R15048 vp_p.n15238 vp_p.n15237 0.296
R15049 vp_p.n15242 vp_p.n15241 0.296
R15050 vp_p.n15252 vp_p.n15251 0.296
R15051 vp_p.n15256 vp_p.n15255 0.296
R15052 vp_p.n15266 vp_p.n15265 0.296
R15053 vp_p.n15270 vp_p.n15269 0.296
R15054 vp_p.n15280 vp_p.n15279 0.296
R15055 vp_p.n15284 vp_p.n15283 0.296
R15056 vp_p.n15294 vp_p.n15293 0.296
R15057 vp_p.n15298 vp_p.n15297 0.296
R15058 vp_p.n15308 vp_p.n15307 0.296
R15059 vp_p.n15312 vp_p.n15311 0.296
R15060 vp_p.n15322 vp_p.n15321 0.296
R15061 vp_p.n15326 vp_p.n15325 0.296
R15062 vp_p.n15336 vp_p.n15335 0.296
R15063 vp_p.n15340 vp_p.n15339 0.296
R15064 vp_p.n15350 vp_p.n15349 0.296
R15065 vp_p.n15354 vp_p.n15353 0.296
R15066 vp_p.n15364 vp_p.n15363 0.296
R15067 vp_p.n15368 vp_p.n15367 0.296
R15068 vp_p.n15378 vp_p.n15377 0.296
R15069 vp_p.n15382 vp_p.n15381 0.296
R15070 vp_p.n15392 vp_p.n15391 0.296
R15071 vp_p.n15396 vp_p.n15395 0.296
R15072 vp_p.n15406 vp_p.n15405 0.296
R15073 vp_p.n15410 vp_p.n15409 0.296
R15074 vp_p.n15420 vp_p.n15419 0.296
R15075 vp_p.n15424 vp_p.n15423 0.296
R15076 vp_p.n15434 vp_p.n15433 0.296
R15077 vp_p.n15438 vp_p.n15437 0.296
R15078 vp_p.n15448 vp_p.n15447 0.296
R15079 vp_p.n15452 vp_p.n15451 0.296
R15080 vp_p.n15462 vp_p.n15461 0.296
R15081 vp_p.n15466 vp_p.n15465 0.296
R15082 vp_p.n15476 vp_p.n15475 0.296
R15083 vp_p.n15480 vp_p.n15479 0.296
R15084 vp_p.n15490 vp_p.n15489 0.296
R15085 vp_p.n15494 vp_p.n15493 0.296
R15086 vp_p.n15504 vp_p.n15503 0.296
R15087 vp_p.n15508 vp_p.n15507 0.296
R15088 vp_p.n15518 vp_p.n15517 0.296
R15089 vp_p.n15522 vp_p.n15521 0.296
R15090 vp_p.n15532 vp_p.n15531 0.296
R15091 vp_p.n15536 vp_p.n15535 0.296
R15092 vp_p.n15546 vp_p.n15545 0.296
R15093 vp_p.n15550 vp_p.n15549 0.296
R15094 vp_p.n15560 vp_p.n15559 0.296
R15095 vp_p.n15564 vp_p.n15563 0.296
R15096 vp_p.n15574 vp_p.n15573 0.296
R15097 vp_p.n15578 vp_p.n15577 0.296
R15098 vp_p.n15588 vp_p.n15587 0.296
R15099 vp_p.n15592 vp_p.n15591 0.296
R15100 vp_p.n15602 vp_p.n15601 0.296
R15101 vp_p.n15606 vp_p.n15605 0.296
R15102 vp_p.n15616 vp_p.n15615 0.296
R15103 vp_p.n15620 vp_p.n15619 0.296
R15104 vp_p.n15630 vp_p.n15629 0.296
R15105 vp_p.n15634 vp_p.n15633 0.296
R15106 vp_p.n15644 vp_p.n15643 0.296
R15107 vp_p.n15648 vp_p.n15647 0.296
R15108 vp_p.n15658 vp_p.n15657 0.296
R15109 vp_p.n15662 vp_p.n15661 0.296
R15110 vp_p.n15672 vp_p.n15671 0.296
R15111 vp_p.n15676 vp_p.n15675 0.296
R15112 vp_p.n15686 vp_p.n15685 0.296
R15113 vp_p.n15690 vp_p.n15689 0.296
R15114 vp_p.n15700 vp_p.n15699 0.296
R15115 vp_p.n15704 vp_p.n15703 0.296
R15116 vp_p.n15714 vp_p.n15713 0.296
R15117 vp_p.n15718 vp_p.n15717 0.296
R15118 vp_p.n15728 vp_p.n15727 0.296
R15119 vp_p.n15732 vp_p.n15731 0.296
R15120 vp_p.n15742 vp_p.n15741 0.296
R15121 vp_p.n15746 vp_p.n15745 0.296
R15122 vp_p.n15756 vp_p.n15755 0.296
R15123 vp_p.n15760 vp_p.n15759 0.296
R15124 vp_p.n15770 vp_p.n15769 0.296
R15125 vp_p.n15774 vp_p.n15773 0.296
R15126 vp_p.n15784 vp_p.n15783 0.296
R15127 vp_p.n15788 vp_p.n15787 0.296
R15128 vp_p.n15798 vp_p.n15797 0.296
R15129 vp_p.n15802 vp_p.n15801 0.296
R15130 vp_p.n15812 vp_p.n15811 0.296
R15131 vp_p.n15816 vp_p.n15815 0.296
R15132 vp_p.n15820 vp_p.n15819 0.296
R15133 vp_p.n15830 vp_p.n15829 0.296
R15134 vp_p.n15835 vp_p.n15834 0.296
R15135 vp_p.n15840 vp_p.n15839 0.296
R15136 vp_p.n15845 vp_p.n15844 0.296
R15137 vp_p.n15850 vp_p.n15849 0.296
R15138 vp_p.n15855 vp_p.n15854 0.296
R15139 vp_p.n15860 vp_p.n15859 0.296
R15140 vp_p.n15865 vp_p.n15864 0.296
R15141 vp_p.n15870 vp_p.n15869 0.296
R15142 vp_p.n15875 vp_p.n15874 0.296
R15143 vp_p.n15880 vp_p.n15879 0.296
R15144 vp_p.n15885 vp_p.n15884 0.296
R15145 vp_p.n15890 vp_p.n15889 0.296
R15146 vp_p.n15895 vp_p.n15894 0.296
R15147 vp_p.n10646 vp_p.n10645 0.296
R15148 vp_p.n10651 vp_p.n10650 0.296
R15149 vp_p.n10661 vp_p.n10660 0.296
R15150 vp_p.n10665 vp_p.n10664 0.296
R15151 vp_p.n10675 vp_p.n10674 0.296
R15152 vp_p.n10679 vp_p.n10678 0.296
R15153 vp_p.n10689 vp_p.n10688 0.296
R15154 vp_p.n10693 vp_p.n10692 0.296
R15155 vp_p.n10703 vp_p.n10702 0.296
R15156 vp_p.n10707 vp_p.n10706 0.296
R15157 vp_p.n10717 vp_p.n10716 0.296
R15158 vp_p.n10721 vp_p.n10720 0.296
R15159 vp_p.n10731 vp_p.n10730 0.296
R15160 vp_p.n10735 vp_p.n10734 0.296
R15161 vp_p.n10745 vp_p.n10744 0.296
R15162 vp_p.n10749 vp_p.n10748 0.296
R15163 vp_p.n10759 vp_p.n10758 0.296
R15164 vp_p.n10763 vp_p.n10762 0.296
R15165 vp_p.n10773 vp_p.n10772 0.296
R15166 vp_p.n10777 vp_p.n10776 0.296
R15167 vp_p.n10787 vp_p.n10786 0.296
R15168 vp_p.n10791 vp_p.n10790 0.296
R15169 vp_p.n10801 vp_p.n10800 0.296
R15170 vp_p.n10805 vp_p.n10804 0.296
R15171 vp_p.n10815 vp_p.n10814 0.296
R15172 vp_p.n10819 vp_p.n10818 0.296
R15173 vp_p.n10829 vp_p.n10828 0.296
R15174 vp_p.n10833 vp_p.n10832 0.296
R15175 vp_p.n10843 vp_p.n10842 0.296
R15176 vp_p.n10847 vp_p.n10846 0.296
R15177 vp_p.n10857 vp_p.n10856 0.296
R15178 vp_p.n10861 vp_p.n10860 0.296
R15179 vp_p.n10871 vp_p.n10870 0.296
R15180 vp_p.n10875 vp_p.n10874 0.296
R15181 vp_p.n10885 vp_p.n10884 0.296
R15182 vp_p.n10889 vp_p.n10888 0.296
R15183 vp_p.n10899 vp_p.n10898 0.296
R15184 vp_p.n10903 vp_p.n10902 0.296
R15185 vp_p.n10913 vp_p.n10912 0.296
R15186 vp_p.n10917 vp_p.n10916 0.296
R15187 vp_p.n10927 vp_p.n10926 0.296
R15188 vp_p.n10931 vp_p.n10930 0.296
R15189 vp_p.n10941 vp_p.n10940 0.296
R15190 vp_p.n10945 vp_p.n10944 0.296
R15191 vp_p.n10955 vp_p.n10954 0.296
R15192 vp_p.n10959 vp_p.n10958 0.296
R15193 vp_p.n10969 vp_p.n10968 0.296
R15194 vp_p.n10973 vp_p.n10972 0.296
R15195 vp_p.n10983 vp_p.n10982 0.296
R15196 vp_p.n10987 vp_p.n10986 0.296
R15197 vp_p.n10997 vp_p.n10996 0.296
R15198 vp_p.n11001 vp_p.n11000 0.296
R15199 vp_p.n11011 vp_p.n11010 0.296
R15200 vp_p.n11015 vp_p.n11014 0.296
R15201 vp_p.n11025 vp_p.n11024 0.296
R15202 vp_p.n11029 vp_p.n11028 0.296
R15203 vp_p.n11039 vp_p.n11038 0.296
R15204 vp_p.n11043 vp_p.n11042 0.296
R15205 vp_p.n11053 vp_p.n11052 0.296
R15206 vp_p.n11057 vp_p.n11056 0.296
R15207 vp_p.n11067 vp_p.n11066 0.296
R15208 vp_p.n11071 vp_p.n11070 0.296
R15209 vp_p.n11081 vp_p.n11080 0.296
R15210 vp_p.n11085 vp_p.n11084 0.296
R15211 vp_p.n11095 vp_p.n11094 0.296
R15212 vp_p.n11099 vp_p.n11098 0.296
R15213 vp_p.n11109 vp_p.n11108 0.296
R15214 vp_p.n11113 vp_p.n11112 0.296
R15215 vp_p.n11123 vp_p.n11122 0.296
R15216 vp_p.n11127 vp_p.n11126 0.296
R15217 vp_p.n11137 vp_p.n11136 0.296
R15218 vp_p.n11141 vp_p.n11140 0.296
R15219 vp_p.n11151 vp_p.n11150 0.296
R15220 vp_p.n11155 vp_p.n11154 0.296
R15221 vp_p.n11165 vp_p.n11164 0.296
R15222 vp_p.n11169 vp_p.n11168 0.296
R15223 vp_p.n11179 vp_p.n11178 0.296
R15224 vp_p.n11183 vp_p.n11182 0.296
R15225 vp_p.n11193 vp_p.n11192 0.296
R15226 vp_p.n11197 vp_p.n11196 0.296
R15227 vp_p.n11207 vp_p.n11206 0.296
R15228 vp_p.n11211 vp_p.n11210 0.296
R15229 vp_p.n11221 vp_p.n11220 0.296
R15230 vp_p.n11225 vp_p.n11224 0.296
R15231 vp_p.n11235 vp_p.n11234 0.296
R15232 vp_p.n11239 vp_p.n11238 0.296
R15233 vp_p.n11249 vp_p.n11248 0.296
R15234 vp_p.n11253 vp_p.n11252 0.296
R15235 vp_p.n11263 vp_p.n11262 0.296
R15236 vp_p.n11267 vp_p.n11266 0.296
R15237 vp_p.n11277 vp_p.n11276 0.296
R15238 vp_p.n11281 vp_p.n11280 0.296
R15239 vp_p.n11291 vp_p.n11290 0.296
R15240 vp_p.n11295 vp_p.n11294 0.296
R15241 vp_p.n11305 vp_p.n11304 0.296
R15242 vp_p.n11309 vp_p.n11308 0.296
R15243 vp_p.n11319 vp_p.n11318 0.296
R15244 vp_p.n11323 vp_p.n11322 0.296
R15245 vp_p.n11333 vp_p.n11332 0.296
R15246 vp_p.n11337 vp_p.n11336 0.296
R15247 vp_p.n11347 vp_p.n11346 0.296
R15248 vp_p.n11351 vp_p.n11350 0.296
R15249 vp_p.n11361 vp_p.n11360 0.296
R15250 vp_p.n11365 vp_p.n11364 0.296
R15251 vp_p.n11375 vp_p.n11374 0.296
R15252 vp_p.n11379 vp_p.n11378 0.296
R15253 vp_p.n11389 vp_p.n11388 0.296
R15254 vp_p.n11393 vp_p.n11392 0.296
R15255 vp_p.n11403 vp_p.n11402 0.296
R15256 vp_p.n11407 vp_p.n11406 0.296
R15257 vp_p.n11417 vp_p.n11416 0.296
R15258 vp_p.n11421 vp_p.n11420 0.296
R15259 vp_p.n11431 vp_p.n11430 0.296
R15260 vp_p.n11435 vp_p.n11434 0.296
R15261 vp_p.n11445 vp_p.n11444 0.296
R15262 vp_p.n11449 vp_p.n11448 0.296
R15263 vp_p.n11459 vp_p.n11458 0.296
R15264 vp_p.n11463 vp_p.n11462 0.296
R15265 vp_p.n11473 vp_p.n11472 0.296
R15266 vp_p.n11477 vp_p.n11476 0.296
R15267 vp_p.n11487 vp_p.n11486 0.296
R15268 vp_p.n11491 vp_p.n11490 0.296
R15269 vp_p.n11501 vp_p.n11500 0.296
R15270 vp_p.n11505 vp_p.n11504 0.296
R15271 vp_p.n11515 vp_p.n11514 0.296
R15272 vp_p.n11519 vp_p.n11518 0.296
R15273 vp_p.n11529 vp_p.n11528 0.296
R15274 vp_p.n11533 vp_p.n11532 0.296
R15275 vp_p.n11543 vp_p.n11542 0.296
R15276 vp_p.n11547 vp_p.n11546 0.296
R15277 vp_p.n11557 vp_p.n11556 0.296
R15278 vp_p.n11561 vp_p.n11560 0.296
R15279 vp_p.n11571 vp_p.n11570 0.296
R15280 vp_p.n11575 vp_p.n11574 0.296
R15281 vp_p.n11585 vp_p.n11584 0.296
R15282 vp_p.n11589 vp_p.n11588 0.296
R15283 vp_p.n11599 vp_p.n11598 0.296
R15284 vp_p.n11604 vp_p.n11603 0.296
R15285 vp_p.n11609 vp_p.n11608 0.296
R15286 vp_p.n11614 vp_p.n11613 0.296
R15287 vp_p.n11619 vp_p.n11618 0.296
R15288 vp_p.n11624 vp_p.n11623 0.296
R15289 vp_p.n11629 vp_p.n11628 0.296
R15290 vp_p.n11634 vp_p.n11633 0.296
R15291 vp_p.n11639 vp_p.n11638 0.296
R15292 vp_p.n11644 vp_p.n11643 0.296
R15293 vp_p.n11649 vp_p.n11648 0.296
R15294 vp_p.n11654 vp_p.n11653 0.296
R15295 vp_p.n11659 vp_p.n11658 0.296
R15296 vp_p.n16315 vp_p.n16314 0.296
R15297 vp_p.n16320 vp_p.n16319 0.296
R15298 vp_p.n16330 vp_p.n16329 0.296
R15299 vp_p.n16334 vp_p.n16333 0.296
R15300 vp_p.n16344 vp_p.n16343 0.296
R15301 vp_p.n16348 vp_p.n16347 0.296
R15302 vp_p.n16358 vp_p.n16357 0.296
R15303 vp_p.n16362 vp_p.n16361 0.296
R15304 vp_p.n16372 vp_p.n16371 0.296
R15305 vp_p.n16376 vp_p.n16375 0.296
R15306 vp_p.n16386 vp_p.n16385 0.296
R15307 vp_p.n16390 vp_p.n16389 0.296
R15308 vp_p.n16400 vp_p.n16399 0.296
R15309 vp_p.n16404 vp_p.n16403 0.296
R15310 vp_p.n16414 vp_p.n16413 0.296
R15311 vp_p.n16418 vp_p.n16417 0.296
R15312 vp_p.n16428 vp_p.n16427 0.296
R15313 vp_p.n16432 vp_p.n16431 0.296
R15314 vp_p.n16442 vp_p.n16441 0.296
R15315 vp_p.n16446 vp_p.n16445 0.296
R15316 vp_p.n16456 vp_p.n16455 0.296
R15317 vp_p.n16460 vp_p.n16459 0.296
R15318 vp_p.n16470 vp_p.n16469 0.296
R15319 vp_p.n16474 vp_p.n16473 0.296
R15320 vp_p.n16484 vp_p.n16483 0.296
R15321 vp_p.n16488 vp_p.n16487 0.296
R15322 vp_p.n16498 vp_p.n16497 0.296
R15323 vp_p.n16502 vp_p.n16501 0.296
R15324 vp_p.n16512 vp_p.n16511 0.296
R15325 vp_p.n16516 vp_p.n16515 0.296
R15326 vp_p.n16526 vp_p.n16525 0.296
R15327 vp_p.n16530 vp_p.n16529 0.296
R15328 vp_p.n16540 vp_p.n16539 0.296
R15329 vp_p.n16544 vp_p.n16543 0.296
R15330 vp_p.n16554 vp_p.n16553 0.296
R15331 vp_p.n16558 vp_p.n16557 0.296
R15332 vp_p.n16568 vp_p.n16567 0.296
R15333 vp_p.n16572 vp_p.n16571 0.296
R15334 vp_p.n16582 vp_p.n16581 0.296
R15335 vp_p.n16586 vp_p.n16585 0.296
R15336 vp_p.n16596 vp_p.n16595 0.296
R15337 vp_p.n16600 vp_p.n16599 0.296
R15338 vp_p.n16610 vp_p.n16609 0.296
R15339 vp_p.n16614 vp_p.n16613 0.296
R15340 vp_p.n16624 vp_p.n16623 0.296
R15341 vp_p.n16628 vp_p.n16627 0.296
R15342 vp_p.n16638 vp_p.n16637 0.296
R15343 vp_p.n16642 vp_p.n16641 0.296
R15344 vp_p.n16652 vp_p.n16651 0.296
R15345 vp_p.n16656 vp_p.n16655 0.296
R15346 vp_p.n16666 vp_p.n16665 0.296
R15347 vp_p.n16670 vp_p.n16669 0.296
R15348 vp_p.n16680 vp_p.n16679 0.296
R15349 vp_p.n16684 vp_p.n16683 0.296
R15350 vp_p.n16694 vp_p.n16693 0.296
R15351 vp_p.n16698 vp_p.n16697 0.296
R15352 vp_p.n16708 vp_p.n16707 0.296
R15353 vp_p.n16712 vp_p.n16711 0.296
R15354 vp_p.n16722 vp_p.n16721 0.296
R15355 vp_p.n16726 vp_p.n16725 0.296
R15356 vp_p.n16736 vp_p.n16735 0.296
R15357 vp_p.n16740 vp_p.n16739 0.296
R15358 vp_p.n16750 vp_p.n16749 0.296
R15359 vp_p.n16754 vp_p.n16753 0.296
R15360 vp_p.n16764 vp_p.n16763 0.296
R15361 vp_p.n16768 vp_p.n16767 0.296
R15362 vp_p.n16778 vp_p.n16777 0.296
R15363 vp_p.n16782 vp_p.n16781 0.296
R15364 vp_p.n16792 vp_p.n16791 0.296
R15365 vp_p.n16796 vp_p.n16795 0.296
R15366 vp_p.n16806 vp_p.n16805 0.296
R15367 vp_p.n16810 vp_p.n16809 0.296
R15368 vp_p.n16820 vp_p.n16819 0.296
R15369 vp_p.n16824 vp_p.n16823 0.296
R15370 vp_p.n16834 vp_p.n16833 0.296
R15371 vp_p.n16838 vp_p.n16837 0.296
R15372 vp_p.n16848 vp_p.n16847 0.296
R15373 vp_p.n16852 vp_p.n16851 0.296
R15374 vp_p.n16862 vp_p.n16861 0.296
R15375 vp_p.n16866 vp_p.n16865 0.296
R15376 vp_p.n16876 vp_p.n16875 0.296
R15377 vp_p.n16880 vp_p.n16879 0.296
R15378 vp_p.n16890 vp_p.n16889 0.296
R15379 vp_p.n16894 vp_p.n16893 0.296
R15380 vp_p.n16904 vp_p.n16903 0.296
R15381 vp_p.n16908 vp_p.n16907 0.296
R15382 vp_p.n16918 vp_p.n16917 0.296
R15383 vp_p.n16922 vp_p.n16921 0.296
R15384 vp_p.n16932 vp_p.n16931 0.296
R15385 vp_p.n16936 vp_p.n16935 0.296
R15386 vp_p.n16946 vp_p.n16945 0.296
R15387 vp_p.n16950 vp_p.n16949 0.296
R15388 vp_p.n16960 vp_p.n16959 0.296
R15389 vp_p.n16964 vp_p.n16963 0.296
R15390 vp_p.n16974 vp_p.n16973 0.296
R15391 vp_p.n16978 vp_p.n16977 0.296
R15392 vp_p.n16988 vp_p.n16987 0.296
R15393 vp_p.n16992 vp_p.n16991 0.296
R15394 vp_p.n17002 vp_p.n17001 0.296
R15395 vp_p.n17006 vp_p.n17005 0.296
R15396 vp_p.n17016 vp_p.n17015 0.296
R15397 vp_p.n17020 vp_p.n17019 0.296
R15398 vp_p.n17030 vp_p.n17029 0.296
R15399 vp_p.n17034 vp_p.n17033 0.296
R15400 vp_p.n17044 vp_p.n17043 0.296
R15401 vp_p.n17048 vp_p.n17047 0.296
R15402 vp_p.n17058 vp_p.n17057 0.296
R15403 vp_p.n17062 vp_p.n17061 0.296
R15404 vp_p.n17072 vp_p.n17071 0.296
R15405 vp_p.n17076 vp_p.n17075 0.296
R15406 vp_p.n17086 vp_p.n17085 0.296
R15407 vp_p.n17090 vp_p.n17089 0.296
R15408 vp_p.n17100 vp_p.n17099 0.296
R15409 vp_p.n17104 vp_p.n17103 0.296
R15410 vp_p.n17114 vp_p.n17113 0.296
R15411 vp_p.n17118 vp_p.n17117 0.296
R15412 vp_p.n17128 vp_p.n17127 0.296
R15413 vp_p.n17132 vp_p.n17131 0.296
R15414 vp_p.n17142 vp_p.n17141 0.296
R15415 vp_p.n17146 vp_p.n17145 0.296
R15416 vp_p.n17156 vp_p.n17155 0.296
R15417 vp_p.n17160 vp_p.n17159 0.296
R15418 vp_p.n17170 vp_p.n17169 0.296
R15419 vp_p.n17174 vp_p.n17173 0.296
R15420 vp_p.n17184 vp_p.n17183 0.296
R15421 vp_p.n17188 vp_p.n17187 0.296
R15422 vp_p.n17198 vp_p.n17197 0.296
R15423 vp_p.n17202 vp_p.n17201 0.296
R15424 vp_p.n17212 vp_p.n17211 0.296
R15425 vp_p.n17216 vp_p.n17215 0.296
R15426 vp_p.n17226 vp_p.n17225 0.296
R15427 vp_p.n17230 vp_p.n17229 0.296
R15428 vp_p.n17240 vp_p.n17239 0.296
R15429 vp_p.n17244 vp_p.n17243 0.296
R15430 vp_p.n17254 vp_p.n17253 0.296
R15431 vp_p.n17258 vp_p.n17257 0.296
R15432 vp_p.n17262 vp_p.n17261 0.296
R15433 vp_p.n17272 vp_p.n17271 0.296
R15434 vp_p.n17277 vp_p.n17276 0.296
R15435 vp_p.n17282 vp_p.n17281 0.296
R15436 vp_p.n17287 vp_p.n17286 0.296
R15437 vp_p.n17292 vp_p.n17291 0.296
R15438 vp_p.n17297 vp_p.n17296 0.296
R15439 vp_p.n17302 vp_p.n17301 0.296
R15440 vp_p.n17307 vp_p.n17306 0.296
R15441 vp_p.n17312 vp_p.n17311 0.296
R15442 vp_p.n17317 vp_p.n17316 0.296
R15443 vp_p.n17322 vp_p.n17321 0.296
R15444 vp_p.n17327 vp_p.n17326 0.296
R15445 vp_p.n9209 vp_p.n9208 0.296
R15446 vp_p.n9214 vp_p.n9213 0.296
R15447 vp_p.n9224 vp_p.n9223 0.296
R15448 vp_p.n9228 vp_p.n9227 0.296
R15449 vp_p.n9238 vp_p.n9237 0.296
R15450 vp_p.n9242 vp_p.n9241 0.296
R15451 vp_p.n9252 vp_p.n9251 0.296
R15452 vp_p.n9256 vp_p.n9255 0.296
R15453 vp_p.n9266 vp_p.n9265 0.296
R15454 vp_p.n9270 vp_p.n9269 0.296
R15455 vp_p.n9280 vp_p.n9279 0.296
R15456 vp_p.n9284 vp_p.n9283 0.296
R15457 vp_p.n9294 vp_p.n9293 0.296
R15458 vp_p.n9298 vp_p.n9297 0.296
R15459 vp_p.n9308 vp_p.n9307 0.296
R15460 vp_p.n9312 vp_p.n9311 0.296
R15461 vp_p.n9322 vp_p.n9321 0.296
R15462 vp_p.n9326 vp_p.n9325 0.296
R15463 vp_p.n9336 vp_p.n9335 0.296
R15464 vp_p.n9340 vp_p.n9339 0.296
R15465 vp_p.n9350 vp_p.n9349 0.296
R15466 vp_p.n9354 vp_p.n9353 0.296
R15467 vp_p.n9364 vp_p.n9363 0.296
R15468 vp_p.n9368 vp_p.n9367 0.296
R15469 vp_p.n9378 vp_p.n9377 0.296
R15470 vp_p.n9382 vp_p.n9381 0.296
R15471 vp_p.n9392 vp_p.n9391 0.296
R15472 vp_p.n9396 vp_p.n9395 0.296
R15473 vp_p.n9406 vp_p.n9405 0.296
R15474 vp_p.n9410 vp_p.n9409 0.296
R15475 vp_p.n9420 vp_p.n9419 0.296
R15476 vp_p.n9424 vp_p.n9423 0.296
R15477 vp_p.n9434 vp_p.n9433 0.296
R15478 vp_p.n9438 vp_p.n9437 0.296
R15479 vp_p.n9448 vp_p.n9447 0.296
R15480 vp_p.n9452 vp_p.n9451 0.296
R15481 vp_p.n9462 vp_p.n9461 0.296
R15482 vp_p.n9466 vp_p.n9465 0.296
R15483 vp_p.n9476 vp_p.n9475 0.296
R15484 vp_p.n9480 vp_p.n9479 0.296
R15485 vp_p.n9490 vp_p.n9489 0.296
R15486 vp_p.n9494 vp_p.n9493 0.296
R15487 vp_p.n9504 vp_p.n9503 0.296
R15488 vp_p.n9508 vp_p.n9507 0.296
R15489 vp_p.n9518 vp_p.n9517 0.296
R15490 vp_p.n9522 vp_p.n9521 0.296
R15491 vp_p.n9532 vp_p.n9531 0.296
R15492 vp_p.n9536 vp_p.n9535 0.296
R15493 vp_p.n9546 vp_p.n9545 0.296
R15494 vp_p.n9550 vp_p.n9549 0.296
R15495 vp_p.n9560 vp_p.n9559 0.296
R15496 vp_p.n9564 vp_p.n9563 0.296
R15497 vp_p.n9574 vp_p.n9573 0.296
R15498 vp_p.n9578 vp_p.n9577 0.296
R15499 vp_p.n9588 vp_p.n9587 0.296
R15500 vp_p.n9592 vp_p.n9591 0.296
R15501 vp_p.n9602 vp_p.n9601 0.296
R15502 vp_p.n9606 vp_p.n9605 0.296
R15503 vp_p.n9616 vp_p.n9615 0.296
R15504 vp_p.n9620 vp_p.n9619 0.296
R15505 vp_p.n9630 vp_p.n9629 0.296
R15506 vp_p.n9634 vp_p.n9633 0.296
R15507 vp_p.n9644 vp_p.n9643 0.296
R15508 vp_p.n9648 vp_p.n9647 0.296
R15509 vp_p.n9658 vp_p.n9657 0.296
R15510 vp_p.n9662 vp_p.n9661 0.296
R15511 vp_p.n9672 vp_p.n9671 0.296
R15512 vp_p.n9676 vp_p.n9675 0.296
R15513 vp_p.n9686 vp_p.n9685 0.296
R15514 vp_p.n9690 vp_p.n9689 0.296
R15515 vp_p.n9700 vp_p.n9699 0.296
R15516 vp_p.n9704 vp_p.n9703 0.296
R15517 vp_p.n9714 vp_p.n9713 0.296
R15518 vp_p.n9718 vp_p.n9717 0.296
R15519 vp_p.n9728 vp_p.n9727 0.296
R15520 vp_p.n9732 vp_p.n9731 0.296
R15521 vp_p.n9742 vp_p.n9741 0.296
R15522 vp_p.n9746 vp_p.n9745 0.296
R15523 vp_p.n9756 vp_p.n9755 0.296
R15524 vp_p.n9760 vp_p.n9759 0.296
R15525 vp_p.n9770 vp_p.n9769 0.296
R15526 vp_p.n9774 vp_p.n9773 0.296
R15527 vp_p.n9784 vp_p.n9783 0.296
R15528 vp_p.n9788 vp_p.n9787 0.296
R15529 vp_p.n9798 vp_p.n9797 0.296
R15530 vp_p.n9802 vp_p.n9801 0.296
R15531 vp_p.n9812 vp_p.n9811 0.296
R15532 vp_p.n9816 vp_p.n9815 0.296
R15533 vp_p.n9826 vp_p.n9825 0.296
R15534 vp_p.n9830 vp_p.n9829 0.296
R15535 vp_p.n9840 vp_p.n9839 0.296
R15536 vp_p.n9844 vp_p.n9843 0.296
R15537 vp_p.n9854 vp_p.n9853 0.296
R15538 vp_p.n9858 vp_p.n9857 0.296
R15539 vp_p.n9868 vp_p.n9867 0.296
R15540 vp_p.n9872 vp_p.n9871 0.296
R15541 vp_p.n9882 vp_p.n9881 0.296
R15542 vp_p.n9886 vp_p.n9885 0.296
R15543 vp_p.n9896 vp_p.n9895 0.296
R15544 vp_p.n9900 vp_p.n9899 0.296
R15545 vp_p.n9910 vp_p.n9909 0.296
R15546 vp_p.n9914 vp_p.n9913 0.296
R15547 vp_p.n9924 vp_p.n9923 0.296
R15548 vp_p.n9928 vp_p.n9927 0.296
R15549 vp_p.n9938 vp_p.n9937 0.296
R15550 vp_p.n9942 vp_p.n9941 0.296
R15551 vp_p.n9952 vp_p.n9951 0.296
R15552 vp_p.n9956 vp_p.n9955 0.296
R15553 vp_p.n9966 vp_p.n9965 0.296
R15554 vp_p.n9970 vp_p.n9969 0.296
R15555 vp_p.n9980 vp_p.n9979 0.296
R15556 vp_p.n9984 vp_p.n9983 0.296
R15557 vp_p.n9994 vp_p.n9993 0.296
R15558 vp_p.n9998 vp_p.n9997 0.296
R15559 vp_p.n10008 vp_p.n10007 0.296
R15560 vp_p.n10012 vp_p.n10011 0.296
R15561 vp_p.n10022 vp_p.n10021 0.296
R15562 vp_p.n10026 vp_p.n10025 0.296
R15563 vp_p.n10036 vp_p.n10035 0.296
R15564 vp_p.n10040 vp_p.n10039 0.296
R15565 vp_p.n10050 vp_p.n10049 0.296
R15566 vp_p.n10054 vp_p.n10053 0.296
R15567 vp_p.n10064 vp_p.n10063 0.296
R15568 vp_p.n10068 vp_p.n10067 0.296
R15569 vp_p.n10078 vp_p.n10077 0.296
R15570 vp_p.n10082 vp_p.n10081 0.296
R15571 vp_p.n10092 vp_p.n10091 0.296
R15572 vp_p.n10096 vp_p.n10095 0.296
R15573 vp_p.n10106 vp_p.n10105 0.296
R15574 vp_p.n10110 vp_p.n10109 0.296
R15575 vp_p.n10120 vp_p.n10119 0.296
R15576 vp_p.n10124 vp_p.n10123 0.296
R15577 vp_p.n10134 vp_p.n10133 0.296
R15578 vp_p.n10138 vp_p.n10137 0.296
R15579 vp_p.n10148 vp_p.n10147 0.296
R15580 vp_p.n10152 vp_p.n10151 0.296
R15581 vp_p.n10162 vp_p.n10161 0.296
R15582 vp_p.n10166 vp_p.n10165 0.296
R15583 vp_p.n10176 vp_p.n10175 0.296
R15584 vp_p.n10181 vp_p.n10180 0.296
R15585 vp_p.n10186 vp_p.n10185 0.296
R15586 vp_p.n10191 vp_p.n10190 0.296
R15587 vp_p.n10196 vp_p.n10195 0.296
R15588 vp_p.n10201 vp_p.n10200 0.296
R15589 vp_p.n10206 vp_p.n10205 0.296
R15590 vp_p.n10211 vp_p.n10210 0.296
R15591 vp_p.n10216 vp_p.n10215 0.296
R15592 vp_p.n10221 vp_p.n10220 0.296
R15593 vp_p.n10226 vp_p.n10225 0.296
R15594 vp_p.n17742 vp_p.n17741 0.296
R15595 vp_p.n17747 vp_p.n17746 0.296
R15596 vp_p.n17757 vp_p.n17756 0.296
R15597 vp_p.n17761 vp_p.n17760 0.296
R15598 vp_p.n17771 vp_p.n17770 0.296
R15599 vp_p.n17775 vp_p.n17774 0.296
R15600 vp_p.n17785 vp_p.n17784 0.296
R15601 vp_p.n17789 vp_p.n17788 0.296
R15602 vp_p.n17799 vp_p.n17798 0.296
R15603 vp_p.n17803 vp_p.n17802 0.296
R15604 vp_p.n17813 vp_p.n17812 0.296
R15605 vp_p.n17817 vp_p.n17816 0.296
R15606 vp_p.n17827 vp_p.n17826 0.296
R15607 vp_p.n17831 vp_p.n17830 0.296
R15608 vp_p.n17841 vp_p.n17840 0.296
R15609 vp_p.n17845 vp_p.n17844 0.296
R15610 vp_p.n17855 vp_p.n17854 0.296
R15611 vp_p.n17859 vp_p.n17858 0.296
R15612 vp_p.n17869 vp_p.n17868 0.296
R15613 vp_p.n17873 vp_p.n17872 0.296
R15614 vp_p.n17883 vp_p.n17882 0.296
R15615 vp_p.n17887 vp_p.n17886 0.296
R15616 vp_p.n17897 vp_p.n17896 0.296
R15617 vp_p.n17901 vp_p.n17900 0.296
R15618 vp_p.n17911 vp_p.n17910 0.296
R15619 vp_p.n17915 vp_p.n17914 0.296
R15620 vp_p.n17925 vp_p.n17924 0.296
R15621 vp_p.n17929 vp_p.n17928 0.296
R15622 vp_p.n17939 vp_p.n17938 0.296
R15623 vp_p.n17943 vp_p.n17942 0.296
R15624 vp_p.n17953 vp_p.n17952 0.296
R15625 vp_p.n17957 vp_p.n17956 0.296
R15626 vp_p.n17967 vp_p.n17966 0.296
R15627 vp_p.n17971 vp_p.n17970 0.296
R15628 vp_p.n17981 vp_p.n17980 0.296
R15629 vp_p.n17985 vp_p.n17984 0.296
R15630 vp_p.n17995 vp_p.n17994 0.296
R15631 vp_p.n17999 vp_p.n17998 0.296
R15632 vp_p.n18009 vp_p.n18008 0.296
R15633 vp_p.n18013 vp_p.n18012 0.296
R15634 vp_p.n18023 vp_p.n18022 0.296
R15635 vp_p.n18027 vp_p.n18026 0.296
R15636 vp_p.n18037 vp_p.n18036 0.296
R15637 vp_p.n18041 vp_p.n18040 0.296
R15638 vp_p.n18051 vp_p.n18050 0.296
R15639 vp_p.n18055 vp_p.n18054 0.296
R15640 vp_p.n18065 vp_p.n18064 0.296
R15641 vp_p.n18069 vp_p.n18068 0.296
R15642 vp_p.n18079 vp_p.n18078 0.296
R15643 vp_p.n18083 vp_p.n18082 0.296
R15644 vp_p.n18093 vp_p.n18092 0.296
R15645 vp_p.n18097 vp_p.n18096 0.296
R15646 vp_p.n18107 vp_p.n18106 0.296
R15647 vp_p.n18111 vp_p.n18110 0.296
R15648 vp_p.n18121 vp_p.n18120 0.296
R15649 vp_p.n18125 vp_p.n18124 0.296
R15650 vp_p.n18135 vp_p.n18134 0.296
R15651 vp_p.n18139 vp_p.n18138 0.296
R15652 vp_p.n18149 vp_p.n18148 0.296
R15653 vp_p.n18153 vp_p.n18152 0.296
R15654 vp_p.n18163 vp_p.n18162 0.296
R15655 vp_p.n18167 vp_p.n18166 0.296
R15656 vp_p.n18177 vp_p.n18176 0.296
R15657 vp_p.n18181 vp_p.n18180 0.296
R15658 vp_p.n18191 vp_p.n18190 0.296
R15659 vp_p.n18195 vp_p.n18194 0.296
R15660 vp_p.n18205 vp_p.n18204 0.296
R15661 vp_p.n18209 vp_p.n18208 0.296
R15662 vp_p.n18219 vp_p.n18218 0.296
R15663 vp_p.n18223 vp_p.n18222 0.296
R15664 vp_p.n18233 vp_p.n18232 0.296
R15665 vp_p.n18237 vp_p.n18236 0.296
R15666 vp_p.n18247 vp_p.n18246 0.296
R15667 vp_p.n18251 vp_p.n18250 0.296
R15668 vp_p.n18261 vp_p.n18260 0.296
R15669 vp_p.n18265 vp_p.n18264 0.296
R15670 vp_p.n18275 vp_p.n18274 0.296
R15671 vp_p.n18279 vp_p.n18278 0.296
R15672 vp_p.n18289 vp_p.n18288 0.296
R15673 vp_p.n18293 vp_p.n18292 0.296
R15674 vp_p.n18303 vp_p.n18302 0.296
R15675 vp_p.n18307 vp_p.n18306 0.296
R15676 vp_p.n18317 vp_p.n18316 0.296
R15677 vp_p.n18321 vp_p.n18320 0.296
R15678 vp_p.n18331 vp_p.n18330 0.296
R15679 vp_p.n18335 vp_p.n18334 0.296
R15680 vp_p.n18345 vp_p.n18344 0.296
R15681 vp_p.n18349 vp_p.n18348 0.296
R15682 vp_p.n18359 vp_p.n18358 0.296
R15683 vp_p.n18363 vp_p.n18362 0.296
R15684 vp_p.n18373 vp_p.n18372 0.296
R15685 vp_p.n18377 vp_p.n18376 0.296
R15686 vp_p.n18387 vp_p.n18386 0.296
R15687 vp_p.n18391 vp_p.n18390 0.296
R15688 vp_p.n18401 vp_p.n18400 0.296
R15689 vp_p.n18405 vp_p.n18404 0.296
R15690 vp_p.n18415 vp_p.n18414 0.296
R15691 vp_p.n18419 vp_p.n18418 0.296
R15692 vp_p.n18429 vp_p.n18428 0.296
R15693 vp_p.n18433 vp_p.n18432 0.296
R15694 vp_p.n18443 vp_p.n18442 0.296
R15695 vp_p.n18447 vp_p.n18446 0.296
R15696 vp_p.n18457 vp_p.n18456 0.296
R15697 vp_p.n18461 vp_p.n18460 0.296
R15698 vp_p.n18471 vp_p.n18470 0.296
R15699 vp_p.n18475 vp_p.n18474 0.296
R15700 vp_p.n18485 vp_p.n18484 0.296
R15701 vp_p.n18489 vp_p.n18488 0.296
R15702 vp_p.n18499 vp_p.n18498 0.296
R15703 vp_p.n18503 vp_p.n18502 0.296
R15704 vp_p.n18513 vp_p.n18512 0.296
R15705 vp_p.n18517 vp_p.n18516 0.296
R15706 vp_p.n18527 vp_p.n18526 0.296
R15707 vp_p.n18531 vp_p.n18530 0.296
R15708 vp_p.n18541 vp_p.n18540 0.296
R15709 vp_p.n18545 vp_p.n18544 0.296
R15710 vp_p.n18555 vp_p.n18554 0.296
R15711 vp_p.n18559 vp_p.n18558 0.296
R15712 vp_p.n18569 vp_p.n18568 0.296
R15713 vp_p.n18573 vp_p.n18572 0.296
R15714 vp_p.n18583 vp_p.n18582 0.296
R15715 vp_p.n18587 vp_p.n18586 0.296
R15716 vp_p.n18597 vp_p.n18596 0.296
R15717 vp_p.n18601 vp_p.n18600 0.296
R15718 vp_p.n18611 vp_p.n18610 0.296
R15719 vp_p.n18615 vp_p.n18614 0.296
R15720 vp_p.n18625 vp_p.n18624 0.296
R15721 vp_p.n18629 vp_p.n18628 0.296
R15722 vp_p.n18639 vp_p.n18638 0.296
R15723 vp_p.n18643 vp_p.n18642 0.296
R15724 vp_p.n18653 vp_p.n18652 0.296
R15725 vp_p.n18657 vp_p.n18656 0.296
R15726 vp_p.n18667 vp_p.n18666 0.296
R15727 vp_p.n18671 vp_p.n18670 0.296
R15728 vp_p.n18681 vp_p.n18680 0.296
R15729 vp_p.n18685 vp_p.n18684 0.296
R15730 vp_p.n18695 vp_p.n18694 0.296
R15731 vp_p.n18699 vp_p.n18698 0.296
R15732 vp_p.n18703 vp_p.n18702 0.296
R15733 vp_p.n18713 vp_p.n18712 0.296
R15734 vp_p.n18718 vp_p.n18717 0.296
R15735 vp_p.n18723 vp_p.n18722 0.296
R15736 vp_p.n18728 vp_p.n18727 0.296
R15737 vp_p.n18733 vp_p.n18732 0.296
R15738 vp_p.n18738 vp_p.n18737 0.296
R15739 vp_p.n18743 vp_p.n18742 0.296
R15740 vp_p.n18748 vp_p.n18747 0.296
R15741 vp_p.n18753 vp_p.n18752 0.296
R15742 vp_p.n18758 vp_p.n18757 0.296
R15743 vp_p.n463 vp_p.n462 0.296
R15744 vp_p.n468 vp_p.n467 0.296
R15745 vp_p.n478 vp_p.n477 0.296
R15746 vp_p.n482 vp_p.n481 0.296
R15747 vp_p.n492 vp_p.n491 0.296
R15748 vp_p.n496 vp_p.n495 0.296
R15749 vp_p.n506 vp_p.n505 0.296
R15750 vp_p.n510 vp_p.n509 0.296
R15751 vp_p.n520 vp_p.n519 0.296
R15752 vp_p.n524 vp_p.n523 0.296
R15753 vp_p.n534 vp_p.n533 0.296
R15754 vp_p.n538 vp_p.n537 0.296
R15755 vp_p.n548 vp_p.n547 0.296
R15756 vp_p.n552 vp_p.n551 0.296
R15757 vp_p.n562 vp_p.n561 0.296
R15758 vp_p.n566 vp_p.n565 0.296
R15759 vp_p.n576 vp_p.n575 0.296
R15760 vp_p.n580 vp_p.n579 0.296
R15761 vp_p.n590 vp_p.n589 0.296
R15762 vp_p.n594 vp_p.n593 0.296
R15763 vp_p.n604 vp_p.n603 0.296
R15764 vp_p.n608 vp_p.n607 0.296
R15765 vp_p.n618 vp_p.n617 0.296
R15766 vp_p.n622 vp_p.n621 0.296
R15767 vp_p.n632 vp_p.n631 0.296
R15768 vp_p.n636 vp_p.n635 0.296
R15769 vp_p.n646 vp_p.n645 0.296
R15770 vp_p.n650 vp_p.n649 0.296
R15771 vp_p.n660 vp_p.n659 0.296
R15772 vp_p.n664 vp_p.n663 0.296
R15773 vp_p.n674 vp_p.n673 0.296
R15774 vp_p.n678 vp_p.n677 0.296
R15775 vp_p.n688 vp_p.n687 0.296
R15776 vp_p.n692 vp_p.n691 0.296
R15777 vp_p.n702 vp_p.n701 0.296
R15778 vp_p.n706 vp_p.n705 0.296
R15779 vp_p.n716 vp_p.n715 0.296
R15780 vp_p.n720 vp_p.n719 0.296
R15781 vp_p.n730 vp_p.n729 0.296
R15782 vp_p.n734 vp_p.n733 0.296
R15783 vp_p.n744 vp_p.n743 0.296
R15784 vp_p.n748 vp_p.n747 0.296
R15785 vp_p.n758 vp_p.n757 0.296
R15786 vp_p.n762 vp_p.n761 0.296
R15787 vp_p.n772 vp_p.n771 0.296
R15788 vp_p.n776 vp_p.n775 0.296
R15789 vp_p.n786 vp_p.n785 0.296
R15790 vp_p.n790 vp_p.n789 0.296
R15791 vp_p.n800 vp_p.n799 0.296
R15792 vp_p.n804 vp_p.n803 0.296
R15793 vp_p.n814 vp_p.n813 0.296
R15794 vp_p.n818 vp_p.n817 0.296
R15795 vp_p.n828 vp_p.n827 0.296
R15796 vp_p.n832 vp_p.n831 0.296
R15797 vp_p.n842 vp_p.n841 0.296
R15798 vp_p.n846 vp_p.n845 0.296
R15799 vp_p.n856 vp_p.n855 0.296
R15800 vp_p.n860 vp_p.n859 0.296
R15801 vp_p.n870 vp_p.n869 0.296
R15802 vp_p.n874 vp_p.n873 0.296
R15803 vp_p.n884 vp_p.n883 0.296
R15804 vp_p.n888 vp_p.n887 0.296
R15805 vp_p.n898 vp_p.n897 0.296
R15806 vp_p.n902 vp_p.n901 0.296
R15807 vp_p.n912 vp_p.n911 0.296
R15808 vp_p.n916 vp_p.n915 0.296
R15809 vp_p.n926 vp_p.n925 0.296
R15810 vp_p.n930 vp_p.n929 0.296
R15811 vp_p.n940 vp_p.n939 0.296
R15812 vp_p.n944 vp_p.n943 0.296
R15813 vp_p.n954 vp_p.n953 0.296
R15814 vp_p.n958 vp_p.n957 0.296
R15815 vp_p.n968 vp_p.n967 0.296
R15816 vp_p.n972 vp_p.n971 0.296
R15817 vp_p.n982 vp_p.n981 0.296
R15818 vp_p.n986 vp_p.n985 0.296
R15819 vp_p.n996 vp_p.n995 0.296
R15820 vp_p.n1000 vp_p.n999 0.296
R15821 vp_p.n1010 vp_p.n1009 0.296
R15822 vp_p.n1014 vp_p.n1013 0.296
R15823 vp_p.n1024 vp_p.n1023 0.296
R15824 vp_p.n1028 vp_p.n1027 0.296
R15825 vp_p.n1038 vp_p.n1037 0.296
R15826 vp_p.n1042 vp_p.n1041 0.296
R15827 vp_p.n1052 vp_p.n1051 0.296
R15828 vp_p.n1056 vp_p.n1055 0.296
R15829 vp_p.n1066 vp_p.n1065 0.296
R15830 vp_p.n1070 vp_p.n1069 0.296
R15831 vp_p.n1080 vp_p.n1079 0.296
R15832 vp_p.n1084 vp_p.n1083 0.296
R15833 vp_p.n1094 vp_p.n1093 0.296
R15834 vp_p.n1098 vp_p.n1097 0.296
R15835 vp_p.n1108 vp_p.n1107 0.296
R15836 vp_p.n1112 vp_p.n1111 0.296
R15837 vp_p.n1122 vp_p.n1121 0.296
R15838 vp_p.n1126 vp_p.n1125 0.296
R15839 vp_p.n1136 vp_p.n1135 0.296
R15840 vp_p.n1140 vp_p.n1139 0.296
R15841 vp_p.n1150 vp_p.n1149 0.296
R15842 vp_p.n1154 vp_p.n1153 0.296
R15843 vp_p.n1164 vp_p.n1163 0.296
R15844 vp_p.n1168 vp_p.n1167 0.296
R15845 vp_p.n1178 vp_p.n1177 0.296
R15846 vp_p.n1182 vp_p.n1181 0.296
R15847 vp_p.n1192 vp_p.n1191 0.296
R15848 vp_p.n1196 vp_p.n1195 0.296
R15849 vp_p.n1206 vp_p.n1205 0.296
R15850 vp_p.n1210 vp_p.n1209 0.296
R15851 vp_p.n1220 vp_p.n1219 0.296
R15852 vp_p.n1224 vp_p.n1223 0.296
R15853 vp_p.n1234 vp_p.n1233 0.296
R15854 vp_p.n1238 vp_p.n1237 0.296
R15855 vp_p.n1248 vp_p.n1247 0.296
R15856 vp_p.n1252 vp_p.n1251 0.296
R15857 vp_p.n1262 vp_p.n1261 0.296
R15858 vp_p.n1266 vp_p.n1265 0.296
R15859 vp_p.n1276 vp_p.n1275 0.296
R15860 vp_p.n1280 vp_p.n1279 0.296
R15861 vp_p.n1290 vp_p.n1289 0.296
R15862 vp_p.n1294 vp_p.n1293 0.296
R15863 vp_p.n1304 vp_p.n1303 0.296
R15864 vp_p.n1308 vp_p.n1307 0.296
R15865 vp_p.n1318 vp_p.n1317 0.296
R15866 vp_p.n1322 vp_p.n1321 0.296
R15867 vp_p.n1332 vp_p.n1331 0.296
R15868 vp_p.n1336 vp_p.n1335 0.296
R15869 vp_p.n1346 vp_p.n1345 0.296
R15870 vp_p.n1350 vp_p.n1349 0.296
R15871 vp_p.n1360 vp_p.n1359 0.296
R15872 vp_p.n1364 vp_p.n1363 0.296
R15873 vp_p.n1374 vp_p.n1373 0.296
R15874 vp_p.n1378 vp_p.n1377 0.296
R15875 vp_p.n1388 vp_p.n1387 0.296
R15876 vp_p.n1392 vp_p.n1391 0.296
R15877 vp_p.n1402 vp_p.n1401 0.296
R15878 vp_p.n1406 vp_p.n1405 0.296
R15879 vp_p.n1416 vp_p.n1415 0.296
R15880 vp_p.n1420 vp_p.n1419 0.296
R15881 vp_p.n1430 vp_p.n1429 0.296
R15882 vp_p.n1434 vp_p.n1433 0.296
R15883 vp_p.n1444 vp_p.n1443 0.296
R15884 vp_p.n1449 vp_p.n1448 0.296
R15885 vp_p.n1454 vp_p.n1453 0.296
R15886 vp_p.n1459 vp_p.n1458 0.296
R15887 vp_p.n1464 vp_p.n1463 0.296
R15888 vp_p.n1469 vp_p.n1468 0.296
R15889 vp_p.n1474 vp_p.n1473 0.296
R15890 vp_p.n1479 vp_p.n1478 0.296
R15891 vp_p.n1484 vp_p.n1483 0.296
R15892 vp_p.n19168 vp_p.n19167 0.296
R15893 vp_p.n19173 vp_p.n19172 0.296
R15894 vp_p.n19183 vp_p.n19182 0.296
R15895 vp_p.n19187 vp_p.n19186 0.296
R15896 vp_p.n19197 vp_p.n19196 0.296
R15897 vp_p.n19201 vp_p.n19200 0.296
R15898 vp_p.n19211 vp_p.n19210 0.296
R15899 vp_p.n19215 vp_p.n19214 0.296
R15900 vp_p.n19225 vp_p.n19224 0.296
R15901 vp_p.n19229 vp_p.n19228 0.296
R15902 vp_p.n19239 vp_p.n19238 0.296
R15903 vp_p.n19243 vp_p.n19242 0.296
R15904 vp_p.n19253 vp_p.n19252 0.296
R15905 vp_p.n19257 vp_p.n19256 0.296
R15906 vp_p.n19267 vp_p.n19266 0.296
R15907 vp_p.n19271 vp_p.n19270 0.296
R15908 vp_p.n19281 vp_p.n19280 0.296
R15909 vp_p.n19285 vp_p.n19284 0.296
R15910 vp_p.n19295 vp_p.n19294 0.296
R15911 vp_p.n19299 vp_p.n19298 0.296
R15912 vp_p.n19309 vp_p.n19308 0.296
R15913 vp_p.n19313 vp_p.n19312 0.296
R15914 vp_p.n19323 vp_p.n19322 0.296
R15915 vp_p.n19327 vp_p.n19326 0.296
R15916 vp_p.n19337 vp_p.n19336 0.296
R15917 vp_p.n19341 vp_p.n19340 0.296
R15918 vp_p.n19351 vp_p.n19350 0.296
R15919 vp_p.n19355 vp_p.n19354 0.296
R15920 vp_p.n19365 vp_p.n19364 0.296
R15921 vp_p.n19369 vp_p.n19368 0.296
R15922 vp_p.n19379 vp_p.n19378 0.296
R15923 vp_p.n19383 vp_p.n19382 0.296
R15924 vp_p.n19393 vp_p.n19392 0.296
R15925 vp_p.n19397 vp_p.n19396 0.296
R15926 vp_p.n19407 vp_p.n19406 0.296
R15927 vp_p.n19411 vp_p.n19410 0.296
R15928 vp_p.n19421 vp_p.n19420 0.296
R15929 vp_p.n19425 vp_p.n19424 0.296
R15930 vp_p.n19435 vp_p.n19434 0.296
R15931 vp_p.n19439 vp_p.n19438 0.296
R15932 vp_p.n19449 vp_p.n19448 0.296
R15933 vp_p.n19453 vp_p.n19452 0.296
R15934 vp_p.n19463 vp_p.n19462 0.296
R15935 vp_p.n19467 vp_p.n19466 0.296
R15936 vp_p.n19477 vp_p.n19476 0.296
R15937 vp_p.n19481 vp_p.n19480 0.296
R15938 vp_p.n19491 vp_p.n19490 0.296
R15939 vp_p.n19495 vp_p.n19494 0.296
R15940 vp_p.n19505 vp_p.n19504 0.296
R15941 vp_p.n19509 vp_p.n19508 0.296
R15942 vp_p.n19519 vp_p.n19518 0.296
R15943 vp_p.n19523 vp_p.n19522 0.296
R15944 vp_p.n19533 vp_p.n19532 0.296
R15945 vp_p.n19537 vp_p.n19536 0.296
R15946 vp_p.n19547 vp_p.n19546 0.296
R15947 vp_p.n19551 vp_p.n19550 0.296
R15948 vp_p.n19561 vp_p.n19560 0.296
R15949 vp_p.n19565 vp_p.n19564 0.296
R15950 vp_p.n19575 vp_p.n19574 0.296
R15951 vp_p.n19579 vp_p.n19578 0.296
R15952 vp_p.n19589 vp_p.n19588 0.296
R15953 vp_p.n19593 vp_p.n19592 0.296
R15954 vp_p.n19603 vp_p.n19602 0.296
R15955 vp_p.n19607 vp_p.n19606 0.296
R15956 vp_p.n19617 vp_p.n19616 0.296
R15957 vp_p.n19621 vp_p.n19620 0.296
R15958 vp_p.n19631 vp_p.n19630 0.296
R15959 vp_p.n19635 vp_p.n19634 0.296
R15960 vp_p.n19645 vp_p.n19644 0.296
R15961 vp_p.n19649 vp_p.n19648 0.296
R15962 vp_p.n19659 vp_p.n19658 0.296
R15963 vp_p.n19663 vp_p.n19662 0.296
R15964 vp_p.n19673 vp_p.n19672 0.296
R15965 vp_p.n19677 vp_p.n19676 0.296
R15966 vp_p.n19687 vp_p.n19686 0.296
R15967 vp_p.n19691 vp_p.n19690 0.296
R15968 vp_p.n19701 vp_p.n19700 0.296
R15969 vp_p.n19705 vp_p.n19704 0.296
R15970 vp_p.n19715 vp_p.n19714 0.296
R15971 vp_p.n19719 vp_p.n19718 0.296
R15972 vp_p.n19729 vp_p.n19728 0.296
R15973 vp_p.n19733 vp_p.n19732 0.296
R15974 vp_p.n19743 vp_p.n19742 0.296
R15975 vp_p.n19747 vp_p.n19746 0.296
R15976 vp_p.n19757 vp_p.n19756 0.296
R15977 vp_p.n19761 vp_p.n19760 0.296
R15978 vp_p.n19771 vp_p.n19770 0.296
R15979 vp_p.n19775 vp_p.n19774 0.296
R15980 vp_p.n19785 vp_p.n19784 0.296
R15981 vp_p.n19789 vp_p.n19788 0.296
R15982 vp_p.n19799 vp_p.n19798 0.296
R15983 vp_p.n19803 vp_p.n19802 0.296
R15984 vp_p.n19813 vp_p.n19812 0.296
R15985 vp_p.n19817 vp_p.n19816 0.296
R15986 vp_p.n19827 vp_p.n19826 0.296
R15987 vp_p.n19831 vp_p.n19830 0.296
R15988 vp_p.n19841 vp_p.n19840 0.296
R15989 vp_p.n19845 vp_p.n19844 0.296
R15990 vp_p.n19855 vp_p.n19854 0.296
R15991 vp_p.n19859 vp_p.n19858 0.296
R15992 vp_p.n19869 vp_p.n19868 0.296
R15993 vp_p.n19873 vp_p.n19872 0.296
R15994 vp_p.n19883 vp_p.n19882 0.296
R15995 vp_p.n19887 vp_p.n19886 0.296
R15996 vp_p.n19897 vp_p.n19896 0.296
R15997 vp_p.n19901 vp_p.n19900 0.296
R15998 vp_p.n19911 vp_p.n19910 0.296
R15999 vp_p.n19915 vp_p.n19914 0.296
R16000 vp_p.n19925 vp_p.n19924 0.296
R16001 vp_p.n19929 vp_p.n19928 0.296
R16002 vp_p.n19939 vp_p.n19938 0.296
R16003 vp_p.n19943 vp_p.n19942 0.296
R16004 vp_p.n19953 vp_p.n19952 0.296
R16005 vp_p.n19957 vp_p.n19956 0.296
R16006 vp_p.n19967 vp_p.n19966 0.296
R16007 vp_p.n19971 vp_p.n19970 0.296
R16008 vp_p.n19981 vp_p.n19980 0.296
R16009 vp_p.n19985 vp_p.n19984 0.296
R16010 vp_p.n19995 vp_p.n19994 0.296
R16011 vp_p.n19999 vp_p.n19998 0.296
R16012 vp_p.n20009 vp_p.n20008 0.296
R16013 vp_p.n20013 vp_p.n20012 0.296
R16014 vp_p.n20023 vp_p.n20022 0.296
R16015 vp_p.n20027 vp_p.n20026 0.296
R16016 vp_p.n20037 vp_p.n20036 0.296
R16017 vp_p.n20041 vp_p.n20040 0.296
R16018 vp_p.n20051 vp_p.n20050 0.296
R16019 vp_p.n20055 vp_p.n20054 0.296
R16020 vp_p.n20065 vp_p.n20064 0.296
R16021 vp_p.n20069 vp_p.n20068 0.296
R16022 vp_p.n20079 vp_p.n20078 0.296
R16023 vp_p.n20083 vp_p.n20082 0.296
R16024 vp_p.n20093 vp_p.n20092 0.296
R16025 vp_p.n20097 vp_p.n20096 0.296
R16026 vp_p.n20107 vp_p.n20106 0.296
R16027 vp_p.n20111 vp_p.n20110 0.296
R16028 vp_p.n20121 vp_p.n20120 0.296
R16029 vp_p.n20125 vp_p.n20124 0.296
R16030 vp_p.n20135 vp_p.n20134 0.296
R16031 vp_p.n20139 vp_p.n20138 0.296
R16032 vp_p.n20143 vp_p.n20142 0.296
R16033 vp_p.n20153 vp_p.n20152 0.296
R16034 vp_p.n20158 vp_p.n20157 0.296
R16035 vp_p.n20163 vp_p.n20162 0.296
R16036 vp_p.n20168 vp_p.n20167 0.296
R16037 vp_p.n20173 vp_p.n20172 0.296
R16038 vp_p.n20178 vp_p.n20177 0.296
R16039 vp_p.n20183 vp_p.n20182 0.296
R16040 vp_p.n20188 vp_p.n20187 0.296
R16041 vp_p.n1889 vp_p.n1888 0.296
R16042 vp_p.n1894 vp_p.n1893 0.296
R16043 vp_p.n1904 vp_p.n1903 0.296
R16044 vp_p.n1908 vp_p.n1907 0.296
R16045 vp_p.n1918 vp_p.n1917 0.296
R16046 vp_p.n1922 vp_p.n1921 0.296
R16047 vp_p.n1932 vp_p.n1931 0.296
R16048 vp_p.n1936 vp_p.n1935 0.296
R16049 vp_p.n1946 vp_p.n1945 0.296
R16050 vp_p.n1950 vp_p.n1949 0.296
R16051 vp_p.n1960 vp_p.n1959 0.296
R16052 vp_p.n1964 vp_p.n1963 0.296
R16053 vp_p.n1974 vp_p.n1973 0.296
R16054 vp_p.n1978 vp_p.n1977 0.296
R16055 vp_p.n1988 vp_p.n1987 0.296
R16056 vp_p.n1992 vp_p.n1991 0.296
R16057 vp_p.n2002 vp_p.n2001 0.296
R16058 vp_p.n2006 vp_p.n2005 0.296
R16059 vp_p.n2016 vp_p.n2015 0.296
R16060 vp_p.n2020 vp_p.n2019 0.296
R16061 vp_p.n2030 vp_p.n2029 0.296
R16062 vp_p.n2034 vp_p.n2033 0.296
R16063 vp_p.n2044 vp_p.n2043 0.296
R16064 vp_p.n2048 vp_p.n2047 0.296
R16065 vp_p.n2058 vp_p.n2057 0.296
R16066 vp_p.n2062 vp_p.n2061 0.296
R16067 vp_p.n2072 vp_p.n2071 0.296
R16068 vp_p.n2076 vp_p.n2075 0.296
R16069 vp_p.n2086 vp_p.n2085 0.296
R16070 vp_p.n2090 vp_p.n2089 0.296
R16071 vp_p.n2100 vp_p.n2099 0.296
R16072 vp_p.n2104 vp_p.n2103 0.296
R16073 vp_p.n2114 vp_p.n2113 0.296
R16074 vp_p.n2118 vp_p.n2117 0.296
R16075 vp_p.n2128 vp_p.n2127 0.296
R16076 vp_p.n2132 vp_p.n2131 0.296
R16077 vp_p.n2142 vp_p.n2141 0.296
R16078 vp_p.n2146 vp_p.n2145 0.296
R16079 vp_p.n2156 vp_p.n2155 0.296
R16080 vp_p.n2160 vp_p.n2159 0.296
R16081 vp_p.n2170 vp_p.n2169 0.296
R16082 vp_p.n2174 vp_p.n2173 0.296
R16083 vp_p.n2184 vp_p.n2183 0.296
R16084 vp_p.n2188 vp_p.n2187 0.296
R16085 vp_p.n2198 vp_p.n2197 0.296
R16086 vp_p.n2202 vp_p.n2201 0.296
R16087 vp_p.n2212 vp_p.n2211 0.296
R16088 vp_p.n2216 vp_p.n2215 0.296
R16089 vp_p.n2226 vp_p.n2225 0.296
R16090 vp_p.n2230 vp_p.n2229 0.296
R16091 vp_p.n2240 vp_p.n2239 0.296
R16092 vp_p.n2244 vp_p.n2243 0.296
R16093 vp_p.n2254 vp_p.n2253 0.296
R16094 vp_p.n2258 vp_p.n2257 0.296
R16095 vp_p.n2268 vp_p.n2267 0.296
R16096 vp_p.n2272 vp_p.n2271 0.296
R16097 vp_p.n2282 vp_p.n2281 0.296
R16098 vp_p.n2286 vp_p.n2285 0.296
R16099 vp_p.n2296 vp_p.n2295 0.296
R16100 vp_p.n2300 vp_p.n2299 0.296
R16101 vp_p.n2310 vp_p.n2309 0.296
R16102 vp_p.n2314 vp_p.n2313 0.296
R16103 vp_p.n2324 vp_p.n2323 0.296
R16104 vp_p.n2328 vp_p.n2327 0.296
R16105 vp_p.n2338 vp_p.n2337 0.296
R16106 vp_p.n2342 vp_p.n2341 0.296
R16107 vp_p.n2352 vp_p.n2351 0.296
R16108 vp_p.n2356 vp_p.n2355 0.296
R16109 vp_p.n2366 vp_p.n2365 0.296
R16110 vp_p.n2370 vp_p.n2369 0.296
R16111 vp_p.n2380 vp_p.n2379 0.296
R16112 vp_p.n2384 vp_p.n2383 0.296
R16113 vp_p.n2394 vp_p.n2393 0.296
R16114 vp_p.n2398 vp_p.n2397 0.296
R16115 vp_p.n2408 vp_p.n2407 0.296
R16116 vp_p.n2412 vp_p.n2411 0.296
R16117 vp_p.n2422 vp_p.n2421 0.296
R16118 vp_p.n2426 vp_p.n2425 0.296
R16119 vp_p.n2436 vp_p.n2435 0.296
R16120 vp_p.n2440 vp_p.n2439 0.296
R16121 vp_p.n2450 vp_p.n2449 0.296
R16122 vp_p.n2454 vp_p.n2453 0.296
R16123 vp_p.n2464 vp_p.n2463 0.296
R16124 vp_p.n2468 vp_p.n2467 0.296
R16125 vp_p.n2478 vp_p.n2477 0.296
R16126 vp_p.n2482 vp_p.n2481 0.296
R16127 vp_p.n2492 vp_p.n2491 0.296
R16128 vp_p.n2496 vp_p.n2495 0.296
R16129 vp_p.n2506 vp_p.n2505 0.296
R16130 vp_p.n2510 vp_p.n2509 0.296
R16131 vp_p.n2520 vp_p.n2519 0.296
R16132 vp_p.n2524 vp_p.n2523 0.296
R16133 vp_p.n2534 vp_p.n2533 0.296
R16134 vp_p.n2538 vp_p.n2537 0.296
R16135 vp_p.n2548 vp_p.n2547 0.296
R16136 vp_p.n2552 vp_p.n2551 0.296
R16137 vp_p.n2562 vp_p.n2561 0.296
R16138 vp_p.n2566 vp_p.n2565 0.296
R16139 vp_p.n2576 vp_p.n2575 0.296
R16140 vp_p.n2580 vp_p.n2579 0.296
R16141 vp_p.n2590 vp_p.n2589 0.296
R16142 vp_p.n2594 vp_p.n2593 0.296
R16143 vp_p.n2604 vp_p.n2603 0.296
R16144 vp_p.n2608 vp_p.n2607 0.296
R16145 vp_p.n2618 vp_p.n2617 0.296
R16146 vp_p.n2622 vp_p.n2621 0.296
R16147 vp_p.n2632 vp_p.n2631 0.296
R16148 vp_p.n2636 vp_p.n2635 0.296
R16149 vp_p.n2646 vp_p.n2645 0.296
R16150 vp_p.n2650 vp_p.n2649 0.296
R16151 vp_p.n2660 vp_p.n2659 0.296
R16152 vp_p.n2664 vp_p.n2663 0.296
R16153 vp_p.n2674 vp_p.n2673 0.296
R16154 vp_p.n2678 vp_p.n2677 0.296
R16155 vp_p.n2688 vp_p.n2687 0.296
R16156 vp_p.n2692 vp_p.n2691 0.296
R16157 vp_p.n2702 vp_p.n2701 0.296
R16158 vp_p.n2706 vp_p.n2705 0.296
R16159 vp_p.n2716 vp_p.n2715 0.296
R16160 vp_p.n2720 vp_p.n2719 0.296
R16161 vp_p.n2730 vp_p.n2729 0.296
R16162 vp_p.n2734 vp_p.n2733 0.296
R16163 vp_p.n2744 vp_p.n2743 0.296
R16164 vp_p.n2748 vp_p.n2747 0.296
R16165 vp_p.n2758 vp_p.n2757 0.296
R16166 vp_p.n2762 vp_p.n2761 0.296
R16167 vp_p.n2772 vp_p.n2771 0.296
R16168 vp_p.n2776 vp_p.n2775 0.296
R16169 vp_p.n2786 vp_p.n2785 0.296
R16170 vp_p.n2790 vp_p.n2789 0.296
R16171 vp_p.n2800 vp_p.n2799 0.296
R16172 vp_p.n2804 vp_p.n2803 0.296
R16173 vp_p.n2814 vp_p.n2813 0.296
R16174 vp_p.n2818 vp_p.n2817 0.296
R16175 vp_p.n2828 vp_p.n2827 0.296
R16176 vp_p.n2832 vp_p.n2831 0.296
R16177 vp_p.n2842 vp_p.n2841 0.296
R16178 vp_p.n2846 vp_p.n2845 0.296
R16179 vp_p.n2856 vp_p.n2855 0.296
R16180 vp_p.n2860 vp_p.n2859 0.296
R16181 vp_p.n2870 vp_p.n2869 0.296
R16182 vp_p.n2874 vp_p.n2873 0.296
R16183 vp_p.n2884 vp_p.n2883 0.296
R16184 vp_p.n2889 vp_p.n2888 0.296
R16185 vp_p.n2894 vp_p.n2893 0.296
R16186 vp_p.n2899 vp_p.n2898 0.296
R16187 vp_p.n2904 vp_p.n2903 0.296
R16188 vp_p.n2909 vp_p.n2908 0.296
R16189 vp_p.n2914 vp_p.n2913 0.296
R16190 vp_p.n20593 vp_p.n20592 0.296
R16191 vp_p.n20598 vp_p.n20597 0.296
R16192 vp_p.n20608 vp_p.n20607 0.296
R16193 vp_p.n20612 vp_p.n20611 0.296
R16194 vp_p.n20622 vp_p.n20621 0.296
R16195 vp_p.n20626 vp_p.n20625 0.296
R16196 vp_p.n20636 vp_p.n20635 0.296
R16197 vp_p.n20640 vp_p.n20639 0.296
R16198 vp_p.n20650 vp_p.n20649 0.296
R16199 vp_p.n20654 vp_p.n20653 0.296
R16200 vp_p.n20664 vp_p.n20663 0.296
R16201 vp_p.n20668 vp_p.n20667 0.296
R16202 vp_p.n20678 vp_p.n20677 0.296
R16203 vp_p.n20682 vp_p.n20681 0.296
R16204 vp_p.n20692 vp_p.n20691 0.296
R16205 vp_p.n20696 vp_p.n20695 0.296
R16206 vp_p.n20706 vp_p.n20705 0.296
R16207 vp_p.n20710 vp_p.n20709 0.296
R16208 vp_p.n20720 vp_p.n20719 0.296
R16209 vp_p.n20724 vp_p.n20723 0.296
R16210 vp_p.n20734 vp_p.n20733 0.296
R16211 vp_p.n20738 vp_p.n20737 0.296
R16212 vp_p.n20748 vp_p.n20747 0.296
R16213 vp_p.n20752 vp_p.n20751 0.296
R16214 vp_p.n20762 vp_p.n20761 0.296
R16215 vp_p.n20766 vp_p.n20765 0.296
R16216 vp_p.n20776 vp_p.n20775 0.296
R16217 vp_p.n20780 vp_p.n20779 0.296
R16218 vp_p.n20790 vp_p.n20789 0.296
R16219 vp_p.n20794 vp_p.n20793 0.296
R16220 vp_p.n20804 vp_p.n20803 0.296
R16221 vp_p.n20808 vp_p.n20807 0.296
R16222 vp_p.n20818 vp_p.n20817 0.296
R16223 vp_p.n20822 vp_p.n20821 0.296
R16224 vp_p.n20832 vp_p.n20831 0.296
R16225 vp_p.n20836 vp_p.n20835 0.296
R16226 vp_p.n20846 vp_p.n20845 0.296
R16227 vp_p.n20850 vp_p.n20849 0.296
R16228 vp_p.n20860 vp_p.n20859 0.296
R16229 vp_p.n20864 vp_p.n20863 0.296
R16230 vp_p.n20874 vp_p.n20873 0.296
R16231 vp_p.n20878 vp_p.n20877 0.296
R16232 vp_p.n20888 vp_p.n20887 0.296
R16233 vp_p.n20892 vp_p.n20891 0.296
R16234 vp_p.n20902 vp_p.n20901 0.296
R16235 vp_p.n20906 vp_p.n20905 0.296
R16236 vp_p.n20916 vp_p.n20915 0.296
R16237 vp_p.n20920 vp_p.n20919 0.296
R16238 vp_p.n20930 vp_p.n20929 0.296
R16239 vp_p.n20934 vp_p.n20933 0.296
R16240 vp_p.n20944 vp_p.n20943 0.296
R16241 vp_p.n20948 vp_p.n20947 0.296
R16242 vp_p.n20958 vp_p.n20957 0.296
R16243 vp_p.n20962 vp_p.n20961 0.296
R16244 vp_p.n20972 vp_p.n20971 0.296
R16245 vp_p.n20976 vp_p.n20975 0.296
R16246 vp_p.n20986 vp_p.n20985 0.296
R16247 vp_p.n20990 vp_p.n20989 0.296
R16248 vp_p.n21000 vp_p.n20999 0.296
R16249 vp_p.n21004 vp_p.n21003 0.296
R16250 vp_p.n21014 vp_p.n21013 0.296
R16251 vp_p.n21018 vp_p.n21017 0.296
R16252 vp_p.n21028 vp_p.n21027 0.296
R16253 vp_p.n21032 vp_p.n21031 0.296
R16254 vp_p.n21042 vp_p.n21041 0.296
R16255 vp_p.n21046 vp_p.n21045 0.296
R16256 vp_p.n21056 vp_p.n21055 0.296
R16257 vp_p.n21060 vp_p.n21059 0.296
R16258 vp_p.n21070 vp_p.n21069 0.296
R16259 vp_p.n21074 vp_p.n21073 0.296
R16260 vp_p.n21084 vp_p.n21083 0.296
R16261 vp_p.n21088 vp_p.n21087 0.296
R16262 vp_p.n21098 vp_p.n21097 0.296
R16263 vp_p.n21102 vp_p.n21101 0.296
R16264 vp_p.n21112 vp_p.n21111 0.296
R16265 vp_p.n21116 vp_p.n21115 0.296
R16266 vp_p.n21126 vp_p.n21125 0.296
R16267 vp_p.n21130 vp_p.n21129 0.296
R16268 vp_p.n21140 vp_p.n21139 0.296
R16269 vp_p.n21144 vp_p.n21143 0.296
R16270 vp_p.n21154 vp_p.n21153 0.296
R16271 vp_p.n21158 vp_p.n21157 0.296
R16272 vp_p.n21168 vp_p.n21167 0.296
R16273 vp_p.n21172 vp_p.n21171 0.296
R16274 vp_p.n21182 vp_p.n21181 0.296
R16275 vp_p.n21186 vp_p.n21185 0.296
R16276 vp_p.n21196 vp_p.n21195 0.296
R16277 vp_p.n21200 vp_p.n21199 0.296
R16278 vp_p.n21210 vp_p.n21209 0.296
R16279 vp_p.n21214 vp_p.n21213 0.296
R16280 vp_p.n21224 vp_p.n21223 0.296
R16281 vp_p.n21228 vp_p.n21227 0.296
R16282 vp_p.n21238 vp_p.n21237 0.296
R16283 vp_p.n21242 vp_p.n21241 0.296
R16284 vp_p.n21252 vp_p.n21251 0.296
R16285 vp_p.n21256 vp_p.n21255 0.296
R16286 vp_p.n21266 vp_p.n21265 0.296
R16287 vp_p.n21270 vp_p.n21269 0.296
R16288 vp_p.n21280 vp_p.n21279 0.296
R16289 vp_p.n21284 vp_p.n21283 0.296
R16290 vp_p.n21294 vp_p.n21293 0.296
R16291 vp_p.n21298 vp_p.n21297 0.296
R16292 vp_p.n21308 vp_p.n21307 0.296
R16293 vp_p.n21312 vp_p.n21311 0.296
R16294 vp_p.n21322 vp_p.n21321 0.296
R16295 vp_p.n21326 vp_p.n21325 0.296
R16296 vp_p.n21336 vp_p.n21335 0.296
R16297 vp_p.n21340 vp_p.n21339 0.296
R16298 vp_p.n21350 vp_p.n21349 0.296
R16299 vp_p.n21354 vp_p.n21353 0.296
R16300 vp_p.n21364 vp_p.n21363 0.296
R16301 vp_p.n21368 vp_p.n21367 0.296
R16302 vp_p.n21378 vp_p.n21377 0.296
R16303 vp_p.n21382 vp_p.n21381 0.296
R16304 vp_p.n21392 vp_p.n21391 0.296
R16305 vp_p.n21396 vp_p.n21395 0.296
R16306 vp_p.n21406 vp_p.n21405 0.296
R16307 vp_p.n21410 vp_p.n21409 0.296
R16308 vp_p.n21420 vp_p.n21419 0.296
R16309 vp_p.n21424 vp_p.n21423 0.296
R16310 vp_p.n21434 vp_p.n21433 0.296
R16311 vp_p.n21438 vp_p.n21437 0.296
R16312 vp_p.n21448 vp_p.n21447 0.296
R16313 vp_p.n21452 vp_p.n21451 0.296
R16314 vp_p.n21462 vp_p.n21461 0.296
R16315 vp_p.n21466 vp_p.n21465 0.296
R16316 vp_p.n21476 vp_p.n21475 0.296
R16317 vp_p.n21480 vp_p.n21479 0.296
R16318 vp_p.n21490 vp_p.n21489 0.296
R16319 vp_p.n21494 vp_p.n21493 0.296
R16320 vp_p.n21504 vp_p.n21503 0.296
R16321 vp_p.n21508 vp_p.n21507 0.296
R16322 vp_p.n21518 vp_p.n21517 0.296
R16323 vp_p.n21522 vp_p.n21521 0.296
R16324 vp_p.n21532 vp_p.n21531 0.296
R16325 vp_p.n21536 vp_p.n21535 0.296
R16326 vp_p.n21546 vp_p.n21545 0.296
R16327 vp_p.n21550 vp_p.n21549 0.296
R16328 vp_p.n21560 vp_p.n21559 0.296
R16329 vp_p.n21564 vp_p.n21563 0.296
R16330 vp_p.n21574 vp_p.n21573 0.296
R16331 vp_p.n21578 vp_p.n21577 0.296
R16332 vp_p.n21582 vp_p.n21581 0.296
R16333 vp_p.n21592 vp_p.n21591 0.296
R16334 vp_p.n21597 vp_p.n21596 0.296
R16335 vp_p.n21602 vp_p.n21601 0.296
R16336 vp_p.n21607 vp_p.n21606 0.296
R16337 vp_p.n21612 vp_p.n21611 0.296
R16338 vp_p.n21617 vp_p.n21616 0.296
R16339 vp_p.n3314 vp_p.n3313 0.296
R16340 vp_p.n3319 vp_p.n3318 0.296
R16341 vp_p.n3329 vp_p.n3328 0.296
R16342 vp_p.n3333 vp_p.n3332 0.296
R16343 vp_p.n3343 vp_p.n3342 0.296
R16344 vp_p.n3347 vp_p.n3346 0.296
R16345 vp_p.n3357 vp_p.n3356 0.296
R16346 vp_p.n3361 vp_p.n3360 0.296
R16347 vp_p.n3371 vp_p.n3370 0.296
R16348 vp_p.n3375 vp_p.n3374 0.296
R16349 vp_p.n3385 vp_p.n3384 0.296
R16350 vp_p.n3389 vp_p.n3388 0.296
R16351 vp_p.n3399 vp_p.n3398 0.296
R16352 vp_p.n3403 vp_p.n3402 0.296
R16353 vp_p.n3413 vp_p.n3412 0.296
R16354 vp_p.n3417 vp_p.n3416 0.296
R16355 vp_p.n3427 vp_p.n3426 0.296
R16356 vp_p.n3431 vp_p.n3430 0.296
R16357 vp_p.n3441 vp_p.n3440 0.296
R16358 vp_p.n3445 vp_p.n3444 0.296
R16359 vp_p.n3455 vp_p.n3454 0.296
R16360 vp_p.n3459 vp_p.n3458 0.296
R16361 vp_p.n3469 vp_p.n3468 0.296
R16362 vp_p.n3473 vp_p.n3472 0.296
R16363 vp_p.n3483 vp_p.n3482 0.296
R16364 vp_p.n3487 vp_p.n3486 0.296
R16365 vp_p.n3497 vp_p.n3496 0.296
R16366 vp_p.n3501 vp_p.n3500 0.296
R16367 vp_p.n3511 vp_p.n3510 0.296
R16368 vp_p.n3515 vp_p.n3514 0.296
R16369 vp_p.n3525 vp_p.n3524 0.296
R16370 vp_p.n3529 vp_p.n3528 0.296
R16371 vp_p.n3539 vp_p.n3538 0.296
R16372 vp_p.n3543 vp_p.n3542 0.296
R16373 vp_p.n3553 vp_p.n3552 0.296
R16374 vp_p.n3557 vp_p.n3556 0.296
R16375 vp_p.n3567 vp_p.n3566 0.296
R16376 vp_p.n3571 vp_p.n3570 0.296
R16377 vp_p.n3581 vp_p.n3580 0.296
R16378 vp_p.n3585 vp_p.n3584 0.296
R16379 vp_p.n3595 vp_p.n3594 0.296
R16380 vp_p.n3599 vp_p.n3598 0.296
R16381 vp_p.n3609 vp_p.n3608 0.296
R16382 vp_p.n3613 vp_p.n3612 0.296
R16383 vp_p.n3623 vp_p.n3622 0.296
R16384 vp_p.n3627 vp_p.n3626 0.296
R16385 vp_p.n3637 vp_p.n3636 0.296
R16386 vp_p.n3641 vp_p.n3640 0.296
R16387 vp_p.n3651 vp_p.n3650 0.296
R16388 vp_p.n3655 vp_p.n3654 0.296
R16389 vp_p.n3665 vp_p.n3664 0.296
R16390 vp_p.n3669 vp_p.n3668 0.296
R16391 vp_p.n3679 vp_p.n3678 0.296
R16392 vp_p.n3683 vp_p.n3682 0.296
R16393 vp_p.n3693 vp_p.n3692 0.296
R16394 vp_p.n3697 vp_p.n3696 0.296
R16395 vp_p.n3707 vp_p.n3706 0.296
R16396 vp_p.n3711 vp_p.n3710 0.296
R16397 vp_p.n3721 vp_p.n3720 0.296
R16398 vp_p.n3725 vp_p.n3724 0.296
R16399 vp_p.n3735 vp_p.n3734 0.296
R16400 vp_p.n3739 vp_p.n3738 0.296
R16401 vp_p.n3749 vp_p.n3748 0.296
R16402 vp_p.n3753 vp_p.n3752 0.296
R16403 vp_p.n3763 vp_p.n3762 0.296
R16404 vp_p.n3767 vp_p.n3766 0.296
R16405 vp_p.n3777 vp_p.n3776 0.296
R16406 vp_p.n3781 vp_p.n3780 0.296
R16407 vp_p.n3791 vp_p.n3790 0.296
R16408 vp_p.n3795 vp_p.n3794 0.296
R16409 vp_p.n3805 vp_p.n3804 0.296
R16410 vp_p.n3809 vp_p.n3808 0.296
R16411 vp_p.n3819 vp_p.n3818 0.296
R16412 vp_p.n3823 vp_p.n3822 0.296
R16413 vp_p.n3833 vp_p.n3832 0.296
R16414 vp_p.n3837 vp_p.n3836 0.296
R16415 vp_p.n3847 vp_p.n3846 0.296
R16416 vp_p.n3851 vp_p.n3850 0.296
R16417 vp_p.n3861 vp_p.n3860 0.296
R16418 vp_p.n3865 vp_p.n3864 0.296
R16419 vp_p.n3875 vp_p.n3874 0.296
R16420 vp_p.n3879 vp_p.n3878 0.296
R16421 vp_p.n3889 vp_p.n3888 0.296
R16422 vp_p.n3893 vp_p.n3892 0.296
R16423 vp_p.n3903 vp_p.n3902 0.296
R16424 vp_p.n3907 vp_p.n3906 0.296
R16425 vp_p.n3917 vp_p.n3916 0.296
R16426 vp_p.n3921 vp_p.n3920 0.296
R16427 vp_p.n3931 vp_p.n3930 0.296
R16428 vp_p.n3935 vp_p.n3934 0.296
R16429 vp_p.n3945 vp_p.n3944 0.296
R16430 vp_p.n3949 vp_p.n3948 0.296
R16431 vp_p.n3959 vp_p.n3958 0.296
R16432 vp_p.n3963 vp_p.n3962 0.296
R16433 vp_p.n3973 vp_p.n3972 0.296
R16434 vp_p.n3977 vp_p.n3976 0.296
R16435 vp_p.n3987 vp_p.n3986 0.296
R16436 vp_p.n3991 vp_p.n3990 0.296
R16437 vp_p.n4001 vp_p.n4000 0.296
R16438 vp_p.n4005 vp_p.n4004 0.296
R16439 vp_p.n4015 vp_p.n4014 0.296
R16440 vp_p.n4019 vp_p.n4018 0.296
R16441 vp_p.n4029 vp_p.n4028 0.296
R16442 vp_p.n4033 vp_p.n4032 0.296
R16443 vp_p.n4043 vp_p.n4042 0.296
R16444 vp_p.n4047 vp_p.n4046 0.296
R16445 vp_p.n4057 vp_p.n4056 0.296
R16446 vp_p.n4061 vp_p.n4060 0.296
R16447 vp_p.n4071 vp_p.n4070 0.296
R16448 vp_p.n4075 vp_p.n4074 0.296
R16449 vp_p.n4085 vp_p.n4084 0.296
R16450 vp_p.n4089 vp_p.n4088 0.296
R16451 vp_p.n4099 vp_p.n4098 0.296
R16452 vp_p.n4103 vp_p.n4102 0.296
R16453 vp_p.n4113 vp_p.n4112 0.296
R16454 vp_p.n4117 vp_p.n4116 0.296
R16455 vp_p.n4127 vp_p.n4126 0.296
R16456 vp_p.n4131 vp_p.n4130 0.296
R16457 vp_p.n4141 vp_p.n4140 0.296
R16458 vp_p.n4145 vp_p.n4144 0.296
R16459 vp_p.n4155 vp_p.n4154 0.296
R16460 vp_p.n4159 vp_p.n4158 0.296
R16461 vp_p.n4169 vp_p.n4168 0.296
R16462 vp_p.n4173 vp_p.n4172 0.296
R16463 vp_p.n4183 vp_p.n4182 0.296
R16464 vp_p.n4187 vp_p.n4186 0.296
R16465 vp_p.n4197 vp_p.n4196 0.296
R16466 vp_p.n4201 vp_p.n4200 0.296
R16467 vp_p.n4211 vp_p.n4210 0.296
R16468 vp_p.n4215 vp_p.n4214 0.296
R16469 vp_p.n4225 vp_p.n4224 0.296
R16470 vp_p.n4229 vp_p.n4228 0.296
R16471 vp_p.n4239 vp_p.n4238 0.296
R16472 vp_p.n4243 vp_p.n4242 0.296
R16473 vp_p.n4253 vp_p.n4252 0.296
R16474 vp_p.n4257 vp_p.n4256 0.296
R16475 vp_p.n4267 vp_p.n4266 0.296
R16476 vp_p.n4271 vp_p.n4270 0.296
R16477 vp_p.n4281 vp_p.n4280 0.296
R16478 vp_p.n4285 vp_p.n4284 0.296
R16479 vp_p.n4295 vp_p.n4294 0.296
R16480 vp_p.n4299 vp_p.n4298 0.296
R16481 vp_p.n4309 vp_p.n4308 0.296
R16482 vp_p.n4313 vp_p.n4312 0.296
R16483 vp_p.n4323 vp_p.n4322 0.296
R16484 vp_p.n4328 vp_p.n4327 0.296
R16485 vp_p.n4333 vp_p.n4332 0.296
R16486 vp_p.n4338 vp_p.n4337 0.296
R16487 vp_p.n4343 vp_p.n4342 0.296
R16488 vp_p.n22017 vp_p.n22016 0.296
R16489 vp_p.n22022 vp_p.n22021 0.296
R16490 vp_p.n22032 vp_p.n22031 0.296
R16491 vp_p.n22036 vp_p.n22035 0.296
R16492 vp_p.n22046 vp_p.n22045 0.296
R16493 vp_p.n22050 vp_p.n22049 0.296
R16494 vp_p.n22060 vp_p.n22059 0.296
R16495 vp_p.n22064 vp_p.n22063 0.296
R16496 vp_p.n22074 vp_p.n22073 0.296
R16497 vp_p.n22078 vp_p.n22077 0.296
R16498 vp_p.n22088 vp_p.n22087 0.296
R16499 vp_p.n22092 vp_p.n22091 0.296
R16500 vp_p.n22102 vp_p.n22101 0.296
R16501 vp_p.n22106 vp_p.n22105 0.296
R16502 vp_p.n22116 vp_p.n22115 0.296
R16503 vp_p.n22120 vp_p.n22119 0.296
R16504 vp_p.n22130 vp_p.n22129 0.296
R16505 vp_p.n22134 vp_p.n22133 0.296
R16506 vp_p.n22144 vp_p.n22143 0.296
R16507 vp_p.n22148 vp_p.n22147 0.296
R16508 vp_p.n22158 vp_p.n22157 0.296
R16509 vp_p.n22162 vp_p.n22161 0.296
R16510 vp_p.n22172 vp_p.n22171 0.296
R16511 vp_p.n22176 vp_p.n22175 0.296
R16512 vp_p.n22186 vp_p.n22185 0.296
R16513 vp_p.n22190 vp_p.n22189 0.296
R16514 vp_p.n22200 vp_p.n22199 0.296
R16515 vp_p.n22204 vp_p.n22203 0.296
R16516 vp_p.n22214 vp_p.n22213 0.296
R16517 vp_p.n22218 vp_p.n22217 0.296
R16518 vp_p.n22228 vp_p.n22227 0.296
R16519 vp_p.n22232 vp_p.n22231 0.296
R16520 vp_p.n22242 vp_p.n22241 0.296
R16521 vp_p.n22246 vp_p.n22245 0.296
R16522 vp_p.n22256 vp_p.n22255 0.296
R16523 vp_p.n22260 vp_p.n22259 0.296
R16524 vp_p.n22270 vp_p.n22269 0.296
R16525 vp_p.n22274 vp_p.n22273 0.296
R16526 vp_p.n22284 vp_p.n22283 0.296
R16527 vp_p.n22288 vp_p.n22287 0.296
R16528 vp_p.n22298 vp_p.n22297 0.296
R16529 vp_p.n22302 vp_p.n22301 0.296
R16530 vp_p.n22312 vp_p.n22311 0.296
R16531 vp_p.n22316 vp_p.n22315 0.296
R16532 vp_p.n22326 vp_p.n22325 0.296
R16533 vp_p.n22330 vp_p.n22329 0.296
R16534 vp_p.n22340 vp_p.n22339 0.296
R16535 vp_p.n22344 vp_p.n22343 0.296
R16536 vp_p.n22354 vp_p.n22353 0.296
R16537 vp_p.n22358 vp_p.n22357 0.296
R16538 vp_p.n22368 vp_p.n22367 0.296
R16539 vp_p.n22372 vp_p.n22371 0.296
R16540 vp_p.n22382 vp_p.n22381 0.296
R16541 vp_p.n22386 vp_p.n22385 0.296
R16542 vp_p.n22396 vp_p.n22395 0.296
R16543 vp_p.n22400 vp_p.n22399 0.296
R16544 vp_p.n22410 vp_p.n22409 0.296
R16545 vp_p.n22414 vp_p.n22413 0.296
R16546 vp_p.n22424 vp_p.n22423 0.296
R16547 vp_p.n22428 vp_p.n22427 0.296
R16548 vp_p.n22438 vp_p.n22437 0.296
R16549 vp_p.n22442 vp_p.n22441 0.296
R16550 vp_p.n22452 vp_p.n22451 0.296
R16551 vp_p.n22456 vp_p.n22455 0.296
R16552 vp_p.n22466 vp_p.n22465 0.296
R16553 vp_p.n22470 vp_p.n22469 0.296
R16554 vp_p.n22480 vp_p.n22479 0.296
R16555 vp_p.n22484 vp_p.n22483 0.296
R16556 vp_p.n22494 vp_p.n22493 0.296
R16557 vp_p.n22498 vp_p.n22497 0.296
R16558 vp_p.n22508 vp_p.n22507 0.296
R16559 vp_p.n22512 vp_p.n22511 0.296
R16560 vp_p.n22522 vp_p.n22521 0.296
R16561 vp_p.n22526 vp_p.n22525 0.296
R16562 vp_p.n22536 vp_p.n22535 0.296
R16563 vp_p.n22540 vp_p.n22539 0.296
R16564 vp_p.n22550 vp_p.n22549 0.296
R16565 vp_p.n22554 vp_p.n22553 0.296
R16566 vp_p.n22564 vp_p.n22563 0.296
R16567 vp_p.n22568 vp_p.n22567 0.296
R16568 vp_p.n22578 vp_p.n22577 0.296
R16569 vp_p.n22582 vp_p.n22581 0.296
R16570 vp_p.n22592 vp_p.n22591 0.296
R16571 vp_p.n22596 vp_p.n22595 0.296
R16572 vp_p.n22606 vp_p.n22605 0.296
R16573 vp_p.n22610 vp_p.n22609 0.296
R16574 vp_p.n22620 vp_p.n22619 0.296
R16575 vp_p.n22624 vp_p.n22623 0.296
R16576 vp_p.n22634 vp_p.n22633 0.296
R16577 vp_p.n22638 vp_p.n22637 0.296
R16578 vp_p.n22648 vp_p.n22647 0.296
R16579 vp_p.n22652 vp_p.n22651 0.296
R16580 vp_p.n22662 vp_p.n22661 0.296
R16581 vp_p.n22666 vp_p.n22665 0.296
R16582 vp_p.n22676 vp_p.n22675 0.296
R16583 vp_p.n22680 vp_p.n22679 0.296
R16584 vp_p.n22690 vp_p.n22689 0.296
R16585 vp_p.n22694 vp_p.n22693 0.296
R16586 vp_p.n22704 vp_p.n22703 0.296
R16587 vp_p.n22708 vp_p.n22707 0.296
R16588 vp_p.n22718 vp_p.n22717 0.296
R16589 vp_p.n22722 vp_p.n22721 0.296
R16590 vp_p.n22732 vp_p.n22731 0.296
R16591 vp_p.n22736 vp_p.n22735 0.296
R16592 vp_p.n22746 vp_p.n22745 0.296
R16593 vp_p.n22750 vp_p.n22749 0.296
R16594 vp_p.n22760 vp_p.n22759 0.296
R16595 vp_p.n22764 vp_p.n22763 0.296
R16596 vp_p.n22774 vp_p.n22773 0.296
R16597 vp_p.n22778 vp_p.n22777 0.296
R16598 vp_p.n22788 vp_p.n22787 0.296
R16599 vp_p.n22792 vp_p.n22791 0.296
R16600 vp_p.n22802 vp_p.n22801 0.296
R16601 vp_p.n22806 vp_p.n22805 0.296
R16602 vp_p.n22816 vp_p.n22815 0.296
R16603 vp_p.n22820 vp_p.n22819 0.296
R16604 vp_p.n22830 vp_p.n22829 0.296
R16605 vp_p.n22834 vp_p.n22833 0.296
R16606 vp_p.n22844 vp_p.n22843 0.296
R16607 vp_p.n22848 vp_p.n22847 0.296
R16608 vp_p.n22858 vp_p.n22857 0.296
R16609 vp_p.n22862 vp_p.n22861 0.296
R16610 vp_p.n22872 vp_p.n22871 0.296
R16611 vp_p.n22876 vp_p.n22875 0.296
R16612 vp_p.n22886 vp_p.n22885 0.296
R16613 vp_p.n22890 vp_p.n22889 0.296
R16614 vp_p.n22900 vp_p.n22899 0.296
R16615 vp_p.n22904 vp_p.n22903 0.296
R16616 vp_p.n22914 vp_p.n22913 0.296
R16617 vp_p.n22918 vp_p.n22917 0.296
R16618 vp_p.n22928 vp_p.n22927 0.296
R16619 vp_p.n22932 vp_p.n22931 0.296
R16620 vp_p.n22942 vp_p.n22941 0.296
R16621 vp_p.n22946 vp_p.n22945 0.296
R16622 vp_p.n22956 vp_p.n22955 0.296
R16623 vp_p.n22960 vp_p.n22959 0.296
R16624 vp_p.n22970 vp_p.n22969 0.296
R16625 vp_p.n22974 vp_p.n22973 0.296
R16626 vp_p.n22984 vp_p.n22983 0.296
R16627 vp_p.n22988 vp_p.n22987 0.296
R16628 vp_p.n22998 vp_p.n22997 0.296
R16629 vp_p.n23002 vp_p.n23001 0.296
R16630 vp_p.n23012 vp_p.n23011 0.296
R16631 vp_p.n23016 vp_p.n23015 0.296
R16632 vp_p.n23020 vp_p.n23019 0.296
R16633 vp_p.n23030 vp_p.n23029 0.296
R16634 vp_p.n23035 vp_p.n23034 0.296
R16635 vp_p.n23040 vp_p.n23039 0.296
R16636 vp_p.n23045 vp_p.n23044 0.296
R16637 vp_p.n4738 vp_p.n4737 0.296
R16638 vp_p.n4743 vp_p.n4742 0.296
R16639 vp_p.n4753 vp_p.n4752 0.296
R16640 vp_p.n4757 vp_p.n4756 0.296
R16641 vp_p.n4767 vp_p.n4766 0.296
R16642 vp_p.n4771 vp_p.n4770 0.296
R16643 vp_p.n4781 vp_p.n4780 0.296
R16644 vp_p.n4785 vp_p.n4784 0.296
R16645 vp_p.n4795 vp_p.n4794 0.296
R16646 vp_p.n4799 vp_p.n4798 0.296
R16647 vp_p.n4809 vp_p.n4808 0.296
R16648 vp_p.n4813 vp_p.n4812 0.296
R16649 vp_p.n4823 vp_p.n4822 0.296
R16650 vp_p.n4827 vp_p.n4826 0.296
R16651 vp_p.n4837 vp_p.n4836 0.296
R16652 vp_p.n4841 vp_p.n4840 0.296
R16653 vp_p.n4851 vp_p.n4850 0.296
R16654 vp_p.n4855 vp_p.n4854 0.296
R16655 vp_p.n4865 vp_p.n4864 0.296
R16656 vp_p.n4869 vp_p.n4868 0.296
R16657 vp_p.n4879 vp_p.n4878 0.296
R16658 vp_p.n4883 vp_p.n4882 0.296
R16659 vp_p.n4893 vp_p.n4892 0.296
R16660 vp_p.n4897 vp_p.n4896 0.296
R16661 vp_p.n4907 vp_p.n4906 0.296
R16662 vp_p.n4911 vp_p.n4910 0.296
R16663 vp_p.n4921 vp_p.n4920 0.296
R16664 vp_p.n4925 vp_p.n4924 0.296
R16665 vp_p.n4935 vp_p.n4934 0.296
R16666 vp_p.n4939 vp_p.n4938 0.296
R16667 vp_p.n4949 vp_p.n4948 0.296
R16668 vp_p.n4953 vp_p.n4952 0.296
R16669 vp_p.n4963 vp_p.n4962 0.296
R16670 vp_p.n4967 vp_p.n4966 0.296
R16671 vp_p.n4977 vp_p.n4976 0.296
R16672 vp_p.n4981 vp_p.n4980 0.296
R16673 vp_p.n4991 vp_p.n4990 0.296
R16674 vp_p.n4995 vp_p.n4994 0.296
R16675 vp_p.n5005 vp_p.n5004 0.296
R16676 vp_p.n5009 vp_p.n5008 0.296
R16677 vp_p.n5019 vp_p.n5018 0.296
R16678 vp_p.n5023 vp_p.n5022 0.296
R16679 vp_p.n5033 vp_p.n5032 0.296
R16680 vp_p.n5037 vp_p.n5036 0.296
R16681 vp_p.n5047 vp_p.n5046 0.296
R16682 vp_p.n5051 vp_p.n5050 0.296
R16683 vp_p.n5061 vp_p.n5060 0.296
R16684 vp_p.n5065 vp_p.n5064 0.296
R16685 vp_p.n5075 vp_p.n5074 0.296
R16686 vp_p.n5079 vp_p.n5078 0.296
R16687 vp_p.n5089 vp_p.n5088 0.296
R16688 vp_p.n5093 vp_p.n5092 0.296
R16689 vp_p.n5103 vp_p.n5102 0.296
R16690 vp_p.n5107 vp_p.n5106 0.296
R16691 vp_p.n5117 vp_p.n5116 0.296
R16692 vp_p.n5121 vp_p.n5120 0.296
R16693 vp_p.n5131 vp_p.n5130 0.296
R16694 vp_p.n5135 vp_p.n5134 0.296
R16695 vp_p.n5145 vp_p.n5144 0.296
R16696 vp_p.n5149 vp_p.n5148 0.296
R16697 vp_p.n5159 vp_p.n5158 0.296
R16698 vp_p.n5163 vp_p.n5162 0.296
R16699 vp_p.n5173 vp_p.n5172 0.296
R16700 vp_p.n5177 vp_p.n5176 0.296
R16701 vp_p.n5187 vp_p.n5186 0.296
R16702 vp_p.n5191 vp_p.n5190 0.296
R16703 vp_p.n5201 vp_p.n5200 0.296
R16704 vp_p.n5205 vp_p.n5204 0.296
R16705 vp_p.n5215 vp_p.n5214 0.296
R16706 vp_p.n5219 vp_p.n5218 0.296
R16707 vp_p.n5229 vp_p.n5228 0.296
R16708 vp_p.n5233 vp_p.n5232 0.296
R16709 vp_p.n5243 vp_p.n5242 0.296
R16710 vp_p.n5247 vp_p.n5246 0.296
R16711 vp_p.n5257 vp_p.n5256 0.296
R16712 vp_p.n5261 vp_p.n5260 0.296
R16713 vp_p.n5271 vp_p.n5270 0.296
R16714 vp_p.n5275 vp_p.n5274 0.296
R16715 vp_p.n5285 vp_p.n5284 0.296
R16716 vp_p.n5289 vp_p.n5288 0.296
R16717 vp_p.n5299 vp_p.n5298 0.296
R16718 vp_p.n5303 vp_p.n5302 0.296
R16719 vp_p.n5313 vp_p.n5312 0.296
R16720 vp_p.n5317 vp_p.n5316 0.296
R16721 vp_p.n5327 vp_p.n5326 0.296
R16722 vp_p.n5331 vp_p.n5330 0.296
R16723 vp_p.n5341 vp_p.n5340 0.296
R16724 vp_p.n5345 vp_p.n5344 0.296
R16725 vp_p.n5355 vp_p.n5354 0.296
R16726 vp_p.n5359 vp_p.n5358 0.296
R16727 vp_p.n5369 vp_p.n5368 0.296
R16728 vp_p.n5373 vp_p.n5372 0.296
R16729 vp_p.n5383 vp_p.n5382 0.296
R16730 vp_p.n5387 vp_p.n5386 0.296
R16731 vp_p.n5397 vp_p.n5396 0.296
R16732 vp_p.n5401 vp_p.n5400 0.296
R16733 vp_p.n5411 vp_p.n5410 0.296
R16734 vp_p.n5415 vp_p.n5414 0.296
R16735 vp_p.n5425 vp_p.n5424 0.296
R16736 vp_p.n5429 vp_p.n5428 0.296
R16737 vp_p.n5439 vp_p.n5438 0.296
R16738 vp_p.n5443 vp_p.n5442 0.296
R16739 vp_p.n5453 vp_p.n5452 0.296
R16740 vp_p.n5457 vp_p.n5456 0.296
R16741 vp_p.n5467 vp_p.n5466 0.296
R16742 vp_p.n5471 vp_p.n5470 0.296
R16743 vp_p.n5481 vp_p.n5480 0.296
R16744 vp_p.n5485 vp_p.n5484 0.296
R16745 vp_p.n5495 vp_p.n5494 0.296
R16746 vp_p.n5499 vp_p.n5498 0.296
R16747 vp_p.n5509 vp_p.n5508 0.296
R16748 vp_p.n5513 vp_p.n5512 0.296
R16749 vp_p.n5523 vp_p.n5522 0.296
R16750 vp_p.n5527 vp_p.n5526 0.296
R16751 vp_p.n5537 vp_p.n5536 0.296
R16752 vp_p.n5541 vp_p.n5540 0.296
R16753 vp_p.n5551 vp_p.n5550 0.296
R16754 vp_p.n5555 vp_p.n5554 0.296
R16755 vp_p.n5565 vp_p.n5564 0.296
R16756 vp_p.n5569 vp_p.n5568 0.296
R16757 vp_p.n5579 vp_p.n5578 0.296
R16758 vp_p.n5583 vp_p.n5582 0.296
R16759 vp_p.n5593 vp_p.n5592 0.296
R16760 vp_p.n5597 vp_p.n5596 0.296
R16761 vp_p.n5607 vp_p.n5606 0.296
R16762 vp_p.n5611 vp_p.n5610 0.296
R16763 vp_p.n5621 vp_p.n5620 0.296
R16764 vp_p.n5625 vp_p.n5624 0.296
R16765 vp_p.n5635 vp_p.n5634 0.296
R16766 vp_p.n5639 vp_p.n5638 0.296
R16767 vp_p.n5649 vp_p.n5648 0.296
R16768 vp_p.n5653 vp_p.n5652 0.296
R16769 vp_p.n5663 vp_p.n5662 0.296
R16770 vp_p.n5667 vp_p.n5666 0.296
R16771 vp_p.n5677 vp_p.n5676 0.296
R16772 vp_p.n5681 vp_p.n5680 0.296
R16773 vp_p.n5691 vp_p.n5690 0.296
R16774 vp_p.n5695 vp_p.n5694 0.296
R16775 vp_p.n5705 vp_p.n5704 0.296
R16776 vp_p.n5709 vp_p.n5708 0.296
R16777 vp_p.n5719 vp_p.n5718 0.296
R16778 vp_p.n5723 vp_p.n5722 0.296
R16779 vp_p.n5733 vp_p.n5732 0.296
R16780 vp_p.n5737 vp_p.n5736 0.296
R16781 vp_p.n5747 vp_p.n5746 0.296
R16782 vp_p.n5751 vp_p.n5750 0.296
R16783 vp_p.n5761 vp_p.n5760 0.296
R16784 vp_p.n5766 vp_p.n5765 0.296
R16785 vp_p.n5771 vp_p.n5770 0.296
R16786 vp_p.n23440 vp_p.n23439 0.296
R16787 vp_p.n23445 vp_p.n23444 0.296
R16788 vp_p.n23455 vp_p.n23454 0.296
R16789 vp_p.n23459 vp_p.n23458 0.296
R16790 vp_p.n23469 vp_p.n23468 0.296
R16791 vp_p.n23473 vp_p.n23472 0.296
R16792 vp_p.n23483 vp_p.n23482 0.296
R16793 vp_p.n23487 vp_p.n23486 0.296
R16794 vp_p.n23497 vp_p.n23496 0.296
R16795 vp_p.n23501 vp_p.n23500 0.296
R16796 vp_p.n23511 vp_p.n23510 0.296
R16797 vp_p.n23515 vp_p.n23514 0.296
R16798 vp_p.n23525 vp_p.n23524 0.296
R16799 vp_p.n23529 vp_p.n23528 0.296
R16800 vp_p.n23539 vp_p.n23538 0.296
R16801 vp_p.n23543 vp_p.n23542 0.296
R16802 vp_p.n23553 vp_p.n23552 0.296
R16803 vp_p.n23557 vp_p.n23556 0.296
R16804 vp_p.n23567 vp_p.n23566 0.296
R16805 vp_p.n23571 vp_p.n23570 0.296
R16806 vp_p.n23581 vp_p.n23580 0.296
R16807 vp_p.n23585 vp_p.n23584 0.296
R16808 vp_p.n23595 vp_p.n23594 0.296
R16809 vp_p.n23599 vp_p.n23598 0.296
R16810 vp_p.n23609 vp_p.n23608 0.296
R16811 vp_p.n23613 vp_p.n23612 0.296
R16812 vp_p.n23623 vp_p.n23622 0.296
R16813 vp_p.n23627 vp_p.n23626 0.296
R16814 vp_p.n23637 vp_p.n23636 0.296
R16815 vp_p.n23641 vp_p.n23640 0.296
R16816 vp_p.n23651 vp_p.n23650 0.296
R16817 vp_p.n23655 vp_p.n23654 0.296
R16818 vp_p.n23665 vp_p.n23664 0.296
R16819 vp_p.n23669 vp_p.n23668 0.296
R16820 vp_p.n23679 vp_p.n23678 0.296
R16821 vp_p.n23683 vp_p.n23682 0.296
R16822 vp_p.n23693 vp_p.n23692 0.296
R16823 vp_p.n23697 vp_p.n23696 0.296
R16824 vp_p.n23707 vp_p.n23706 0.296
R16825 vp_p.n23711 vp_p.n23710 0.296
R16826 vp_p.n23721 vp_p.n23720 0.296
R16827 vp_p.n23725 vp_p.n23724 0.296
R16828 vp_p.n23735 vp_p.n23734 0.296
R16829 vp_p.n23739 vp_p.n23738 0.296
R16830 vp_p.n23749 vp_p.n23748 0.296
R16831 vp_p.n23753 vp_p.n23752 0.296
R16832 vp_p.n23763 vp_p.n23762 0.296
R16833 vp_p.n23767 vp_p.n23766 0.296
R16834 vp_p.n23777 vp_p.n23776 0.296
R16835 vp_p.n23781 vp_p.n23780 0.296
R16836 vp_p.n23791 vp_p.n23790 0.296
R16837 vp_p.n23795 vp_p.n23794 0.296
R16838 vp_p.n23805 vp_p.n23804 0.296
R16839 vp_p.n23809 vp_p.n23808 0.296
R16840 vp_p.n23819 vp_p.n23818 0.296
R16841 vp_p.n23823 vp_p.n23822 0.296
R16842 vp_p.n23833 vp_p.n23832 0.296
R16843 vp_p.n23837 vp_p.n23836 0.296
R16844 vp_p.n23847 vp_p.n23846 0.296
R16845 vp_p.n23851 vp_p.n23850 0.296
R16846 vp_p.n23861 vp_p.n23860 0.296
R16847 vp_p.n23865 vp_p.n23864 0.296
R16848 vp_p.n23875 vp_p.n23874 0.296
R16849 vp_p.n23879 vp_p.n23878 0.296
R16850 vp_p.n23889 vp_p.n23888 0.296
R16851 vp_p.n23893 vp_p.n23892 0.296
R16852 vp_p.n23903 vp_p.n23902 0.296
R16853 vp_p.n23907 vp_p.n23906 0.296
R16854 vp_p.n23917 vp_p.n23916 0.296
R16855 vp_p.n23921 vp_p.n23920 0.296
R16856 vp_p.n23931 vp_p.n23930 0.296
R16857 vp_p.n23935 vp_p.n23934 0.296
R16858 vp_p.n23945 vp_p.n23944 0.296
R16859 vp_p.n23949 vp_p.n23948 0.296
R16860 vp_p.n23959 vp_p.n23958 0.296
R16861 vp_p.n23963 vp_p.n23962 0.296
R16862 vp_p.n23973 vp_p.n23972 0.296
R16863 vp_p.n23977 vp_p.n23976 0.296
R16864 vp_p.n23987 vp_p.n23986 0.296
R16865 vp_p.n23991 vp_p.n23990 0.296
R16866 vp_p.n24001 vp_p.n24000 0.296
R16867 vp_p.n24005 vp_p.n24004 0.296
R16868 vp_p.n24015 vp_p.n24014 0.296
R16869 vp_p.n24019 vp_p.n24018 0.296
R16870 vp_p.n24029 vp_p.n24028 0.296
R16871 vp_p.n24033 vp_p.n24032 0.296
R16872 vp_p.n24043 vp_p.n24042 0.296
R16873 vp_p.n24047 vp_p.n24046 0.296
R16874 vp_p.n24057 vp_p.n24056 0.296
R16875 vp_p.n24061 vp_p.n24060 0.296
R16876 vp_p.n24071 vp_p.n24070 0.296
R16877 vp_p.n24075 vp_p.n24074 0.296
R16878 vp_p.n24085 vp_p.n24084 0.296
R16879 vp_p.n24089 vp_p.n24088 0.296
R16880 vp_p.n24099 vp_p.n24098 0.296
R16881 vp_p.n24103 vp_p.n24102 0.296
R16882 vp_p.n24113 vp_p.n24112 0.296
R16883 vp_p.n24117 vp_p.n24116 0.296
R16884 vp_p.n24127 vp_p.n24126 0.296
R16885 vp_p.n24131 vp_p.n24130 0.296
R16886 vp_p.n24141 vp_p.n24140 0.296
R16887 vp_p.n24145 vp_p.n24144 0.296
R16888 vp_p.n24155 vp_p.n24154 0.296
R16889 vp_p.n24159 vp_p.n24158 0.296
R16890 vp_p.n24169 vp_p.n24168 0.296
R16891 vp_p.n24173 vp_p.n24172 0.296
R16892 vp_p.n24183 vp_p.n24182 0.296
R16893 vp_p.n24187 vp_p.n24186 0.296
R16894 vp_p.n24197 vp_p.n24196 0.296
R16895 vp_p.n24201 vp_p.n24200 0.296
R16896 vp_p.n24211 vp_p.n24210 0.296
R16897 vp_p.n24215 vp_p.n24214 0.296
R16898 vp_p.n24225 vp_p.n24224 0.296
R16899 vp_p.n24229 vp_p.n24228 0.296
R16900 vp_p.n24239 vp_p.n24238 0.296
R16901 vp_p.n24243 vp_p.n24242 0.296
R16902 vp_p.n24253 vp_p.n24252 0.296
R16903 vp_p.n24257 vp_p.n24256 0.296
R16904 vp_p.n24267 vp_p.n24266 0.296
R16905 vp_p.n24271 vp_p.n24270 0.296
R16906 vp_p.n24281 vp_p.n24280 0.296
R16907 vp_p.n24285 vp_p.n24284 0.296
R16908 vp_p.n24295 vp_p.n24294 0.296
R16909 vp_p.n24299 vp_p.n24298 0.296
R16910 vp_p.n24309 vp_p.n24308 0.296
R16911 vp_p.n24313 vp_p.n24312 0.296
R16912 vp_p.n24323 vp_p.n24322 0.296
R16913 vp_p.n24327 vp_p.n24326 0.296
R16914 vp_p.n24337 vp_p.n24336 0.296
R16915 vp_p.n24341 vp_p.n24340 0.296
R16916 vp_p.n24351 vp_p.n24350 0.296
R16917 vp_p.n24355 vp_p.n24354 0.296
R16918 vp_p.n24365 vp_p.n24364 0.296
R16919 vp_p.n24369 vp_p.n24368 0.296
R16920 vp_p.n24379 vp_p.n24378 0.296
R16921 vp_p.n24383 vp_p.n24382 0.296
R16922 vp_p.n24393 vp_p.n24392 0.296
R16923 vp_p.n24397 vp_p.n24396 0.296
R16924 vp_p.n24407 vp_p.n24406 0.296
R16925 vp_p.n24411 vp_p.n24410 0.296
R16926 vp_p.n24421 vp_p.n24420 0.296
R16927 vp_p.n24425 vp_p.n24424 0.296
R16928 vp_p.n24435 vp_p.n24434 0.296
R16929 vp_p.n24439 vp_p.n24438 0.296
R16930 vp_p.n24449 vp_p.n24448 0.296
R16931 vp_p.n24453 vp_p.n24452 0.296
R16932 vp_p.n24457 vp_p.n24456 0.296
R16933 vp_p.n24467 vp_p.n24466 0.296
R16934 vp_p.n24472 vp_p.n24471 0.296
R16935 vp_p.n6161 vp_p.n6160 0.296
R16936 vp_p.n6166 vp_p.n6165 0.296
R16937 vp_p.n6176 vp_p.n6175 0.296
R16938 vp_p.n6180 vp_p.n6179 0.296
R16939 vp_p.n6190 vp_p.n6189 0.296
R16940 vp_p.n6194 vp_p.n6193 0.296
R16941 vp_p.n6204 vp_p.n6203 0.296
R16942 vp_p.n6208 vp_p.n6207 0.296
R16943 vp_p.n6218 vp_p.n6217 0.296
R16944 vp_p.n6222 vp_p.n6221 0.296
R16945 vp_p.n6232 vp_p.n6231 0.296
R16946 vp_p.n6236 vp_p.n6235 0.296
R16947 vp_p.n6246 vp_p.n6245 0.296
R16948 vp_p.n6250 vp_p.n6249 0.296
R16949 vp_p.n6260 vp_p.n6259 0.296
R16950 vp_p.n6264 vp_p.n6263 0.296
R16951 vp_p.n6274 vp_p.n6273 0.296
R16952 vp_p.n6278 vp_p.n6277 0.296
R16953 vp_p.n6288 vp_p.n6287 0.296
R16954 vp_p.n6292 vp_p.n6291 0.296
R16955 vp_p.n6302 vp_p.n6301 0.296
R16956 vp_p.n6306 vp_p.n6305 0.296
R16957 vp_p.n6316 vp_p.n6315 0.296
R16958 vp_p.n6320 vp_p.n6319 0.296
R16959 vp_p.n6330 vp_p.n6329 0.296
R16960 vp_p.n6334 vp_p.n6333 0.296
R16961 vp_p.n6344 vp_p.n6343 0.296
R16962 vp_p.n6348 vp_p.n6347 0.296
R16963 vp_p.n6358 vp_p.n6357 0.296
R16964 vp_p.n6362 vp_p.n6361 0.296
R16965 vp_p.n6372 vp_p.n6371 0.296
R16966 vp_p.n6376 vp_p.n6375 0.296
R16967 vp_p.n6386 vp_p.n6385 0.296
R16968 vp_p.n6390 vp_p.n6389 0.296
R16969 vp_p.n6400 vp_p.n6399 0.296
R16970 vp_p.n6404 vp_p.n6403 0.296
R16971 vp_p.n6414 vp_p.n6413 0.296
R16972 vp_p.n6418 vp_p.n6417 0.296
R16973 vp_p.n6428 vp_p.n6427 0.296
R16974 vp_p.n6432 vp_p.n6431 0.296
R16975 vp_p.n6442 vp_p.n6441 0.296
R16976 vp_p.n6446 vp_p.n6445 0.296
R16977 vp_p.n6456 vp_p.n6455 0.296
R16978 vp_p.n6460 vp_p.n6459 0.296
R16979 vp_p.n6470 vp_p.n6469 0.296
R16980 vp_p.n6474 vp_p.n6473 0.296
R16981 vp_p.n6484 vp_p.n6483 0.296
R16982 vp_p.n6488 vp_p.n6487 0.296
R16983 vp_p.n6498 vp_p.n6497 0.296
R16984 vp_p.n6502 vp_p.n6501 0.296
R16985 vp_p.n6512 vp_p.n6511 0.296
R16986 vp_p.n6516 vp_p.n6515 0.296
R16987 vp_p.n6526 vp_p.n6525 0.296
R16988 vp_p.n6530 vp_p.n6529 0.296
R16989 vp_p.n6540 vp_p.n6539 0.296
R16990 vp_p.n6544 vp_p.n6543 0.296
R16991 vp_p.n6554 vp_p.n6553 0.296
R16992 vp_p.n6558 vp_p.n6557 0.296
R16993 vp_p.n6568 vp_p.n6567 0.296
R16994 vp_p.n6572 vp_p.n6571 0.296
R16995 vp_p.n6582 vp_p.n6581 0.296
R16996 vp_p.n6586 vp_p.n6585 0.296
R16997 vp_p.n6596 vp_p.n6595 0.296
R16998 vp_p.n6600 vp_p.n6599 0.296
R16999 vp_p.n6610 vp_p.n6609 0.296
R17000 vp_p.n6614 vp_p.n6613 0.296
R17001 vp_p.n6624 vp_p.n6623 0.296
R17002 vp_p.n6628 vp_p.n6627 0.296
R17003 vp_p.n6638 vp_p.n6637 0.296
R17004 vp_p.n6642 vp_p.n6641 0.296
R17005 vp_p.n6652 vp_p.n6651 0.296
R17006 vp_p.n6656 vp_p.n6655 0.296
R17007 vp_p.n6666 vp_p.n6665 0.296
R17008 vp_p.n6670 vp_p.n6669 0.296
R17009 vp_p.n6680 vp_p.n6679 0.296
R17010 vp_p.n6684 vp_p.n6683 0.296
R17011 vp_p.n6694 vp_p.n6693 0.296
R17012 vp_p.n6698 vp_p.n6697 0.296
R17013 vp_p.n6708 vp_p.n6707 0.296
R17014 vp_p.n6712 vp_p.n6711 0.296
R17015 vp_p.n6722 vp_p.n6721 0.296
R17016 vp_p.n6726 vp_p.n6725 0.296
R17017 vp_p.n6736 vp_p.n6735 0.296
R17018 vp_p.n6740 vp_p.n6739 0.296
R17019 vp_p.n6750 vp_p.n6749 0.296
R17020 vp_p.n6754 vp_p.n6753 0.296
R17021 vp_p.n6764 vp_p.n6763 0.296
R17022 vp_p.n6768 vp_p.n6767 0.296
R17023 vp_p.n6778 vp_p.n6777 0.296
R17024 vp_p.n6782 vp_p.n6781 0.296
R17025 vp_p.n6792 vp_p.n6791 0.296
R17026 vp_p.n6796 vp_p.n6795 0.296
R17027 vp_p.n6806 vp_p.n6805 0.296
R17028 vp_p.n6810 vp_p.n6809 0.296
R17029 vp_p.n6820 vp_p.n6819 0.296
R17030 vp_p.n6824 vp_p.n6823 0.296
R17031 vp_p.n6834 vp_p.n6833 0.296
R17032 vp_p.n6838 vp_p.n6837 0.296
R17033 vp_p.n6848 vp_p.n6847 0.296
R17034 vp_p.n6852 vp_p.n6851 0.296
R17035 vp_p.n6862 vp_p.n6861 0.296
R17036 vp_p.n6866 vp_p.n6865 0.296
R17037 vp_p.n6876 vp_p.n6875 0.296
R17038 vp_p.n6880 vp_p.n6879 0.296
R17039 vp_p.n6890 vp_p.n6889 0.296
R17040 vp_p.n6894 vp_p.n6893 0.296
R17041 vp_p.n6904 vp_p.n6903 0.296
R17042 vp_p.n6908 vp_p.n6907 0.296
R17043 vp_p.n6918 vp_p.n6917 0.296
R17044 vp_p.n6922 vp_p.n6921 0.296
R17045 vp_p.n6932 vp_p.n6931 0.296
R17046 vp_p.n6936 vp_p.n6935 0.296
R17047 vp_p.n6946 vp_p.n6945 0.296
R17048 vp_p.n6950 vp_p.n6949 0.296
R17049 vp_p.n6960 vp_p.n6959 0.296
R17050 vp_p.n6964 vp_p.n6963 0.296
R17051 vp_p.n6974 vp_p.n6973 0.296
R17052 vp_p.n6978 vp_p.n6977 0.296
R17053 vp_p.n6988 vp_p.n6987 0.296
R17054 vp_p.n6992 vp_p.n6991 0.296
R17055 vp_p.n7002 vp_p.n7001 0.296
R17056 vp_p.n7006 vp_p.n7005 0.296
R17057 vp_p.n7016 vp_p.n7015 0.296
R17058 vp_p.n7020 vp_p.n7019 0.296
R17059 vp_p.n7030 vp_p.n7029 0.296
R17060 vp_p.n7034 vp_p.n7033 0.296
R17061 vp_p.n7044 vp_p.n7043 0.296
R17062 vp_p.n7048 vp_p.n7047 0.296
R17063 vp_p.n7058 vp_p.n7057 0.296
R17064 vp_p.n7062 vp_p.n7061 0.296
R17065 vp_p.n7072 vp_p.n7071 0.296
R17066 vp_p.n7076 vp_p.n7075 0.296
R17067 vp_p.n7086 vp_p.n7085 0.296
R17068 vp_p.n7090 vp_p.n7089 0.296
R17069 vp_p.n7100 vp_p.n7099 0.296
R17070 vp_p.n7104 vp_p.n7103 0.296
R17071 vp_p.n7114 vp_p.n7113 0.296
R17072 vp_p.n7118 vp_p.n7117 0.296
R17073 vp_p.n7128 vp_p.n7127 0.296
R17074 vp_p.n7132 vp_p.n7131 0.296
R17075 vp_p.n7142 vp_p.n7141 0.296
R17076 vp_p.n7146 vp_p.n7145 0.296
R17077 vp_p.n7156 vp_p.n7155 0.296
R17078 vp_p.n7160 vp_p.n7159 0.296
R17079 vp_p.n7170 vp_p.n7169 0.296
R17080 vp_p.n7174 vp_p.n7173 0.296
R17081 vp_p.n7184 vp_p.n7183 0.296
R17082 vp_p.n7188 vp_p.n7187 0.296
R17083 vp_p.n7198 vp_p.n7197 0.296
R17084 vp_p.n24862 vp_p.n24861 0.296
R17085 vp_p.n24867 vp_p.n24866 0.296
R17086 vp_p.n24877 vp_p.n24876 0.296
R17087 vp_p.n24881 vp_p.n24880 0.296
R17088 vp_p.n24891 vp_p.n24890 0.296
R17089 vp_p.n24895 vp_p.n24894 0.296
R17090 vp_p.n24905 vp_p.n24904 0.296
R17091 vp_p.n24909 vp_p.n24908 0.296
R17092 vp_p.n24919 vp_p.n24918 0.296
R17093 vp_p.n24923 vp_p.n24922 0.296
R17094 vp_p.n24933 vp_p.n24932 0.296
R17095 vp_p.n24937 vp_p.n24936 0.296
R17096 vp_p.n24947 vp_p.n24946 0.296
R17097 vp_p.n24951 vp_p.n24950 0.296
R17098 vp_p.n24961 vp_p.n24960 0.296
R17099 vp_p.n24965 vp_p.n24964 0.296
R17100 vp_p.n24975 vp_p.n24974 0.296
R17101 vp_p.n24979 vp_p.n24978 0.296
R17102 vp_p.n24989 vp_p.n24988 0.296
R17103 vp_p.n24993 vp_p.n24992 0.296
R17104 vp_p.n25003 vp_p.n25002 0.296
R17105 vp_p.n25007 vp_p.n25006 0.296
R17106 vp_p.n25017 vp_p.n25016 0.296
R17107 vp_p.n25021 vp_p.n25020 0.296
R17108 vp_p.n25031 vp_p.n25030 0.296
R17109 vp_p.n25035 vp_p.n25034 0.296
R17110 vp_p.n25045 vp_p.n25044 0.296
R17111 vp_p.n25049 vp_p.n25048 0.296
R17112 vp_p.n25059 vp_p.n25058 0.296
R17113 vp_p.n25063 vp_p.n25062 0.296
R17114 vp_p.n25073 vp_p.n25072 0.296
R17115 vp_p.n25077 vp_p.n25076 0.296
R17116 vp_p.n25087 vp_p.n25086 0.296
R17117 vp_p.n25091 vp_p.n25090 0.296
R17118 vp_p.n25101 vp_p.n25100 0.296
R17119 vp_p.n25105 vp_p.n25104 0.296
R17120 vp_p.n25115 vp_p.n25114 0.296
R17121 vp_p.n25119 vp_p.n25118 0.296
R17122 vp_p.n25129 vp_p.n25128 0.296
R17123 vp_p.n25133 vp_p.n25132 0.296
R17124 vp_p.n25143 vp_p.n25142 0.296
R17125 vp_p.n25147 vp_p.n25146 0.296
R17126 vp_p.n25157 vp_p.n25156 0.296
R17127 vp_p.n25161 vp_p.n25160 0.296
R17128 vp_p.n25171 vp_p.n25170 0.296
R17129 vp_p.n25175 vp_p.n25174 0.296
R17130 vp_p.n25185 vp_p.n25184 0.296
R17131 vp_p.n25189 vp_p.n25188 0.296
R17132 vp_p.n25199 vp_p.n25198 0.296
R17133 vp_p.n25203 vp_p.n25202 0.296
R17134 vp_p.n25213 vp_p.n25212 0.296
R17135 vp_p.n25217 vp_p.n25216 0.296
R17136 vp_p.n25227 vp_p.n25226 0.296
R17137 vp_p.n25231 vp_p.n25230 0.296
R17138 vp_p.n25241 vp_p.n25240 0.296
R17139 vp_p.n25245 vp_p.n25244 0.296
R17140 vp_p.n25255 vp_p.n25254 0.296
R17141 vp_p.n25259 vp_p.n25258 0.296
R17142 vp_p.n25269 vp_p.n25268 0.296
R17143 vp_p.n25273 vp_p.n25272 0.296
R17144 vp_p.n25283 vp_p.n25282 0.296
R17145 vp_p.n25287 vp_p.n25286 0.296
R17146 vp_p.n25297 vp_p.n25296 0.296
R17147 vp_p.n25301 vp_p.n25300 0.296
R17148 vp_p.n25311 vp_p.n25310 0.296
R17149 vp_p.n25315 vp_p.n25314 0.296
R17150 vp_p.n25325 vp_p.n25324 0.296
R17151 vp_p.n25329 vp_p.n25328 0.296
R17152 vp_p.n25339 vp_p.n25338 0.296
R17153 vp_p.n25343 vp_p.n25342 0.296
R17154 vp_p.n25353 vp_p.n25352 0.296
R17155 vp_p.n25357 vp_p.n25356 0.296
R17156 vp_p.n25367 vp_p.n25366 0.296
R17157 vp_p.n25371 vp_p.n25370 0.296
R17158 vp_p.n25381 vp_p.n25380 0.296
R17159 vp_p.n25385 vp_p.n25384 0.296
R17160 vp_p.n25395 vp_p.n25394 0.296
R17161 vp_p.n25399 vp_p.n25398 0.296
R17162 vp_p.n25409 vp_p.n25408 0.296
R17163 vp_p.n25413 vp_p.n25412 0.296
R17164 vp_p.n25423 vp_p.n25422 0.296
R17165 vp_p.n25427 vp_p.n25426 0.296
R17166 vp_p.n25437 vp_p.n25436 0.296
R17167 vp_p.n25441 vp_p.n25440 0.296
R17168 vp_p.n25451 vp_p.n25450 0.296
R17169 vp_p.n25455 vp_p.n25454 0.296
R17170 vp_p.n25465 vp_p.n25464 0.296
R17171 vp_p.n25469 vp_p.n25468 0.296
R17172 vp_p.n25479 vp_p.n25478 0.296
R17173 vp_p.n25483 vp_p.n25482 0.296
R17174 vp_p.n25493 vp_p.n25492 0.296
R17175 vp_p.n25497 vp_p.n25496 0.296
R17176 vp_p.n25507 vp_p.n25506 0.296
R17177 vp_p.n25511 vp_p.n25510 0.296
R17178 vp_p.n25521 vp_p.n25520 0.296
R17179 vp_p.n25525 vp_p.n25524 0.296
R17180 vp_p.n25535 vp_p.n25534 0.296
R17181 vp_p.n25539 vp_p.n25538 0.296
R17182 vp_p.n25549 vp_p.n25548 0.296
R17183 vp_p.n25553 vp_p.n25552 0.296
R17184 vp_p.n25563 vp_p.n25562 0.296
R17185 vp_p.n25567 vp_p.n25566 0.296
R17186 vp_p.n25577 vp_p.n25576 0.296
R17187 vp_p.n25581 vp_p.n25580 0.296
R17188 vp_p.n25591 vp_p.n25590 0.296
R17189 vp_p.n25595 vp_p.n25594 0.296
R17190 vp_p.n25605 vp_p.n25604 0.296
R17191 vp_p.n25609 vp_p.n25608 0.296
R17192 vp_p.n25619 vp_p.n25618 0.296
R17193 vp_p.n25623 vp_p.n25622 0.296
R17194 vp_p.n25633 vp_p.n25632 0.296
R17195 vp_p.n25637 vp_p.n25636 0.296
R17196 vp_p.n25647 vp_p.n25646 0.296
R17197 vp_p.n25651 vp_p.n25650 0.296
R17198 vp_p.n25661 vp_p.n25660 0.296
R17199 vp_p.n25665 vp_p.n25664 0.296
R17200 vp_p.n25675 vp_p.n25674 0.296
R17201 vp_p.n25679 vp_p.n25678 0.296
R17202 vp_p.n25689 vp_p.n25688 0.296
R17203 vp_p.n25693 vp_p.n25692 0.296
R17204 vp_p.n25703 vp_p.n25702 0.296
R17205 vp_p.n25707 vp_p.n25706 0.296
R17206 vp_p.n25717 vp_p.n25716 0.296
R17207 vp_p.n25721 vp_p.n25720 0.296
R17208 vp_p.n25731 vp_p.n25730 0.296
R17209 vp_p.n25735 vp_p.n25734 0.296
R17210 vp_p.n25745 vp_p.n25744 0.296
R17211 vp_p.n25749 vp_p.n25748 0.296
R17212 vp_p.n25759 vp_p.n25758 0.296
R17213 vp_p.n25763 vp_p.n25762 0.296
R17214 vp_p.n25773 vp_p.n25772 0.296
R17215 vp_p.n25777 vp_p.n25776 0.296
R17216 vp_p.n25787 vp_p.n25786 0.296
R17217 vp_p.n25791 vp_p.n25790 0.296
R17218 vp_p.n25801 vp_p.n25800 0.296
R17219 vp_p.n25805 vp_p.n25804 0.296
R17220 vp_p.n25815 vp_p.n25814 0.296
R17221 vp_p.n25819 vp_p.n25818 0.296
R17222 vp_p.n25829 vp_p.n25828 0.296
R17223 vp_p.n25833 vp_p.n25832 0.296
R17224 vp_p.n25843 vp_p.n25842 0.296
R17225 vp_p.n25847 vp_p.n25846 0.296
R17226 vp_p.n25857 vp_p.n25856 0.296
R17227 vp_p.n25861 vp_p.n25860 0.296
R17228 vp_p.n25871 vp_p.n25870 0.296
R17229 vp_p.n25875 vp_p.n25874 0.296
R17230 vp_p.n25885 vp_p.n25884 0.296
R17231 vp_p.n25889 vp_p.n25888 0.296
R17232 vp_p.n25893 vp_p.n25892 0.296
R17233 vp_p.n7578 vp_p.n7577 0.296
R17234 vp_p.n7588 vp_p.n7587 0.296
R17235 vp_p.n7598 vp_p.n7597 0.296
R17236 vp_p.n7602 vp_p.n7601 0.296
R17237 vp_p.n7612 vp_p.n7611 0.296
R17238 vp_p.n7616 vp_p.n7615 0.296
R17239 vp_p.n7626 vp_p.n7625 0.296
R17240 vp_p.n7630 vp_p.n7629 0.296
R17241 vp_p.n7640 vp_p.n7639 0.296
R17242 vp_p.n7644 vp_p.n7643 0.296
R17243 vp_p.n7654 vp_p.n7653 0.296
R17244 vp_p.n7658 vp_p.n7657 0.296
R17245 vp_p.n7668 vp_p.n7667 0.296
R17246 vp_p.n7672 vp_p.n7671 0.296
R17247 vp_p.n7682 vp_p.n7681 0.296
R17248 vp_p.n7686 vp_p.n7685 0.296
R17249 vp_p.n7696 vp_p.n7695 0.296
R17250 vp_p.n7700 vp_p.n7699 0.296
R17251 vp_p.n7710 vp_p.n7709 0.296
R17252 vp_p.n7714 vp_p.n7713 0.296
R17253 vp_p.n7724 vp_p.n7723 0.296
R17254 vp_p.n7728 vp_p.n7727 0.296
R17255 vp_p.n7738 vp_p.n7737 0.296
R17256 vp_p.n7742 vp_p.n7741 0.296
R17257 vp_p.n7752 vp_p.n7751 0.296
R17258 vp_p.n7756 vp_p.n7755 0.296
R17259 vp_p.n7766 vp_p.n7765 0.296
R17260 vp_p.n7770 vp_p.n7769 0.296
R17261 vp_p.n7780 vp_p.n7779 0.296
R17262 vp_p.n7784 vp_p.n7783 0.296
R17263 vp_p.n7794 vp_p.n7793 0.296
R17264 vp_p.n7798 vp_p.n7797 0.296
R17265 vp_p.n7808 vp_p.n7807 0.296
R17266 vp_p.n7812 vp_p.n7811 0.296
R17267 vp_p.n7822 vp_p.n7821 0.296
R17268 vp_p.n7826 vp_p.n7825 0.296
R17269 vp_p.n7836 vp_p.n7835 0.296
R17270 vp_p.n7840 vp_p.n7839 0.296
R17271 vp_p.n7850 vp_p.n7849 0.296
R17272 vp_p.n7854 vp_p.n7853 0.296
R17273 vp_p.n7864 vp_p.n7863 0.296
R17274 vp_p.n7868 vp_p.n7867 0.296
R17275 vp_p.n7878 vp_p.n7877 0.296
R17276 vp_p.n7882 vp_p.n7881 0.296
R17277 vp_p.n7892 vp_p.n7891 0.296
R17278 vp_p.n7896 vp_p.n7895 0.296
R17279 vp_p.n7906 vp_p.n7905 0.296
R17280 vp_p.n7910 vp_p.n7909 0.296
R17281 vp_p.n7920 vp_p.n7919 0.296
R17282 vp_p.n7924 vp_p.n7923 0.296
R17283 vp_p.n7934 vp_p.n7933 0.296
R17284 vp_p.n7938 vp_p.n7937 0.296
R17285 vp_p.n7948 vp_p.n7947 0.296
R17286 vp_p.n7952 vp_p.n7951 0.296
R17287 vp_p.n7962 vp_p.n7961 0.296
R17288 vp_p.n7966 vp_p.n7965 0.296
R17289 vp_p.n7976 vp_p.n7975 0.296
R17290 vp_p.n7980 vp_p.n7979 0.296
R17291 vp_p.n7990 vp_p.n7989 0.296
R17292 vp_p.n7994 vp_p.n7993 0.296
R17293 vp_p.n8004 vp_p.n8003 0.296
R17294 vp_p.n8008 vp_p.n8007 0.296
R17295 vp_p.n8018 vp_p.n8017 0.296
R17296 vp_p.n8022 vp_p.n8021 0.296
R17297 vp_p.n8032 vp_p.n8031 0.296
R17298 vp_p.n8036 vp_p.n8035 0.296
R17299 vp_p.n8046 vp_p.n8045 0.296
R17300 vp_p.n8050 vp_p.n8049 0.296
R17301 vp_p.n8060 vp_p.n8059 0.296
R17302 vp_p.n8064 vp_p.n8063 0.296
R17303 vp_p.n8074 vp_p.n8073 0.296
R17304 vp_p.n8078 vp_p.n8077 0.296
R17305 vp_p.n8088 vp_p.n8087 0.296
R17306 vp_p.n8092 vp_p.n8091 0.296
R17307 vp_p.n8102 vp_p.n8101 0.296
R17308 vp_p.n8106 vp_p.n8105 0.296
R17309 vp_p.n8116 vp_p.n8115 0.296
R17310 vp_p.n8120 vp_p.n8119 0.296
R17311 vp_p.n8130 vp_p.n8129 0.296
R17312 vp_p.n8134 vp_p.n8133 0.296
R17313 vp_p.n8144 vp_p.n8143 0.296
R17314 vp_p.n8148 vp_p.n8147 0.296
R17315 vp_p.n8158 vp_p.n8157 0.296
R17316 vp_p.n8162 vp_p.n8161 0.296
R17317 vp_p.n8172 vp_p.n8171 0.296
R17318 vp_p.n8176 vp_p.n8175 0.296
R17319 vp_p.n8186 vp_p.n8185 0.296
R17320 vp_p.n8190 vp_p.n8189 0.296
R17321 vp_p.n8200 vp_p.n8199 0.296
R17322 vp_p.n8204 vp_p.n8203 0.296
R17323 vp_p.n8214 vp_p.n8213 0.296
R17324 vp_p.n8218 vp_p.n8217 0.296
R17325 vp_p.n8228 vp_p.n8227 0.296
R17326 vp_p.n8232 vp_p.n8231 0.296
R17327 vp_p.n8242 vp_p.n8241 0.296
R17328 vp_p.n8246 vp_p.n8245 0.296
R17329 vp_p.n8256 vp_p.n8255 0.296
R17330 vp_p.n8260 vp_p.n8259 0.296
R17331 vp_p.n8270 vp_p.n8269 0.296
R17332 vp_p.n8274 vp_p.n8273 0.296
R17333 vp_p.n8284 vp_p.n8283 0.296
R17334 vp_p.n8288 vp_p.n8287 0.296
R17335 vp_p.n8298 vp_p.n8297 0.296
R17336 vp_p.n8302 vp_p.n8301 0.296
R17337 vp_p.n8312 vp_p.n8311 0.296
R17338 vp_p.n8316 vp_p.n8315 0.296
R17339 vp_p.n8326 vp_p.n8325 0.296
R17340 vp_p.n8330 vp_p.n8329 0.296
R17341 vp_p.n8340 vp_p.n8339 0.296
R17342 vp_p.n8344 vp_p.n8343 0.296
R17343 vp_p.n8354 vp_p.n8353 0.296
R17344 vp_p.n8358 vp_p.n8357 0.296
R17345 vp_p.n8368 vp_p.n8367 0.296
R17346 vp_p.n8372 vp_p.n8371 0.296
R17347 vp_p.n8382 vp_p.n8381 0.296
R17348 vp_p.n8386 vp_p.n8385 0.296
R17349 vp_p.n8396 vp_p.n8395 0.296
R17350 vp_p.n8400 vp_p.n8399 0.296
R17351 vp_p.n8410 vp_p.n8409 0.296
R17352 vp_p.n8414 vp_p.n8413 0.296
R17353 vp_p.n8424 vp_p.n8423 0.296
R17354 vp_p.n8428 vp_p.n8427 0.296
R17355 vp_p.n8438 vp_p.n8437 0.296
R17356 vp_p.n8442 vp_p.n8441 0.296
R17357 vp_p.n8452 vp_p.n8451 0.296
R17358 vp_p.n8456 vp_p.n8455 0.296
R17359 vp_p.n8466 vp_p.n8465 0.296
R17360 vp_p.n8470 vp_p.n8469 0.296
R17361 vp_p.n8480 vp_p.n8479 0.296
R17362 vp_p.n8484 vp_p.n8483 0.296
R17363 vp_p.n8494 vp_p.n8493 0.296
R17364 vp_p.n8498 vp_p.n8497 0.296
R17365 vp_p.n8508 vp_p.n8507 0.296
R17366 vp_p.n8512 vp_p.n8511 0.296
R17367 vp_p.n8522 vp_p.n8521 0.296
R17368 vp_p.n8526 vp_p.n8525 0.296
R17369 vp_p.n8536 vp_p.n8535 0.296
R17370 vp_p.n8540 vp_p.n8539 0.296
R17371 vp_p.n8550 vp_p.n8549 0.296
R17372 vp_p.n8554 vp_p.n8553 0.296
R17373 vp_p.n8564 vp_p.n8563 0.296
R17374 vp_p.n8568 vp_p.n8567 0.296
R17375 vp_p.n8578 vp_p.n8577 0.296
R17376 vp_p.n8582 vp_p.n8581 0.296
R17377 vp_p.n8592 vp_p.n8591 0.296
R17378 vp_p.n8596 vp_p.n8595 0.296
R17379 vp_p.n8606 vp_p.n8605 0.296
R17380 vp_p.n8610 vp_p.n8609 0.296
R17381 vp_p.n8620 vp_p.n8619 0.296
R17382 vp_p.n26288 vp_p.n26287 0.296
R17383 vp_p.n26292 vp_p.n26291 0.296
R17384 vp_p.n26302 vp_p.n26301 0.296
R17385 vp_p.n26306 vp_p.n26305 0.296
R17386 vp_p.n26316 vp_p.n26315 0.296
R17387 vp_p.n26320 vp_p.n26319 0.296
R17388 vp_p.n26330 vp_p.n26329 0.296
R17389 vp_p.n26334 vp_p.n26333 0.296
R17390 vp_p.n26344 vp_p.n26343 0.296
R17391 vp_p.n26348 vp_p.n26347 0.296
R17392 vp_p.n26358 vp_p.n26357 0.296
R17393 vp_p.n26362 vp_p.n26361 0.296
R17394 vp_p.n26372 vp_p.n26371 0.296
R17395 vp_p.n26376 vp_p.n26375 0.296
R17396 vp_p.n26386 vp_p.n26385 0.296
R17397 vp_p.n26390 vp_p.n26389 0.296
R17398 vp_p.n26400 vp_p.n26399 0.296
R17399 vp_p.n26404 vp_p.n26403 0.296
R17400 vp_p.n26414 vp_p.n26413 0.296
R17401 vp_p.n26418 vp_p.n26417 0.296
R17402 vp_p.n26428 vp_p.n26427 0.296
R17403 vp_p.n26432 vp_p.n26431 0.296
R17404 vp_p.n26442 vp_p.n26441 0.296
R17405 vp_p.n26446 vp_p.n26445 0.296
R17406 vp_p.n26456 vp_p.n26455 0.296
R17407 vp_p.n26460 vp_p.n26459 0.296
R17408 vp_p.n26470 vp_p.n26469 0.296
R17409 vp_p.n26474 vp_p.n26473 0.296
R17410 vp_p.n26484 vp_p.n26483 0.296
R17411 vp_p.n26488 vp_p.n26487 0.296
R17412 vp_p.n26498 vp_p.n26497 0.296
R17413 vp_p.n26502 vp_p.n26501 0.296
R17414 vp_p.n26512 vp_p.n26511 0.296
R17415 vp_p.n26516 vp_p.n26515 0.296
R17416 vp_p.n26526 vp_p.n26525 0.296
R17417 vp_p.n26530 vp_p.n26529 0.296
R17418 vp_p.n26540 vp_p.n26539 0.296
R17419 vp_p.n26544 vp_p.n26543 0.296
R17420 vp_p.n26554 vp_p.n26553 0.296
R17421 vp_p.n26558 vp_p.n26557 0.296
R17422 vp_p.n26568 vp_p.n26567 0.296
R17423 vp_p.n26572 vp_p.n26571 0.296
R17424 vp_p.n26582 vp_p.n26581 0.296
R17425 vp_p.n26586 vp_p.n26585 0.296
R17426 vp_p.n26596 vp_p.n26595 0.296
R17427 vp_p.n26600 vp_p.n26599 0.296
R17428 vp_p.n26610 vp_p.n26609 0.296
R17429 vp_p.n26614 vp_p.n26613 0.296
R17430 vp_p.n26624 vp_p.n26623 0.296
R17431 vp_p.n26628 vp_p.n26627 0.296
R17432 vp_p.n26638 vp_p.n26637 0.296
R17433 vp_p.n26642 vp_p.n26641 0.296
R17434 vp_p.n26652 vp_p.n26651 0.296
R17435 vp_p.n26656 vp_p.n26655 0.296
R17436 vp_p.n26666 vp_p.n26665 0.296
R17437 vp_p.n26670 vp_p.n26669 0.296
R17438 vp_p.n26680 vp_p.n26679 0.296
R17439 vp_p.n26684 vp_p.n26683 0.296
R17440 vp_p.n26694 vp_p.n26693 0.296
R17441 vp_p.n26698 vp_p.n26697 0.296
R17442 vp_p.n26708 vp_p.n26707 0.296
R17443 vp_p.n26712 vp_p.n26711 0.296
R17444 vp_p.n26722 vp_p.n26721 0.296
R17445 vp_p.n26726 vp_p.n26725 0.296
R17446 vp_p.n26736 vp_p.n26735 0.296
R17447 vp_p.n26740 vp_p.n26739 0.296
R17448 vp_p.n26750 vp_p.n26749 0.296
R17449 vp_p.n26754 vp_p.n26753 0.296
R17450 vp_p.n26764 vp_p.n26763 0.296
R17451 vp_p.n26768 vp_p.n26767 0.296
R17452 vp_p.n26778 vp_p.n26777 0.296
R17453 vp_p.n26782 vp_p.n26781 0.296
R17454 vp_p.n26792 vp_p.n26791 0.296
R17455 vp_p.n26796 vp_p.n26795 0.296
R17456 vp_p.n26806 vp_p.n26805 0.296
R17457 vp_p.n26810 vp_p.n26809 0.296
R17458 vp_p.n26820 vp_p.n26819 0.296
R17459 vp_p.n26824 vp_p.n26823 0.296
R17460 vp_p.n26834 vp_p.n26833 0.296
R17461 vp_p.n26838 vp_p.n26837 0.296
R17462 vp_p.n26848 vp_p.n26847 0.296
R17463 vp_p.n26852 vp_p.n26851 0.296
R17464 vp_p.n26862 vp_p.n26861 0.296
R17465 vp_p.n26866 vp_p.n26865 0.296
R17466 vp_p.n26876 vp_p.n26875 0.296
R17467 vp_p.n26880 vp_p.n26879 0.296
R17468 vp_p.n26890 vp_p.n26889 0.296
R17469 vp_p.n26894 vp_p.n26893 0.296
R17470 vp_p.n26904 vp_p.n26903 0.296
R17471 vp_p.n26908 vp_p.n26907 0.296
R17472 vp_p.n26918 vp_p.n26917 0.296
R17473 vp_p.n26922 vp_p.n26921 0.296
R17474 vp_p.n26932 vp_p.n26931 0.296
R17475 vp_p.n26936 vp_p.n26935 0.296
R17476 vp_p.n26946 vp_p.n26945 0.296
R17477 vp_p.n26950 vp_p.n26949 0.296
R17478 vp_p.n26960 vp_p.n26959 0.296
R17479 vp_p.n26964 vp_p.n26963 0.296
R17480 vp_p.n26974 vp_p.n26973 0.296
R17481 vp_p.n26978 vp_p.n26977 0.296
R17482 vp_p.n26988 vp_p.n26987 0.296
R17483 vp_p.n26992 vp_p.n26991 0.296
R17484 vp_p.n27002 vp_p.n27001 0.296
R17485 vp_p.n27006 vp_p.n27005 0.296
R17486 vp_p.n27016 vp_p.n27015 0.296
R17487 vp_p.n27020 vp_p.n27019 0.296
R17488 vp_p.n27030 vp_p.n27029 0.296
R17489 vp_p.n27034 vp_p.n27033 0.296
R17490 vp_p.n27044 vp_p.n27043 0.296
R17491 vp_p.n27048 vp_p.n27047 0.296
R17492 vp_p.n27058 vp_p.n27057 0.296
R17493 vp_p.n27062 vp_p.n27061 0.296
R17494 vp_p.n27072 vp_p.n27071 0.296
R17495 vp_p.n27076 vp_p.n27075 0.296
R17496 vp_p.n27086 vp_p.n27085 0.296
R17497 vp_p.n27090 vp_p.n27089 0.296
R17498 vp_p.n27100 vp_p.n27099 0.296
R17499 vp_p.n27104 vp_p.n27103 0.296
R17500 vp_p.n27114 vp_p.n27113 0.296
R17501 vp_p.n27118 vp_p.n27117 0.296
R17502 vp_p.n27128 vp_p.n27127 0.296
R17503 vp_p.n27132 vp_p.n27131 0.296
R17504 vp_p.n27142 vp_p.n27141 0.296
R17505 vp_p.n27146 vp_p.n27145 0.296
R17506 vp_p.n27156 vp_p.n27155 0.296
R17507 vp_p.n27160 vp_p.n27159 0.296
R17508 vp_p.n27170 vp_p.n27169 0.296
R17509 vp_p.n27174 vp_p.n27173 0.296
R17510 vp_p.n27184 vp_p.n27183 0.296
R17511 vp_p.n27188 vp_p.n27187 0.296
R17512 vp_p.n27198 vp_p.n27197 0.296
R17513 vp_p.n27202 vp_p.n27201 0.296
R17514 vp_p.n27212 vp_p.n27211 0.296
R17515 vp_p.n27216 vp_p.n27215 0.296
R17516 vp_p.n27226 vp_p.n27225 0.296
R17517 vp_p.n27230 vp_p.n27229 0.296
R17518 vp_p.n27240 vp_p.n27239 0.296
R17519 vp_p.n27244 vp_p.n27243 0.296
R17520 vp_p.n27254 vp_p.n27253 0.296
R17521 vp_p.n27258 vp_p.n27257 0.296
R17522 vp_p.n27268 vp_p.n27267 0.296
R17523 vp_p.n27272 vp_p.n27271 0.296
R17524 vp_p.n27282 vp_p.n27281 0.296
R17525 vp_p.n27286 vp_p.n27285 0.296
R17526 vp_p.n27296 vp_p.n27295 0.296
R17527 vp_p.n27300 vp_p.n27299 0.296
R17528 vp_p.n27310 vp_p.n27309 0.296
R17529 vp_p.n27314 vp_p.n27313 0.296
R17530 vp_p.n27324 vp_p.n27323 0.296
R17531 vp_p.n9204 vp_p.n9203 0.289
R17532 vp_p.n458 vp_p.n457 0.289
R17533 vp_p.n27435 vp_p.n14466 0.227
R17534 vp_p.n27436 vp_p.n13097 0.227
R17535 vp_p.n27434 vp_p.n15899 0.227
R17536 vp_p.n27437 vp_p.n11663 0.227
R17537 vp_p.n27433 vp_p.n17331 0.227
R17538 vp_p.n27438 vp_p.n10230 0.227
R17539 vp_p.n27432 vp_p.n18762 0.227
R17540 vp_p.n8733 vp_p.n1488 0.227
R17541 vp_p.n27431 vp_p.n20192 0.227
R17542 vp_p.n8732 vp_p.n2918 0.227
R17543 vp_p.n27430 vp_p.n21621 0.227
R17544 vp_p.n8731 vp_p.n4347 0.227
R17545 vp_p.n27429 vp_p.n23049 0.227
R17546 vp_p.n8730 vp_p.n5775 0.227
R17547 vp_p.n27428 vp_p.n24476 0.227
R17548 vp_p.n8729 vp_p.n7202 0.227
R17549 vp_p.n27427 vp_p.n25902 0.227
R17550 vp_p.n8728 vp_p.n8629 0.227
R17551 vp_p.n27426 vp_p.n27327 0.227
R17552 vp_p.n8729 vp_p.n8728 0.212
R17553 vp_p.n8730 vp_p.n8729 0.212
R17554 vp_p.n8731 vp_p.n8730 0.212
R17555 vp_p.n8732 vp_p.n8731 0.212
R17556 vp_p.n8733 vp_p.n8732 0.212
R17557 vp_p.n27438 vp_p.n27437 0.212
R17558 vp_p.n27437 vp_p.n27436 0.212
R17559 vp_p.n27436 vp_p.n27435 0.212
R17560 vp_p.n27435 vp_p.n27434 0.212
R17561 vp_p.n27434 vp_p.n27433 0.212
R17562 vp_p.n27433 vp_p.n27432 0.212
R17563 vp_p.n27432 vp_p.n27431 0.212
R17564 vp_p.n27431 vp_p.n27430 0.212
R17565 vp_p.n27430 vp_p.n27429 0.212
R17566 vp_p.n27429 vp_p.n27428 0.212
R17567 vp_p.n27428 vp_p.n27427 0.212
R17568 vp_p.n27427 vp_p.n27426 0.212
R17569 vp_p.n453 vp_p.n452 0.201
R17570 vp_p.n454 vp_p.n453 0.201
R17571 vp_p.n455 vp_p.n454 0.201
R17572 vp_p.n456 vp_p.n455 0.201
R17573 vp_p.n457 vp_p.n456 0.201
R17574 vp_p.n9203 vp_p.n9202 0.201
R17575 vp_p.n9202 vp_p.n9201 0.201
R17576 vp_p.n9201 vp_p.n9200 0.201
R17577 vp_p.n9200 vp_p.n9199 0.201
R17578 vp_p.n9199 vp_p.n9198 0.201
R17579 vp_p.n9198 vp_p.n9197 0.201
R17580 vp_p.n9197 vp_p.n9196 0.201
R17581 vp_p.n9196 vp_p.n9195 0.201
R17582 vp_p.n9195 vp_p.n9194 0.201
R17583 vp_p.n9194 vp_p.n9193 0.201
R17584 vp_p.n9193 vp_p.n9192 0.201
R17585 vp_p.n9192 vp_p.n9191 0.201
R17586 vp_p vp_p.n27438 0.149
R17587 vp_p vp_p.n8733 0.063
R17588 vp_p.n13856 vp_p.n13855 0.013
R17589 vp_p.n13860 vp_p.n13859 0.013
R17590 vp_p.n13864 vp_p.n13863 0.013
R17591 vp_p.n13868 vp_p.n13867 0.013
R17592 vp_p.n13872 vp_p.n13871 0.013
R17593 vp_p.n13876 vp_p.n13875 0.013
R17594 vp_p.n13880 vp_p.n13879 0.013
R17595 vp_p.n13884 vp_p.n13883 0.013
R17596 vp_p.n13888 vp_p.n13887 0.013
R17597 vp_p.n13892 vp_p.n13891 0.013
R17598 vp_p.n13896 vp_p.n13895 0.013
R17599 vp_p.n13900 vp_p.n13899 0.013
R17600 vp_p.n13904 vp_p.n13903 0.013
R17601 vp_p.n13908 vp_p.n13907 0.013
R17602 vp_p.n13912 vp_p.n13911 0.013
R17603 vp_p.n13916 vp_p.n13915 0.013
R17604 vp_p.n13920 vp_p.n13919 0.013
R17605 vp_p.n13924 vp_p.n13923 0.013
R17606 vp_p.n13928 vp_p.n13927 0.013
R17607 vp_p.n13932 vp_p.n13931 0.013
R17608 vp_p.n13936 vp_p.n13935 0.013
R17609 vp_p.n13940 vp_p.n13939 0.013
R17610 vp_p.n13944 vp_p.n13943 0.013
R17611 vp_p.n13948 vp_p.n13947 0.013
R17612 vp_p.n13952 vp_p.n13951 0.013
R17613 vp_p.n13956 vp_p.n13955 0.013
R17614 vp_p.n13960 vp_p.n13959 0.013
R17615 vp_p.n13964 vp_p.n13963 0.013
R17616 vp_p.n13968 vp_p.n13967 0.013
R17617 vp_p.n13972 vp_p.n13971 0.013
R17618 vp_p.n13976 vp_p.n13975 0.013
R17619 vp_p.n13980 vp_p.n13979 0.013
R17620 vp_p.n13984 vp_p.n13983 0.013
R17621 vp_p.n13988 vp_p.n13987 0.013
R17622 vp_p.n13992 vp_p.n13991 0.013
R17623 vp_p.n13996 vp_p.n13995 0.013
R17624 vp_p.n14000 vp_p.n13999 0.013
R17625 vp_p.n14004 vp_p.n14003 0.013
R17626 vp_p.n14008 vp_p.n14007 0.013
R17627 vp_p.n14012 vp_p.n14011 0.013
R17628 vp_p.n14016 vp_p.n14015 0.013
R17629 vp_p.n14020 vp_p.n14019 0.013
R17630 vp_p.n14024 vp_p.n14023 0.013
R17631 vp_p.n14028 vp_p.n14027 0.013
R17632 vp_p.n14032 vp_p.n14031 0.013
R17633 vp_p.n14036 vp_p.n14035 0.013
R17634 vp_p.n14040 vp_p.n14039 0.013
R17635 vp_p.n14044 vp_p.n14043 0.013
R17636 vp_p.n14048 vp_p.n14047 0.013
R17637 vp_p.n14052 vp_p.n14051 0.013
R17638 vp_p.n14056 vp_p.n14055 0.013
R17639 vp_p.n14060 vp_p.n14059 0.013
R17640 vp_p.n14064 vp_p.n14063 0.013
R17641 vp_p.n14068 vp_p.n14067 0.013
R17642 vp_p.n14072 vp_p.n14071 0.013
R17643 vp_p.n14076 vp_p.n14075 0.013
R17644 vp_p.n14080 vp_p.n14079 0.013
R17645 vp_p.n14084 vp_p.n14083 0.013
R17646 vp_p.n14088 vp_p.n14087 0.013
R17647 vp_p.n14092 vp_p.n14091 0.013
R17648 vp_p.n14096 vp_p.n14095 0.013
R17649 vp_p.n14100 vp_p.n14099 0.013
R17650 vp_p.n14104 vp_p.n14103 0.013
R17651 vp_p.n14108 vp_p.n14107 0.013
R17652 vp_p.n14112 vp_p.n14111 0.013
R17653 vp_p.n14116 vp_p.n14115 0.013
R17654 vp_p.n14120 vp_p.n14119 0.013
R17655 vp_p.n14124 vp_p.n14123 0.013
R17656 vp_p.n14128 vp_p.n14127 0.013
R17657 vp_p.n14132 vp_p.n14131 0.013
R17658 vp_p.n14136 vp_p.n14135 0.013
R17659 vp_p.n14140 vp_p.n14139 0.013
R17660 vp_p.n14144 vp_p.n14143 0.013
R17661 vp_p.n14148 vp_p.n14147 0.013
R17662 vp_p.n14152 vp_p.n14151 0.013
R17663 vp_p.n14156 vp_p.n14155 0.013
R17664 vp_p.n14160 vp_p.n14159 0.013
R17665 vp_p.n14164 vp_p.n14163 0.013
R17666 vp_p.n14168 vp_p.n14167 0.013
R17667 vp_p.n14172 vp_p.n14171 0.013
R17668 vp_p.n14176 vp_p.n14175 0.013
R17669 vp_p.n14180 vp_p.n14179 0.013
R17670 vp_p.n14184 vp_p.n14183 0.013
R17671 vp_p.n14188 vp_p.n14187 0.013
R17672 vp_p.n14192 vp_p.n14191 0.013
R17673 vp_p.n14196 vp_p.n14195 0.013
R17674 vp_p.n14200 vp_p.n14199 0.013
R17675 vp_p.n14204 vp_p.n14203 0.013
R17676 vp_p.n14208 vp_p.n14207 0.013
R17677 vp_p.n14212 vp_p.n14211 0.013
R17678 vp_p.n14216 vp_p.n14215 0.013
R17679 vp_p.n14220 vp_p.n14219 0.013
R17680 vp_p.n14224 vp_p.n14223 0.013
R17681 vp_p.n14228 vp_p.n14227 0.013
R17682 vp_p.n14232 vp_p.n14231 0.013
R17683 vp_p.n14236 vp_p.n14235 0.013
R17684 vp_p.n14240 vp_p.n14239 0.013
R17685 vp_p.n14244 vp_p.n14243 0.013
R17686 vp_p.n14248 vp_p.n14247 0.013
R17687 vp_p.n14252 vp_p.n14251 0.013
R17688 vp_p.n14256 vp_p.n14255 0.013
R17689 vp_p.n14260 vp_p.n14259 0.013
R17690 vp_p.n14264 vp_p.n14263 0.013
R17691 vp_p.n14268 vp_p.n14267 0.013
R17692 vp_p.n14272 vp_p.n14271 0.013
R17693 vp_p.n14276 vp_p.n14275 0.013
R17694 vp_p.n14280 vp_p.n14279 0.013
R17695 vp_p.n14284 vp_p.n14283 0.013
R17696 vp_p.n14288 vp_p.n14287 0.013
R17697 vp_p.n14292 vp_p.n14291 0.013
R17698 vp_p.n14296 vp_p.n14295 0.013
R17699 vp_p.n14300 vp_p.n14299 0.013
R17700 vp_p.n14304 vp_p.n14303 0.013
R17701 vp_p.n14308 vp_p.n14307 0.013
R17702 vp_p.n14312 vp_p.n14311 0.013
R17703 vp_p.n14316 vp_p.n14315 0.013
R17704 vp_p.n14320 vp_p.n14319 0.013
R17705 vp_p.n14324 vp_p.n14323 0.013
R17706 vp_p.n14328 vp_p.n14327 0.013
R17707 vp_p.n14332 vp_p.n14331 0.013
R17708 vp_p.n14336 vp_p.n14335 0.013
R17709 vp_p.n14340 vp_p.n14339 0.013
R17710 vp_p.n14344 vp_p.n14343 0.013
R17711 vp_p.n14348 vp_p.n14347 0.013
R17712 vp_p.n14352 vp_p.n14351 0.013
R17713 vp_p.n14356 vp_p.n14355 0.013
R17714 vp_p.n14360 vp_p.n14359 0.013
R17715 vp_p.n14364 vp_p.n14363 0.013
R17716 vp_p.n14368 vp_p.n14367 0.013
R17717 vp_p.n14372 vp_p.n14371 0.013
R17718 vp_p.n14376 vp_p.n14375 0.013
R17719 vp_p.n12102 vp_p.n12101 0.013
R17720 vp_p.n12116 vp_p.n12115 0.013
R17721 vp_p.n12130 vp_p.n12129 0.013
R17722 vp_p.n12144 vp_p.n12143 0.013
R17723 vp_p.n12158 vp_p.n12157 0.013
R17724 vp_p.n12172 vp_p.n12171 0.013
R17725 vp_p.n12186 vp_p.n12185 0.013
R17726 vp_p.n12200 vp_p.n12199 0.013
R17727 vp_p.n12214 vp_p.n12213 0.013
R17728 vp_p.n12228 vp_p.n12227 0.013
R17729 vp_p.n12242 vp_p.n12241 0.013
R17730 vp_p.n12256 vp_p.n12255 0.013
R17731 vp_p.n12270 vp_p.n12269 0.013
R17732 vp_p.n12284 vp_p.n12283 0.013
R17733 vp_p.n12298 vp_p.n12297 0.013
R17734 vp_p.n12312 vp_p.n12311 0.013
R17735 vp_p.n12326 vp_p.n12325 0.013
R17736 vp_p.n12340 vp_p.n12339 0.013
R17737 vp_p.n12354 vp_p.n12353 0.013
R17738 vp_p.n12368 vp_p.n12367 0.013
R17739 vp_p.n12382 vp_p.n12381 0.013
R17740 vp_p.n12396 vp_p.n12395 0.013
R17741 vp_p.n12410 vp_p.n12409 0.013
R17742 vp_p.n12424 vp_p.n12423 0.013
R17743 vp_p.n12438 vp_p.n12437 0.013
R17744 vp_p.n12452 vp_p.n12451 0.013
R17745 vp_p.n12466 vp_p.n12465 0.013
R17746 vp_p.n12480 vp_p.n12479 0.013
R17747 vp_p.n12494 vp_p.n12493 0.013
R17748 vp_p.n12508 vp_p.n12507 0.013
R17749 vp_p.n12522 vp_p.n12521 0.013
R17750 vp_p.n12536 vp_p.n12535 0.013
R17751 vp_p.n12550 vp_p.n12549 0.013
R17752 vp_p.n12564 vp_p.n12563 0.013
R17753 vp_p.n12578 vp_p.n12577 0.013
R17754 vp_p.n12592 vp_p.n12591 0.013
R17755 vp_p.n12606 vp_p.n12605 0.013
R17756 vp_p.n12620 vp_p.n12619 0.013
R17757 vp_p.n12634 vp_p.n12633 0.013
R17758 vp_p.n12648 vp_p.n12647 0.013
R17759 vp_p.n12662 vp_p.n12661 0.013
R17760 vp_p.n12676 vp_p.n12675 0.013
R17761 vp_p.n12690 vp_p.n12689 0.013
R17762 vp_p.n12704 vp_p.n12703 0.013
R17763 vp_p.n12718 vp_p.n12717 0.013
R17764 vp_p.n12732 vp_p.n12731 0.013
R17765 vp_p.n12746 vp_p.n12745 0.013
R17766 vp_p.n12760 vp_p.n12759 0.013
R17767 vp_p.n12774 vp_p.n12773 0.013
R17768 vp_p.n12788 vp_p.n12787 0.013
R17769 vp_p.n12802 vp_p.n12801 0.013
R17770 vp_p.n12816 vp_p.n12815 0.013
R17771 vp_p.n12830 vp_p.n12829 0.013
R17772 vp_p.n12844 vp_p.n12843 0.013
R17773 vp_p.n12858 vp_p.n12857 0.013
R17774 vp_p.n12872 vp_p.n12871 0.013
R17775 vp_p.n12886 vp_p.n12885 0.013
R17776 vp_p.n12900 vp_p.n12899 0.013
R17777 vp_p.n12914 vp_p.n12913 0.013
R17778 vp_p.n12928 vp_p.n12927 0.013
R17779 vp_p.n12942 vp_p.n12941 0.013
R17780 vp_p.n12956 vp_p.n12955 0.013
R17781 vp_p.n12970 vp_p.n12969 0.013
R17782 vp_p.n12984 vp_p.n12983 0.013
R17783 vp_p.n12998 vp_p.n12997 0.013
R17784 vp_p.n13012 vp_p.n13011 0.013
R17785 vp_p.n14905 vp_p.n14904 0.013
R17786 vp_p.n14919 vp_p.n14918 0.013
R17787 vp_p.n14933 vp_p.n14932 0.013
R17788 vp_p.n14947 vp_p.n14946 0.013
R17789 vp_p.n14961 vp_p.n14960 0.013
R17790 vp_p.n14975 vp_p.n14974 0.013
R17791 vp_p.n14989 vp_p.n14988 0.013
R17792 vp_p.n15003 vp_p.n15002 0.013
R17793 vp_p.n15017 vp_p.n15016 0.013
R17794 vp_p.n15031 vp_p.n15030 0.013
R17795 vp_p.n15045 vp_p.n15044 0.013
R17796 vp_p.n15059 vp_p.n15058 0.013
R17797 vp_p.n15073 vp_p.n15072 0.013
R17798 vp_p.n15087 vp_p.n15086 0.013
R17799 vp_p.n15101 vp_p.n15100 0.013
R17800 vp_p.n15115 vp_p.n15114 0.013
R17801 vp_p.n15129 vp_p.n15128 0.013
R17802 vp_p.n15143 vp_p.n15142 0.013
R17803 vp_p.n15157 vp_p.n15156 0.013
R17804 vp_p.n15171 vp_p.n15170 0.013
R17805 vp_p.n15185 vp_p.n15184 0.013
R17806 vp_p.n15199 vp_p.n15198 0.013
R17807 vp_p.n15213 vp_p.n15212 0.013
R17808 vp_p.n15227 vp_p.n15226 0.013
R17809 vp_p.n15241 vp_p.n15240 0.013
R17810 vp_p.n15255 vp_p.n15254 0.013
R17811 vp_p.n15269 vp_p.n15268 0.013
R17812 vp_p.n15283 vp_p.n15282 0.013
R17813 vp_p.n15297 vp_p.n15296 0.013
R17814 vp_p.n15311 vp_p.n15310 0.013
R17815 vp_p.n15325 vp_p.n15324 0.013
R17816 vp_p.n15339 vp_p.n15338 0.013
R17817 vp_p.n15353 vp_p.n15352 0.013
R17818 vp_p.n15367 vp_p.n15366 0.013
R17819 vp_p.n15381 vp_p.n15380 0.013
R17820 vp_p.n15395 vp_p.n15394 0.013
R17821 vp_p.n15409 vp_p.n15408 0.013
R17822 vp_p.n15423 vp_p.n15422 0.013
R17823 vp_p.n15437 vp_p.n15436 0.013
R17824 vp_p.n15451 vp_p.n15450 0.013
R17825 vp_p.n15465 vp_p.n15464 0.013
R17826 vp_p.n15479 vp_p.n15478 0.013
R17827 vp_p.n15493 vp_p.n15492 0.013
R17828 vp_p.n15507 vp_p.n15506 0.013
R17829 vp_p.n15521 vp_p.n15520 0.013
R17830 vp_p.n15535 vp_p.n15534 0.013
R17831 vp_p.n15549 vp_p.n15548 0.013
R17832 vp_p.n15563 vp_p.n15562 0.013
R17833 vp_p.n15577 vp_p.n15576 0.013
R17834 vp_p.n15591 vp_p.n15590 0.013
R17835 vp_p.n15605 vp_p.n15604 0.013
R17836 vp_p.n15619 vp_p.n15618 0.013
R17837 vp_p.n15633 vp_p.n15632 0.013
R17838 vp_p.n15647 vp_p.n15646 0.013
R17839 vp_p.n15661 vp_p.n15660 0.013
R17840 vp_p.n15675 vp_p.n15674 0.013
R17841 vp_p.n15689 vp_p.n15688 0.013
R17842 vp_p.n15703 vp_p.n15702 0.013
R17843 vp_p.n15717 vp_p.n15716 0.013
R17844 vp_p.n15731 vp_p.n15730 0.013
R17845 vp_p.n15745 vp_p.n15744 0.013
R17846 vp_p.n15759 vp_p.n15758 0.013
R17847 vp_p.n15773 vp_p.n15772 0.013
R17848 vp_p.n15787 vp_p.n15786 0.013
R17849 vp_p.n15801 vp_p.n15800 0.013
R17850 vp_p.n15815 vp_p.n15814 0.013
R17851 vp_p.n15819 vp_p.n15818 0.013
R17852 vp_p.n10664 vp_p.n10663 0.013
R17853 vp_p.n10678 vp_p.n10677 0.013
R17854 vp_p.n10692 vp_p.n10691 0.013
R17855 vp_p.n10706 vp_p.n10705 0.013
R17856 vp_p.n10720 vp_p.n10719 0.013
R17857 vp_p.n10734 vp_p.n10733 0.013
R17858 vp_p.n10748 vp_p.n10747 0.013
R17859 vp_p.n10762 vp_p.n10761 0.013
R17860 vp_p.n10776 vp_p.n10775 0.013
R17861 vp_p.n10790 vp_p.n10789 0.013
R17862 vp_p.n10804 vp_p.n10803 0.013
R17863 vp_p.n10818 vp_p.n10817 0.013
R17864 vp_p.n10832 vp_p.n10831 0.013
R17865 vp_p.n10846 vp_p.n10845 0.013
R17866 vp_p.n10860 vp_p.n10859 0.013
R17867 vp_p.n10874 vp_p.n10873 0.013
R17868 vp_p.n10888 vp_p.n10887 0.013
R17869 vp_p.n10902 vp_p.n10901 0.013
R17870 vp_p.n10916 vp_p.n10915 0.013
R17871 vp_p.n10930 vp_p.n10929 0.013
R17872 vp_p.n10944 vp_p.n10943 0.013
R17873 vp_p.n10958 vp_p.n10957 0.013
R17874 vp_p.n10972 vp_p.n10971 0.013
R17875 vp_p.n10986 vp_p.n10985 0.013
R17876 vp_p.n11000 vp_p.n10999 0.013
R17877 vp_p.n11014 vp_p.n11013 0.013
R17878 vp_p.n11028 vp_p.n11027 0.013
R17879 vp_p.n11042 vp_p.n11041 0.013
R17880 vp_p.n11056 vp_p.n11055 0.013
R17881 vp_p.n11070 vp_p.n11069 0.013
R17882 vp_p.n11084 vp_p.n11083 0.013
R17883 vp_p.n11098 vp_p.n11097 0.013
R17884 vp_p.n11112 vp_p.n11111 0.013
R17885 vp_p.n11126 vp_p.n11125 0.013
R17886 vp_p.n11140 vp_p.n11139 0.013
R17887 vp_p.n11154 vp_p.n11153 0.013
R17888 vp_p.n11168 vp_p.n11167 0.013
R17889 vp_p.n11182 vp_p.n11181 0.013
R17890 vp_p.n11196 vp_p.n11195 0.013
R17891 vp_p.n11210 vp_p.n11209 0.013
R17892 vp_p.n11224 vp_p.n11223 0.013
R17893 vp_p.n11238 vp_p.n11237 0.013
R17894 vp_p.n11252 vp_p.n11251 0.013
R17895 vp_p.n11266 vp_p.n11265 0.013
R17896 vp_p.n11280 vp_p.n11279 0.013
R17897 vp_p.n11294 vp_p.n11293 0.013
R17898 vp_p.n11308 vp_p.n11307 0.013
R17899 vp_p.n11322 vp_p.n11321 0.013
R17900 vp_p.n11336 vp_p.n11335 0.013
R17901 vp_p.n11350 vp_p.n11349 0.013
R17902 vp_p.n11364 vp_p.n11363 0.013
R17903 vp_p.n11378 vp_p.n11377 0.013
R17904 vp_p.n11392 vp_p.n11391 0.013
R17905 vp_p.n11406 vp_p.n11405 0.013
R17906 vp_p.n11420 vp_p.n11419 0.013
R17907 vp_p.n11434 vp_p.n11433 0.013
R17908 vp_p.n11448 vp_p.n11447 0.013
R17909 vp_p.n11462 vp_p.n11461 0.013
R17910 vp_p.n11476 vp_p.n11475 0.013
R17911 vp_p.n11490 vp_p.n11489 0.013
R17912 vp_p.n11504 vp_p.n11503 0.013
R17913 vp_p.n11518 vp_p.n11517 0.013
R17914 vp_p.n11532 vp_p.n11531 0.013
R17915 vp_p.n11546 vp_p.n11545 0.013
R17916 vp_p.n11560 vp_p.n11559 0.013
R17917 vp_p.n11574 vp_p.n11573 0.013
R17918 vp_p.n11588 vp_p.n11587 0.013
R17919 vp_p.n16333 vp_p.n16332 0.013
R17920 vp_p.n16347 vp_p.n16346 0.013
R17921 vp_p.n16361 vp_p.n16360 0.013
R17922 vp_p.n16375 vp_p.n16374 0.013
R17923 vp_p.n16389 vp_p.n16388 0.013
R17924 vp_p.n16403 vp_p.n16402 0.013
R17925 vp_p.n16417 vp_p.n16416 0.013
R17926 vp_p.n16431 vp_p.n16430 0.013
R17927 vp_p.n16445 vp_p.n16444 0.013
R17928 vp_p.n16459 vp_p.n16458 0.013
R17929 vp_p.n16473 vp_p.n16472 0.013
R17930 vp_p.n16487 vp_p.n16486 0.013
R17931 vp_p.n16501 vp_p.n16500 0.013
R17932 vp_p.n16515 vp_p.n16514 0.013
R17933 vp_p.n16529 vp_p.n16528 0.013
R17934 vp_p.n16543 vp_p.n16542 0.013
R17935 vp_p.n16557 vp_p.n16556 0.013
R17936 vp_p.n16571 vp_p.n16570 0.013
R17937 vp_p.n16585 vp_p.n16584 0.013
R17938 vp_p.n16599 vp_p.n16598 0.013
R17939 vp_p.n16613 vp_p.n16612 0.013
R17940 vp_p.n16627 vp_p.n16626 0.013
R17941 vp_p.n16641 vp_p.n16640 0.013
R17942 vp_p.n16655 vp_p.n16654 0.013
R17943 vp_p.n16669 vp_p.n16668 0.013
R17944 vp_p.n16683 vp_p.n16682 0.013
R17945 vp_p.n16697 vp_p.n16696 0.013
R17946 vp_p.n16711 vp_p.n16710 0.013
R17947 vp_p.n16725 vp_p.n16724 0.013
R17948 vp_p.n16739 vp_p.n16738 0.013
R17949 vp_p.n16753 vp_p.n16752 0.013
R17950 vp_p.n16767 vp_p.n16766 0.013
R17951 vp_p.n16781 vp_p.n16780 0.013
R17952 vp_p.n16795 vp_p.n16794 0.013
R17953 vp_p.n16809 vp_p.n16808 0.013
R17954 vp_p.n16823 vp_p.n16822 0.013
R17955 vp_p.n16837 vp_p.n16836 0.013
R17956 vp_p.n16851 vp_p.n16850 0.013
R17957 vp_p.n16865 vp_p.n16864 0.013
R17958 vp_p.n16879 vp_p.n16878 0.013
R17959 vp_p.n16893 vp_p.n16892 0.013
R17960 vp_p.n16907 vp_p.n16906 0.013
R17961 vp_p.n16921 vp_p.n16920 0.013
R17962 vp_p.n16935 vp_p.n16934 0.013
R17963 vp_p.n16949 vp_p.n16948 0.013
R17964 vp_p.n16963 vp_p.n16962 0.013
R17965 vp_p.n16977 vp_p.n16976 0.013
R17966 vp_p.n16991 vp_p.n16990 0.013
R17967 vp_p.n17005 vp_p.n17004 0.013
R17968 vp_p.n17019 vp_p.n17018 0.013
R17969 vp_p.n17033 vp_p.n17032 0.013
R17970 vp_p.n17047 vp_p.n17046 0.013
R17971 vp_p.n17061 vp_p.n17060 0.013
R17972 vp_p.n17075 vp_p.n17074 0.013
R17973 vp_p.n17089 vp_p.n17088 0.013
R17974 vp_p.n17103 vp_p.n17102 0.013
R17975 vp_p.n17117 vp_p.n17116 0.013
R17976 vp_p.n17131 vp_p.n17130 0.013
R17977 vp_p.n17145 vp_p.n17144 0.013
R17978 vp_p.n17159 vp_p.n17158 0.013
R17979 vp_p.n17173 vp_p.n17172 0.013
R17980 vp_p.n17187 vp_p.n17186 0.013
R17981 vp_p.n17201 vp_p.n17200 0.013
R17982 vp_p.n17215 vp_p.n17214 0.013
R17983 vp_p.n17229 vp_p.n17228 0.013
R17984 vp_p.n17243 vp_p.n17242 0.013
R17985 vp_p.n17257 vp_p.n17256 0.013
R17986 vp_p.n17261 vp_p.n17260 0.013
R17987 vp_p.n9227 vp_p.n9226 0.013
R17988 vp_p.n9241 vp_p.n9240 0.013
R17989 vp_p.n9255 vp_p.n9254 0.013
R17990 vp_p.n9269 vp_p.n9268 0.013
R17991 vp_p.n9283 vp_p.n9282 0.013
R17992 vp_p.n9297 vp_p.n9296 0.013
R17993 vp_p.n9311 vp_p.n9310 0.013
R17994 vp_p.n9325 vp_p.n9324 0.013
R17995 vp_p.n9339 vp_p.n9338 0.013
R17996 vp_p.n9353 vp_p.n9352 0.013
R17997 vp_p.n9367 vp_p.n9366 0.013
R17998 vp_p.n9381 vp_p.n9380 0.013
R17999 vp_p.n9395 vp_p.n9394 0.013
R18000 vp_p.n9409 vp_p.n9408 0.013
R18001 vp_p.n9423 vp_p.n9422 0.013
R18002 vp_p.n9437 vp_p.n9436 0.013
R18003 vp_p.n9451 vp_p.n9450 0.013
R18004 vp_p.n9465 vp_p.n9464 0.013
R18005 vp_p.n9479 vp_p.n9478 0.013
R18006 vp_p.n9493 vp_p.n9492 0.013
R18007 vp_p.n9507 vp_p.n9506 0.013
R18008 vp_p.n9521 vp_p.n9520 0.013
R18009 vp_p.n9535 vp_p.n9534 0.013
R18010 vp_p.n9549 vp_p.n9548 0.013
R18011 vp_p.n9563 vp_p.n9562 0.013
R18012 vp_p.n9577 vp_p.n9576 0.013
R18013 vp_p.n9591 vp_p.n9590 0.013
R18014 vp_p.n9605 vp_p.n9604 0.013
R18015 vp_p.n9619 vp_p.n9618 0.013
R18016 vp_p.n9633 vp_p.n9632 0.013
R18017 vp_p.n9647 vp_p.n9646 0.013
R18018 vp_p.n9661 vp_p.n9660 0.013
R18019 vp_p.n9675 vp_p.n9674 0.013
R18020 vp_p.n9689 vp_p.n9688 0.013
R18021 vp_p.n9703 vp_p.n9702 0.013
R18022 vp_p.n9717 vp_p.n9716 0.013
R18023 vp_p.n9731 vp_p.n9730 0.013
R18024 vp_p.n9745 vp_p.n9744 0.013
R18025 vp_p.n9759 vp_p.n9758 0.013
R18026 vp_p.n9773 vp_p.n9772 0.013
R18027 vp_p.n9787 vp_p.n9786 0.013
R18028 vp_p.n9801 vp_p.n9800 0.013
R18029 vp_p.n9815 vp_p.n9814 0.013
R18030 vp_p.n9829 vp_p.n9828 0.013
R18031 vp_p.n9843 vp_p.n9842 0.013
R18032 vp_p.n9857 vp_p.n9856 0.013
R18033 vp_p.n9871 vp_p.n9870 0.013
R18034 vp_p.n9885 vp_p.n9884 0.013
R18035 vp_p.n9899 vp_p.n9898 0.013
R18036 vp_p.n9913 vp_p.n9912 0.013
R18037 vp_p.n9927 vp_p.n9926 0.013
R18038 vp_p.n9941 vp_p.n9940 0.013
R18039 vp_p.n9955 vp_p.n9954 0.013
R18040 vp_p.n9969 vp_p.n9968 0.013
R18041 vp_p.n9983 vp_p.n9982 0.013
R18042 vp_p.n9997 vp_p.n9996 0.013
R18043 vp_p.n10011 vp_p.n10010 0.013
R18044 vp_p.n10025 vp_p.n10024 0.013
R18045 vp_p.n10039 vp_p.n10038 0.013
R18046 vp_p.n10053 vp_p.n10052 0.013
R18047 vp_p.n10067 vp_p.n10066 0.013
R18048 vp_p.n10081 vp_p.n10080 0.013
R18049 vp_p.n10095 vp_p.n10094 0.013
R18050 vp_p.n10109 vp_p.n10108 0.013
R18051 vp_p.n10123 vp_p.n10122 0.013
R18052 vp_p.n10137 vp_p.n10136 0.013
R18053 vp_p.n10151 vp_p.n10150 0.013
R18054 vp_p.n10165 vp_p.n10164 0.013
R18055 vp_p.n17760 vp_p.n17759 0.013
R18056 vp_p.n17774 vp_p.n17773 0.013
R18057 vp_p.n17788 vp_p.n17787 0.013
R18058 vp_p.n17802 vp_p.n17801 0.013
R18059 vp_p.n17816 vp_p.n17815 0.013
R18060 vp_p.n17830 vp_p.n17829 0.013
R18061 vp_p.n17844 vp_p.n17843 0.013
R18062 vp_p.n17858 vp_p.n17857 0.013
R18063 vp_p.n17872 vp_p.n17871 0.013
R18064 vp_p.n17886 vp_p.n17885 0.013
R18065 vp_p.n17900 vp_p.n17899 0.013
R18066 vp_p.n17914 vp_p.n17913 0.013
R18067 vp_p.n17928 vp_p.n17927 0.013
R18068 vp_p.n17942 vp_p.n17941 0.013
R18069 vp_p.n17956 vp_p.n17955 0.013
R18070 vp_p.n17970 vp_p.n17969 0.013
R18071 vp_p.n17984 vp_p.n17983 0.013
R18072 vp_p.n17998 vp_p.n17997 0.013
R18073 vp_p.n18012 vp_p.n18011 0.013
R18074 vp_p.n18026 vp_p.n18025 0.013
R18075 vp_p.n18040 vp_p.n18039 0.013
R18076 vp_p.n18054 vp_p.n18053 0.013
R18077 vp_p.n18068 vp_p.n18067 0.013
R18078 vp_p.n18082 vp_p.n18081 0.013
R18079 vp_p.n18096 vp_p.n18095 0.013
R18080 vp_p.n18110 vp_p.n18109 0.013
R18081 vp_p.n18124 vp_p.n18123 0.013
R18082 vp_p.n18138 vp_p.n18137 0.013
R18083 vp_p.n18152 vp_p.n18151 0.013
R18084 vp_p.n18166 vp_p.n18165 0.013
R18085 vp_p.n18180 vp_p.n18179 0.013
R18086 vp_p.n18194 vp_p.n18193 0.013
R18087 vp_p.n18208 vp_p.n18207 0.013
R18088 vp_p.n18222 vp_p.n18221 0.013
R18089 vp_p.n18236 vp_p.n18235 0.013
R18090 vp_p.n18250 vp_p.n18249 0.013
R18091 vp_p.n18264 vp_p.n18263 0.013
R18092 vp_p.n18278 vp_p.n18277 0.013
R18093 vp_p.n18292 vp_p.n18291 0.013
R18094 vp_p.n18306 vp_p.n18305 0.013
R18095 vp_p.n18320 vp_p.n18319 0.013
R18096 vp_p.n18334 vp_p.n18333 0.013
R18097 vp_p.n18348 vp_p.n18347 0.013
R18098 vp_p.n18362 vp_p.n18361 0.013
R18099 vp_p.n18376 vp_p.n18375 0.013
R18100 vp_p.n18390 vp_p.n18389 0.013
R18101 vp_p.n18404 vp_p.n18403 0.013
R18102 vp_p.n18418 vp_p.n18417 0.013
R18103 vp_p.n18432 vp_p.n18431 0.013
R18104 vp_p.n18446 vp_p.n18445 0.013
R18105 vp_p.n18460 vp_p.n18459 0.013
R18106 vp_p.n18474 vp_p.n18473 0.013
R18107 vp_p.n18488 vp_p.n18487 0.013
R18108 vp_p.n18502 vp_p.n18501 0.013
R18109 vp_p.n18516 vp_p.n18515 0.013
R18110 vp_p.n18530 vp_p.n18529 0.013
R18111 vp_p.n18544 vp_p.n18543 0.013
R18112 vp_p.n18558 vp_p.n18557 0.013
R18113 vp_p.n18572 vp_p.n18571 0.013
R18114 vp_p.n18586 vp_p.n18585 0.013
R18115 vp_p.n18600 vp_p.n18599 0.013
R18116 vp_p.n18614 vp_p.n18613 0.013
R18117 vp_p.n18628 vp_p.n18627 0.013
R18118 vp_p.n18642 vp_p.n18641 0.013
R18119 vp_p.n18656 vp_p.n18655 0.013
R18120 vp_p.n18670 vp_p.n18669 0.013
R18121 vp_p.n18684 vp_p.n18683 0.013
R18122 vp_p.n18698 vp_p.n18697 0.013
R18123 vp_p.n18702 vp_p.n18701 0.013
R18124 vp_p.n481 vp_p.n480 0.013
R18125 vp_p.n495 vp_p.n494 0.013
R18126 vp_p.n509 vp_p.n508 0.013
R18127 vp_p.n523 vp_p.n522 0.013
R18128 vp_p.n537 vp_p.n536 0.013
R18129 vp_p.n551 vp_p.n550 0.013
R18130 vp_p.n565 vp_p.n564 0.013
R18131 vp_p.n579 vp_p.n578 0.013
R18132 vp_p.n593 vp_p.n592 0.013
R18133 vp_p.n607 vp_p.n606 0.013
R18134 vp_p.n621 vp_p.n620 0.013
R18135 vp_p.n635 vp_p.n634 0.013
R18136 vp_p.n649 vp_p.n648 0.013
R18137 vp_p.n663 vp_p.n662 0.013
R18138 vp_p.n677 vp_p.n676 0.013
R18139 vp_p.n691 vp_p.n690 0.013
R18140 vp_p.n705 vp_p.n704 0.013
R18141 vp_p.n719 vp_p.n718 0.013
R18142 vp_p.n733 vp_p.n732 0.013
R18143 vp_p.n747 vp_p.n746 0.013
R18144 vp_p.n761 vp_p.n760 0.013
R18145 vp_p.n775 vp_p.n774 0.013
R18146 vp_p.n789 vp_p.n788 0.013
R18147 vp_p.n803 vp_p.n802 0.013
R18148 vp_p.n817 vp_p.n816 0.013
R18149 vp_p.n831 vp_p.n830 0.013
R18150 vp_p.n845 vp_p.n844 0.013
R18151 vp_p.n859 vp_p.n858 0.013
R18152 vp_p.n873 vp_p.n872 0.013
R18153 vp_p.n887 vp_p.n886 0.013
R18154 vp_p.n901 vp_p.n900 0.013
R18155 vp_p.n915 vp_p.n914 0.013
R18156 vp_p.n929 vp_p.n928 0.013
R18157 vp_p.n943 vp_p.n942 0.013
R18158 vp_p.n957 vp_p.n956 0.013
R18159 vp_p.n971 vp_p.n970 0.013
R18160 vp_p.n985 vp_p.n984 0.013
R18161 vp_p.n999 vp_p.n998 0.013
R18162 vp_p.n1013 vp_p.n1012 0.013
R18163 vp_p.n1027 vp_p.n1026 0.013
R18164 vp_p.n1041 vp_p.n1040 0.013
R18165 vp_p.n1055 vp_p.n1054 0.013
R18166 vp_p.n1069 vp_p.n1068 0.013
R18167 vp_p.n1083 vp_p.n1082 0.013
R18168 vp_p.n1097 vp_p.n1096 0.013
R18169 vp_p.n1111 vp_p.n1110 0.013
R18170 vp_p.n1125 vp_p.n1124 0.013
R18171 vp_p.n1139 vp_p.n1138 0.013
R18172 vp_p.n1153 vp_p.n1152 0.013
R18173 vp_p.n1167 vp_p.n1166 0.013
R18174 vp_p.n1181 vp_p.n1180 0.013
R18175 vp_p.n1195 vp_p.n1194 0.013
R18176 vp_p.n1209 vp_p.n1208 0.013
R18177 vp_p.n1223 vp_p.n1222 0.013
R18178 vp_p.n1237 vp_p.n1236 0.013
R18179 vp_p.n1251 vp_p.n1250 0.013
R18180 vp_p.n1265 vp_p.n1264 0.013
R18181 vp_p.n1279 vp_p.n1278 0.013
R18182 vp_p.n1293 vp_p.n1292 0.013
R18183 vp_p.n1307 vp_p.n1306 0.013
R18184 vp_p.n1321 vp_p.n1320 0.013
R18185 vp_p.n1335 vp_p.n1334 0.013
R18186 vp_p.n1349 vp_p.n1348 0.013
R18187 vp_p.n1363 vp_p.n1362 0.013
R18188 vp_p.n1377 vp_p.n1376 0.013
R18189 vp_p.n1391 vp_p.n1390 0.013
R18190 vp_p.n1405 vp_p.n1404 0.013
R18191 vp_p.n1419 vp_p.n1418 0.013
R18192 vp_p.n1433 vp_p.n1432 0.013
R18193 vp_p.n19186 vp_p.n19185 0.013
R18194 vp_p.n19200 vp_p.n19199 0.013
R18195 vp_p.n19214 vp_p.n19213 0.013
R18196 vp_p.n19228 vp_p.n19227 0.013
R18197 vp_p.n19242 vp_p.n19241 0.013
R18198 vp_p.n19256 vp_p.n19255 0.013
R18199 vp_p.n19270 vp_p.n19269 0.013
R18200 vp_p.n19284 vp_p.n19283 0.013
R18201 vp_p.n19298 vp_p.n19297 0.013
R18202 vp_p.n19312 vp_p.n19311 0.013
R18203 vp_p.n19326 vp_p.n19325 0.013
R18204 vp_p.n19340 vp_p.n19339 0.013
R18205 vp_p.n19354 vp_p.n19353 0.013
R18206 vp_p.n19368 vp_p.n19367 0.013
R18207 vp_p.n19382 vp_p.n19381 0.013
R18208 vp_p.n19396 vp_p.n19395 0.013
R18209 vp_p.n19410 vp_p.n19409 0.013
R18210 vp_p.n19424 vp_p.n19423 0.013
R18211 vp_p.n19438 vp_p.n19437 0.013
R18212 vp_p.n19452 vp_p.n19451 0.013
R18213 vp_p.n19466 vp_p.n19465 0.013
R18214 vp_p.n19480 vp_p.n19479 0.013
R18215 vp_p.n19494 vp_p.n19493 0.013
R18216 vp_p.n19508 vp_p.n19507 0.013
R18217 vp_p.n19522 vp_p.n19521 0.013
R18218 vp_p.n19536 vp_p.n19535 0.013
R18219 vp_p.n19550 vp_p.n19549 0.013
R18220 vp_p.n19564 vp_p.n19563 0.013
R18221 vp_p.n19578 vp_p.n19577 0.013
R18222 vp_p.n19592 vp_p.n19591 0.013
R18223 vp_p.n19606 vp_p.n19605 0.013
R18224 vp_p.n19620 vp_p.n19619 0.013
R18225 vp_p.n19634 vp_p.n19633 0.013
R18226 vp_p.n19648 vp_p.n19647 0.013
R18227 vp_p.n19662 vp_p.n19661 0.013
R18228 vp_p.n19676 vp_p.n19675 0.013
R18229 vp_p.n19690 vp_p.n19689 0.013
R18230 vp_p.n19704 vp_p.n19703 0.013
R18231 vp_p.n19718 vp_p.n19717 0.013
R18232 vp_p.n19732 vp_p.n19731 0.013
R18233 vp_p.n19746 vp_p.n19745 0.013
R18234 vp_p.n19760 vp_p.n19759 0.013
R18235 vp_p.n19774 vp_p.n19773 0.013
R18236 vp_p.n19788 vp_p.n19787 0.013
R18237 vp_p.n19802 vp_p.n19801 0.013
R18238 vp_p.n19816 vp_p.n19815 0.013
R18239 vp_p.n19830 vp_p.n19829 0.013
R18240 vp_p.n19844 vp_p.n19843 0.013
R18241 vp_p.n19858 vp_p.n19857 0.013
R18242 vp_p.n19872 vp_p.n19871 0.013
R18243 vp_p.n19886 vp_p.n19885 0.013
R18244 vp_p.n19900 vp_p.n19899 0.013
R18245 vp_p.n19914 vp_p.n19913 0.013
R18246 vp_p.n19928 vp_p.n19927 0.013
R18247 vp_p.n19942 vp_p.n19941 0.013
R18248 vp_p.n19956 vp_p.n19955 0.013
R18249 vp_p.n19970 vp_p.n19969 0.013
R18250 vp_p.n19984 vp_p.n19983 0.013
R18251 vp_p.n19998 vp_p.n19997 0.013
R18252 vp_p.n20012 vp_p.n20011 0.013
R18253 vp_p.n20026 vp_p.n20025 0.013
R18254 vp_p.n20040 vp_p.n20039 0.013
R18255 vp_p.n20054 vp_p.n20053 0.013
R18256 vp_p.n20068 vp_p.n20067 0.013
R18257 vp_p.n20082 vp_p.n20081 0.013
R18258 vp_p.n20096 vp_p.n20095 0.013
R18259 vp_p.n20110 vp_p.n20109 0.013
R18260 vp_p.n20124 vp_p.n20123 0.013
R18261 vp_p.n20138 vp_p.n20137 0.013
R18262 vp_p.n20142 vp_p.n20141 0.013
R18263 vp_p.n1907 vp_p.n1906 0.013
R18264 vp_p.n1921 vp_p.n1920 0.013
R18265 vp_p.n1935 vp_p.n1934 0.013
R18266 vp_p.n1949 vp_p.n1948 0.013
R18267 vp_p.n1963 vp_p.n1962 0.013
R18268 vp_p.n1977 vp_p.n1976 0.013
R18269 vp_p.n1991 vp_p.n1990 0.013
R18270 vp_p.n2005 vp_p.n2004 0.013
R18271 vp_p.n2019 vp_p.n2018 0.013
R18272 vp_p.n2033 vp_p.n2032 0.013
R18273 vp_p.n2047 vp_p.n2046 0.013
R18274 vp_p.n2061 vp_p.n2060 0.013
R18275 vp_p.n2075 vp_p.n2074 0.013
R18276 vp_p.n2089 vp_p.n2088 0.013
R18277 vp_p.n2103 vp_p.n2102 0.013
R18278 vp_p.n2117 vp_p.n2116 0.013
R18279 vp_p.n2131 vp_p.n2130 0.013
R18280 vp_p.n2145 vp_p.n2144 0.013
R18281 vp_p.n2159 vp_p.n2158 0.013
R18282 vp_p.n2173 vp_p.n2172 0.013
R18283 vp_p.n2187 vp_p.n2186 0.013
R18284 vp_p.n2201 vp_p.n2200 0.013
R18285 vp_p.n2215 vp_p.n2214 0.013
R18286 vp_p.n2229 vp_p.n2228 0.013
R18287 vp_p.n2243 vp_p.n2242 0.013
R18288 vp_p.n2257 vp_p.n2256 0.013
R18289 vp_p.n2271 vp_p.n2270 0.013
R18290 vp_p.n2285 vp_p.n2284 0.013
R18291 vp_p.n2299 vp_p.n2298 0.013
R18292 vp_p.n2313 vp_p.n2312 0.013
R18293 vp_p.n2327 vp_p.n2326 0.013
R18294 vp_p.n2341 vp_p.n2340 0.013
R18295 vp_p.n2355 vp_p.n2354 0.013
R18296 vp_p.n2369 vp_p.n2368 0.013
R18297 vp_p.n2383 vp_p.n2382 0.013
R18298 vp_p.n2397 vp_p.n2396 0.013
R18299 vp_p.n2411 vp_p.n2410 0.013
R18300 vp_p.n2425 vp_p.n2424 0.013
R18301 vp_p.n2439 vp_p.n2438 0.013
R18302 vp_p.n2453 vp_p.n2452 0.013
R18303 vp_p.n2467 vp_p.n2466 0.013
R18304 vp_p.n2481 vp_p.n2480 0.013
R18305 vp_p.n2495 vp_p.n2494 0.013
R18306 vp_p.n2509 vp_p.n2508 0.013
R18307 vp_p.n2523 vp_p.n2522 0.013
R18308 vp_p.n2537 vp_p.n2536 0.013
R18309 vp_p.n2551 vp_p.n2550 0.013
R18310 vp_p.n2565 vp_p.n2564 0.013
R18311 vp_p.n2579 vp_p.n2578 0.013
R18312 vp_p.n2593 vp_p.n2592 0.013
R18313 vp_p.n2607 vp_p.n2606 0.013
R18314 vp_p.n2621 vp_p.n2620 0.013
R18315 vp_p.n2635 vp_p.n2634 0.013
R18316 vp_p.n2649 vp_p.n2648 0.013
R18317 vp_p.n2663 vp_p.n2662 0.013
R18318 vp_p.n2677 vp_p.n2676 0.013
R18319 vp_p.n2691 vp_p.n2690 0.013
R18320 vp_p.n2705 vp_p.n2704 0.013
R18321 vp_p.n2719 vp_p.n2718 0.013
R18322 vp_p.n2733 vp_p.n2732 0.013
R18323 vp_p.n2747 vp_p.n2746 0.013
R18324 vp_p.n2761 vp_p.n2760 0.013
R18325 vp_p.n2775 vp_p.n2774 0.013
R18326 vp_p.n2789 vp_p.n2788 0.013
R18327 vp_p.n2803 vp_p.n2802 0.013
R18328 vp_p.n2817 vp_p.n2816 0.013
R18329 vp_p.n2831 vp_p.n2830 0.013
R18330 vp_p.n2845 vp_p.n2844 0.013
R18331 vp_p.n2859 vp_p.n2858 0.013
R18332 vp_p.n2873 vp_p.n2872 0.013
R18333 vp_p.n20611 vp_p.n20610 0.013
R18334 vp_p.n20625 vp_p.n20624 0.013
R18335 vp_p.n20639 vp_p.n20638 0.013
R18336 vp_p.n20653 vp_p.n20652 0.013
R18337 vp_p.n20667 vp_p.n20666 0.013
R18338 vp_p.n20681 vp_p.n20680 0.013
R18339 vp_p.n20695 vp_p.n20694 0.013
R18340 vp_p.n20709 vp_p.n20708 0.013
R18341 vp_p.n20723 vp_p.n20722 0.013
R18342 vp_p.n20737 vp_p.n20736 0.013
R18343 vp_p.n20751 vp_p.n20750 0.013
R18344 vp_p.n20765 vp_p.n20764 0.013
R18345 vp_p.n20779 vp_p.n20778 0.013
R18346 vp_p.n20793 vp_p.n20792 0.013
R18347 vp_p.n20807 vp_p.n20806 0.013
R18348 vp_p.n20821 vp_p.n20820 0.013
R18349 vp_p.n20835 vp_p.n20834 0.013
R18350 vp_p.n20849 vp_p.n20848 0.013
R18351 vp_p.n20863 vp_p.n20862 0.013
R18352 vp_p.n20877 vp_p.n20876 0.013
R18353 vp_p.n20891 vp_p.n20890 0.013
R18354 vp_p.n20905 vp_p.n20904 0.013
R18355 vp_p.n20919 vp_p.n20918 0.013
R18356 vp_p.n20933 vp_p.n20932 0.013
R18357 vp_p.n20947 vp_p.n20946 0.013
R18358 vp_p.n20961 vp_p.n20960 0.013
R18359 vp_p.n20975 vp_p.n20974 0.013
R18360 vp_p.n20989 vp_p.n20988 0.013
R18361 vp_p.n21003 vp_p.n21002 0.013
R18362 vp_p.n21017 vp_p.n21016 0.013
R18363 vp_p.n21031 vp_p.n21030 0.013
R18364 vp_p.n21045 vp_p.n21044 0.013
R18365 vp_p.n21059 vp_p.n21058 0.013
R18366 vp_p.n21073 vp_p.n21072 0.013
R18367 vp_p.n21087 vp_p.n21086 0.013
R18368 vp_p.n21101 vp_p.n21100 0.013
R18369 vp_p.n21115 vp_p.n21114 0.013
R18370 vp_p.n21129 vp_p.n21128 0.013
R18371 vp_p.n21143 vp_p.n21142 0.013
R18372 vp_p.n21157 vp_p.n21156 0.013
R18373 vp_p.n21171 vp_p.n21170 0.013
R18374 vp_p.n21185 vp_p.n21184 0.013
R18375 vp_p.n21199 vp_p.n21198 0.013
R18376 vp_p.n21213 vp_p.n21212 0.013
R18377 vp_p.n21227 vp_p.n21226 0.013
R18378 vp_p.n21241 vp_p.n21240 0.013
R18379 vp_p.n21255 vp_p.n21254 0.013
R18380 vp_p.n21269 vp_p.n21268 0.013
R18381 vp_p.n21283 vp_p.n21282 0.013
R18382 vp_p.n21297 vp_p.n21296 0.013
R18383 vp_p.n21311 vp_p.n21310 0.013
R18384 vp_p.n21325 vp_p.n21324 0.013
R18385 vp_p.n21339 vp_p.n21338 0.013
R18386 vp_p.n21353 vp_p.n21352 0.013
R18387 vp_p.n21367 vp_p.n21366 0.013
R18388 vp_p.n21381 vp_p.n21380 0.013
R18389 vp_p.n21395 vp_p.n21394 0.013
R18390 vp_p.n21409 vp_p.n21408 0.013
R18391 vp_p.n21423 vp_p.n21422 0.013
R18392 vp_p.n21437 vp_p.n21436 0.013
R18393 vp_p.n21451 vp_p.n21450 0.013
R18394 vp_p.n21465 vp_p.n21464 0.013
R18395 vp_p.n21479 vp_p.n21478 0.013
R18396 vp_p.n21493 vp_p.n21492 0.013
R18397 vp_p.n21507 vp_p.n21506 0.013
R18398 vp_p.n21521 vp_p.n21520 0.013
R18399 vp_p.n21535 vp_p.n21534 0.013
R18400 vp_p.n21549 vp_p.n21548 0.013
R18401 vp_p.n21563 vp_p.n21562 0.013
R18402 vp_p.n21577 vp_p.n21576 0.013
R18403 vp_p.n21581 vp_p.n21580 0.013
R18404 vp_p.n3332 vp_p.n3331 0.013
R18405 vp_p.n3346 vp_p.n3345 0.013
R18406 vp_p.n3360 vp_p.n3359 0.013
R18407 vp_p.n3374 vp_p.n3373 0.013
R18408 vp_p.n3388 vp_p.n3387 0.013
R18409 vp_p.n3402 vp_p.n3401 0.013
R18410 vp_p.n3416 vp_p.n3415 0.013
R18411 vp_p.n3430 vp_p.n3429 0.013
R18412 vp_p.n3444 vp_p.n3443 0.013
R18413 vp_p.n3458 vp_p.n3457 0.013
R18414 vp_p.n3472 vp_p.n3471 0.013
R18415 vp_p.n3486 vp_p.n3485 0.013
R18416 vp_p.n3500 vp_p.n3499 0.013
R18417 vp_p.n3514 vp_p.n3513 0.013
R18418 vp_p.n3528 vp_p.n3527 0.013
R18419 vp_p.n3542 vp_p.n3541 0.013
R18420 vp_p.n3556 vp_p.n3555 0.013
R18421 vp_p.n3570 vp_p.n3569 0.013
R18422 vp_p.n3584 vp_p.n3583 0.013
R18423 vp_p.n3598 vp_p.n3597 0.013
R18424 vp_p.n3612 vp_p.n3611 0.013
R18425 vp_p.n3626 vp_p.n3625 0.013
R18426 vp_p.n3640 vp_p.n3639 0.013
R18427 vp_p.n3654 vp_p.n3653 0.013
R18428 vp_p.n3668 vp_p.n3667 0.013
R18429 vp_p.n3682 vp_p.n3681 0.013
R18430 vp_p.n3696 vp_p.n3695 0.013
R18431 vp_p.n3710 vp_p.n3709 0.013
R18432 vp_p.n3724 vp_p.n3723 0.013
R18433 vp_p.n3738 vp_p.n3737 0.013
R18434 vp_p.n3752 vp_p.n3751 0.013
R18435 vp_p.n3766 vp_p.n3765 0.013
R18436 vp_p.n3780 vp_p.n3779 0.013
R18437 vp_p.n3794 vp_p.n3793 0.013
R18438 vp_p.n3808 vp_p.n3807 0.013
R18439 vp_p.n3822 vp_p.n3821 0.013
R18440 vp_p.n3836 vp_p.n3835 0.013
R18441 vp_p.n3850 vp_p.n3849 0.013
R18442 vp_p.n3864 vp_p.n3863 0.013
R18443 vp_p.n3878 vp_p.n3877 0.013
R18444 vp_p.n3892 vp_p.n3891 0.013
R18445 vp_p.n3906 vp_p.n3905 0.013
R18446 vp_p.n3920 vp_p.n3919 0.013
R18447 vp_p.n3934 vp_p.n3933 0.013
R18448 vp_p.n3948 vp_p.n3947 0.013
R18449 vp_p.n3962 vp_p.n3961 0.013
R18450 vp_p.n3976 vp_p.n3975 0.013
R18451 vp_p.n3990 vp_p.n3989 0.013
R18452 vp_p.n4004 vp_p.n4003 0.013
R18453 vp_p.n4018 vp_p.n4017 0.013
R18454 vp_p.n4032 vp_p.n4031 0.013
R18455 vp_p.n4046 vp_p.n4045 0.013
R18456 vp_p.n4060 vp_p.n4059 0.013
R18457 vp_p.n4074 vp_p.n4073 0.013
R18458 vp_p.n4088 vp_p.n4087 0.013
R18459 vp_p.n4102 vp_p.n4101 0.013
R18460 vp_p.n4116 vp_p.n4115 0.013
R18461 vp_p.n4130 vp_p.n4129 0.013
R18462 vp_p.n4144 vp_p.n4143 0.013
R18463 vp_p.n4158 vp_p.n4157 0.013
R18464 vp_p.n4172 vp_p.n4171 0.013
R18465 vp_p.n4186 vp_p.n4185 0.013
R18466 vp_p.n4200 vp_p.n4199 0.013
R18467 vp_p.n4214 vp_p.n4213 0.013
R18468 vp_p.n4228 vp_p.n4227 0.013
R18469 vp_p.n4242 vp_p.n4241 0.013
R18470 vp_p.n4256 vp_p.n4255 0.013
R18471 vp_p.n4270 vp_p.n4269 0.013
R18472 vp_p.n4284 vp_p.n4283 0.013
R18473 vp_p.n4298 vp_p.n4297 0.013
R18474 vp_p.n4312 vp_p.n4311 0.013
R18475 vp_p.n22035 vp_p.n22034 0.013
R18476 vp_p.n22049 vp_p.n22048 0.013
R18477 vp_p.n22063 vp_p.n22062 0.013
R18478 vp_p.n22077 vp_p.n22076 0.013
R18479 vp_p.n22091 vp_p.n22090 0.013
R18480 vp_p.n22105 vp_p.n22104 0.013
R18481 vp_p.n22119 vp_p.n22118 0.013
R18482 vp_p.n22133 vp_p.n22132 0.013
R18483 vp_p.n22147 vp_p.n22146 0.013
R18484 vp_p.n22161 vp_p.n22160 0.013
R18485 vp_p.n22175 vp_p.n22174 0.013
R18486 vp_p.n22189 vp_p.n22188 0.013
R18487 vp_p.n22203 vp_p.n22202 0.013
R18488 vp_p.n22217 vp_p.n22216 0.013
R18489 vp_p.n22231 vp_p.n22230 0.013
R18490 vp_p.n22245 vp_p.n22244 0.013
R18491 vp_p.n22259 vp_p.n22258 0.013
R18492 vp_p.n22273 vp_p.n22272 0.013
R18493 vp_p.n22287 vp_p.n22286 0.013
R18494 vp_p.n22301 vp_p.n22300 0.013
R18495 vp_p.n22315 vp_p.n22314 0.013
R18496 vp_p.n22329 vp_p.n22328 0.013
R18497 vp_p.n22343 vp_p.n22342 0.013
R18498 vp_p.n22357 vp_p.n22356 0.013
R18499 vp_p.n22371 vp_p.n22370 0.013
R18500 vp_p.n22385 vp_p.n22384 0.013
R18501 vp_p.n22399 vp_p.n22398 0.013
R18502 vp_p.n22413 vp_p.n22412 0.013
R18503 vp_p.n22427 vp_p.n22426 0.013
R18504 vp_p.n22441 vp_p.n22440 0.013
R18505 vp_p.n22455 vp_p.n22454 0.013
R18506 vp_p.n22469 vp_p.n22468 0.013
R18507 vp_p.n22483 vp_p.n22482 0.013
R18508 vp_p.n22497 vp_p.n22496 0.013
R18509 vp_p.n22511 vp_p.n22510 0.013
R18510 vp_p.n22525 vp_p.n22524 0.013
R18511 vp_p.n22539 vp_p.n22538 0.013
R18512 vp_p.n22553 vp_p.n22552 0.013
R18513 vp_p.n22567 vp_p.n22566 0.013
R18514 vp_p.n22581 vp_p.n22580 0.013
R18515 vp_p.n22595 vp_p.n22594 0.013
R18516 vp_p.n22609 vp_p.n22608 0.013
R18517 vp_p.n22623 vp_p.n22622 0.013
R18518 vp_p.n22637 vp_p.n22636 0.013
R18519 vp_p.n22651 vp_p.n22650 0.013
R18520 vp_p.n22665 vp_p.n22664 0.013
R18521 vp_p.n22679 vp_p.n22678 0.013
R18522 vp_p.n22693 vp_p.n22692 0.013
R18523 vp_p.n22707 vp_p.n22706 0.013
R18524 vp_p.n22721 vp_p.n22720 0.013
R18525 vp_p.n22735 vp_p.n22734 0.013
R18526 vp_p.n22749 vp_p.n22748 0.013
R18527 vp_p.n22763 vp_p.n22762 0.013
R18528 vp_p.n22777 vp_p.n22776 0.013
R18529 vp_p.n22791 vp_p.n22790 0.013
R18530 vp_p.n22805 vp_p.n22804 0.013
R18531 vp_p.n22819 vp_p.n22818 0.013
R18532 vp_p.n22833 vp_p.n22832 0.013
R18533 vp_p.n22847 vp_p.n22846 0.013
R18534 vp_p.n22861 vp_p.n22860 0.013
R18535 vp_p.n22875 vp_p.n22874 0.013
R18536 vp_p.n22889 vp_p.n22888 0.013
R18537 vp_p.n22903 vp_p.n22902 0.013
R18538 vp_p.n22917 vp_p.n22916 0.013
R18539 vp_p.n22931 vp_p.n22930 0.013
R18540 vp_p.n22945 vp_p.n22944 0.013
R18541 vp_p.n22959 vp_p.n22958 0.013
R18542 vp_p.n22973 vp_p.n22972 0.013
R18543 vp_p.n22987 vp_p.n22986 0.013
R18544 vp_p.n23001 vp_p.n23000 0.013
R18545 vp_p.n23015 vp_p.n23014 0.013
R18546 vp_p.n23019 vp_p.n23018 0.013
R18547 vp_p.n4756 vp_p.n4755 0.013
R18548 vp_p.n4770 vp_p.n4769 0.013
R18549 vp_p.n4784 vp_p.n4783 0.013
R18550 vp_p.n4798 vp_p.n4797 0.013
R18551 vp_p.n4812 vp_p.n4811 0.013
R18552 vp_p.n4826 vp_p.n4825 0.013
R18553 vp_p.n4840 vp_p.n4839 0.013
R18554 vp_p.n4854 vp_p.n4853 0.013
R18555 vp_p.n4868 vp_p.n4867 0.013
R18556 vp_p.n4882 vp_p.n4881 0.013
R18557 vp_p.n4896 vp_p.n4895 0.013
R18558 vp_p.n4910 vp_p.n4909 0.013
R18559 vp_p.n4924 vp_p.n4923 0.013
R18560 vp_p.n4938 vp_p.n4937 0.013
R18561 vp_p.n4952 vp_p.n4951 0.013
R18562 vp_p.n4966 vp_p.n4965 0.013
R18563 vp_p.n4980 vp_p.n4979 0.013
R18564 vp_p.n4994 vp_p.n4993 0.013
R18565 vp_p.n5008 vp_p.n5007 0.013
R18566 vp_p.n5022 vp_p.n5021 0.013
R18567 vp_p.n5036 vp_p.n5035 0.013
R18568 vp_p.n5050 vp_p.n5049 0.013
R18569 vp_p.n5064 vp_p.n5063 0.013
R18570 vp_p.n5078 vp_p.n5077 0.013
R18571 vp_p.n5092 vp_p.n5091 0.013
R18572 vp_p.n5106 vp_p.n5105 0.013
R18573 vp_p.n5120 vp_p.n5119 0.013
R18574 vp_p.n5134 vp_p.n5133 0.013
R18575 vp_p.n5148 vp_p.n5147 0.013
R18576 vp_p.n5162 vp_p.n5161 0.013
R18577 vp_p.n5176 vp_p.n5175 0.013
R18578 vp_p.n5190 vp_p.n5189 0.013
R18579 vp_p.n5204 vp_p.n5203 0.013
R18580 vp_p.n5218 vp_p.n5217 0.013
R18581 vp_p.n5232 vp_p.n5231 0.013
R18582 vp_p.n5246 vp_p.n5245 0.013
R18583 vp_p.n5260 vp_p.n5259 0.013
R18584 vp_p.n5274 vp_p.n5273 0.013
R18585 vp_p.n5288 vp_p.n5287 0.013
R18586 vp_p.n5302 vp_p.n5301 0.013
R18587 vp_p.n5316 vp_p.n5315 0.013
R18588 vp_p.n5330 vp_p.n5329 0.013
R18589 vp_p.n5344 vp_p.n5343 0.013
R18590 vp_p.n5358 vp_p.n5357 0.013
R18591 vp_p.n5372 vp_p.n5371 0.013
R18592 vp_p.n5386 vp_p.n5385 0.013
R18593 vp_p.n5400 vp_p.n5399 0.013
R18594 vp_p.n5414 vp_p.n5413 0.013
R18595 vp_p.n5428 vp_p.n5427 0.013
R18596 vp_p.n5442 vp_p.n5441 0.013
R18597 vp_p.n5456 vp_p.n5455 0.013
R18598 vp_p.n5470 vp_p.n5469 0.013
R18599 vp_p.n5484 vp_p.n5483 0.013
R18600 vp_p.n5498 vp_p.n5497 0.013
R18601 vp_p.n5512 vp_p.n5511 0.013
R18602 vp_p.n5526 vp_p.n5525 0.013
R18603 vp_p.n5540 vp_p.n5539 0.013
R18604 vp_p.n5554 vp_p.n5553 0.013
R18605 vp_p.n5568 vp_p.n5567 0.013
R18606 vp_p.n5582 vp_p.n5581 0.013
R18607 vp_p.n5596 vp_p.n5595 0.013
R18608 vp_p.n5610 vp_p.n5609 0.013
R18609 vp_p.n5624 vp_p.n5623 0.013
R18610 vp_p.n5638 vp_p.n5637 0.013
R18611 vp_p.n5652 vp_p.n5651 0.013
R18612 vp_p.n5666 vp_p.n5665 0.013
R18613 vp_p.n5680 vp_p.n5679 0.013
R18614 vp_p.n5694 vp_p.n5693 0.013
R18615 vp_p.n5708 vp_p.n5707 0.013
R18616 vp_p.n5722 vp_p.n5721 0.013
R18617 vp_p.n5736 vp_p.n5735 0.013
R18618 vp_p.n5750 vp_p.n5749 0.013
R18619 vp_p.n23458 vp_p.n23457 0.013
R18620 vp_p.n23472 vp_p.n23471 0.013
R18621 vp_p.n23486 vp_p.n23485 0.013
R18622 vp_p.n23500 vp_p.n23499 0.013
R18623 vp_p.n23514 vp_p.n23513 0.013
R18624 vp_p.n23528 vp_p.n23527 0.013
R18625 vp_p.n23542 vp_p.n23541 0.013
R18626 vp_p.n23556 vp_p.n23555 0.013
R18627 vp_p.n23570 vp_p.n23569 0.013
R18628 vp_p.n23584 vp_p.n23583 0.013
R18629 vp_p.n23598 vp_p.n23597 0.013
R18630 vp_p.n23612 vp_p.n23611 0.013
R18631 vp_p.n23626 vp_p.n23625 0.013
R18632 vp_p.n23640 vp_p.n23639 0.013
R18633 vp_p.n23654 vp_p.n23653 0.013
R18634 vp_p.n23668 vp_p.n23667 0.013
R18635 vp_p.n23682 vp_p.n23681 0.013
R18636 vp_p.n23696 vp_p.n23695 0.013
R18637 vp_p.n23710 vp_p.n23709 0.013
R18638 vp_p.n23724 vp_p.n23723 0.013
R18639 vp_p.n23738 vp_p.n23737 0.013
R18640 vp_p.n23752 vp_p.n23751 0.013
R18641 vp_p.n23766 vp_p.n23765 0.013
R18642 vp_p.n23780 vp_p.n23779 0.013
R18643 vp_p.n23794 vp_p.n23793 0.013
R18644 vp_p.n23808 vp_p.n23807 0.013
R18645 vp_p.n23822 vp_p.n23821 0.013
R18646 vp_p.n23836 vp_p.n23835 0.013
R18647 vp_p.n23850 vp_p.n23849 0.013
R18648 vp_p.n23864 vp_p.n23863 0.013
R18649 vp_p.n23878 vp_p.n23877 0.013
R18650 vp_p.n23892 vp_p.n23891 0.013
R18651 vp_p.n23906 vp_p.n23905 0.013
R18652 vp_p.n23920 vp_p.n23919 0.013
R18653 vp_p.n23934 vp_p.n23933 0.013
R18654 vp_p.n23948 vp_p.n23947 0.013
R18655 vp_p.n23962 vp_p.n23961 0.013
R18656 vp_p.n23976 vp_p.n23975 0.013
R18657 vp_p.n23990 vp_p.n23989 0.013
R18658 vp_p.n24004 vp_p.n24003 0.013
R18659 vp_p.n24018 vp_p.n24017 0.013
R18660 vp_p.n24032 vp_p.n24031 0.013
R18661 vp_p.n24046 vp_p.n24045 0.013
R18662 vp_p.n24060 vp_p.n24059 0.013
R18663 vp_p.n24074 vp_p.n24073 0.013
R18664 vp_p.n24088 vp_p.n24087 0.013
R18665 vp_p.n24102 vp_p.n24101 0.013
R18666 vp_p.n24116 vp_p.n24115 0.013
R18667 vp_p.n24130 vp_p.n24129 0.013
R18668 vp_p.n24144 vp_p.n24143 0.013
R18669 vp_p.n24158 vp_p.n24157 0.013
R18670 vp_p.n24172 vp_p.n24171 0.013
R18671 vp_p.n24186 vp_p.n24185 0.013
R18672 vp_p.n24200 vp_p.n24199 0.013
R18673 vp_p.n24214 vp_p.n24213 0.013
R18674 vp_p.n24228 vp_p.n24227 0.013
R18675 vp_p.n24242 vp_p.n24241 0.013
R18676 vp_p.n24256 vp_p.n24255 0.013
R18677 vp_p.n24270 vp_p.n24269 0.013
R18678 vp_p.n24284 vp_p.n24283 0.013
R18679 vp_p.n24298 vp_p.n24297 0.013
R18680 vp_p.n24312 vp_p.n24311 0.013
R18681 vp_p.n24326 vp_p.n24325 0.013
R18682 vp_p.n24340 vp_p.n24339 0.013
R18683 vp_p.n24354 vp_p.n24353 0.013
R18684 vp_p.n24368 vp_p.n24367 0.013
R18685 vp_p.n24382 vp_p.n24381 0.013
R18686 vp_p.n24396 vp_p.n24395 0.013
R18687 vp_p.n24410 vp_p.n24409 0.013
R18688 vp_p.n24424 vp_p.n24423 0.013
R18689 vp_p.n24438 vp_p.n24437 0.013
R18690 vp_p.n24452 vp_p.n24451 0.013
R18691 vp_p.n24456 vp_p.n24455 0.013
R18692 vp_p.n6179 vp_p.n6178 0.013
R18693 vp_p.n6193 vp_p.n6192 0.013
R18694 vp_p.n6207 vp_p.n6206 0.013
R18695 vp_p.n6221 vp_p.n6220 0.013
R18696 vp_p.n6235 vp_p.n6234 0.013
R18697 vp_p.n6249 vp_p.n6248 0.013
R18698 vp_p.n6263 vp_p.n6262 0.013
R18699 vp_p.n6277 vp_p.n6276 0.013
R18700 vp_p.n6291 vp_p.n6290 0.013
R18701 vp_p.n6305 vp_p.n6304 0.013
R18702 vp_p.n6319 vp_p.n6318 0.013
R18703 vp_p.n6333 vp_p.n6332 0.013
R18704 vp_p.n6347 vp_p.n6346 0.013
R18705 vp_p.n6361 vp_p.n6360 0.013
R18706 vp_p.n6375 vp_p.n6374 0.013
R18707 vp_p.n6389 vp_p.n6388 0.013
R18708 vp_p.n6403 vp_p.n6402 0.013
R18709 vp_p.n6417 vp_p.n6416 0.013
R18710 vp_p.n6431 vp_p.n6430 0.013
R18711 vp_p.n6445 vp_p.n6444 0.013
R18712 vp_p.n6459 vp_p.n6458 0.013
R18713 vp_p.n6473 vp_p.n6472 0.013
R18714 vp_p.n6487 vp_p.n6486 0.013
R18715 vp_p.n6501 vp_p.n6500 0.013
R18716 vp_p.n6515 vp_p.n6514 0.013
R18717 vp_p.n6529 vp_p.n6528 0.013
R18718 vp_p.n6543 vp_p.n6542 0.013
R18719 vp_p.n6557 vp_p.n6556 0.013
R18720 vp_p.n6571 vp_p.n6570 0.013
R18721 vp_p.n6585 vp_p.n6584 0.013
R18722 vp_p.n6599 vp_p.n6598 0.013
R18723 vp_p.n6613 vp_p.n6612 0.013
R18724 vp_p.n6627 vp_p.n6626 0.013
R18725 vp_p.n6641 vp_p.n6640 0.013
R18726 vp_p.n6655 vp_p.n6654 0.013
R18727 vp_p.n6669 vp_p.n6668 0.013
R18728 vp_p.n6683 vp_p.n6682 0.013
R18729 vp_p.n6697 vp_p.n6696 0.013
R18730 vp_p.n6711 vp_p.n6710 0.013
R18731 vp_p.n6725 vp_p.n6724 0.013
R18732 vp_p.n6739 vp_p.n6738 0.013
R18733 vp_p.n6753 vp_p.n6752 0.013
R18734 vp_p.n6767 vp_p.n6766 0.013
R18735 vp_p.n6781 vp_p.n6780 0.013
R18736 vp_p.n6795 vp_p.n6794 0.013
R18737 vp_p.n6809 vp_p.n6808 0.013
R18738 vp_p.n6823 vp_p.n6822 0.013
R18739 vp_p.n6837 vp_p.n6836 0.013
R18740 vp_p.n6851 vp_p.n6850 0.013
R18741 vp_p.n6865 vp_p.n6864 0.013
R18742 vp_p.n6879 vp_p.n6878 0.013
R18743 vp_p.n6893 vp_p.n6892 0.013
R18744 vp_p.n6907 vp_p.n6906 0.013
R18745 vp_p.n6921 vp_p.n6920 0.013
R18746 vp_p.n6935 vp_p.n6934 0.013
R18747 vp_p.n6949 vp_p.n6948 0.013
R18748 vp_p.n6963 vp_p.n6962 0.013
R18749 vp_p.n6977 vp_p.n6976 0.013
R18750 vp_p.n6991 vp_p.n6990 0.013
R18751 vp_p.n7005 vp_p.n7004 0.013
R18752 vp_p.n7019 vp_p.n7018 0.013
R18753 vp_p.n7033 vp_p.n7032 0.013
R18754 vp_p.n7047 vp_p.n7046 0.013
R18755 vp_p.n7061 vp_p.n7060 0.013
R18756 vp_p.n7075 vp_p.n7074 0.013
R18757 vp_p.n7089 vp_p.n7088 0.013
R18758 vp_p.n7103 vp_p.n7102 0.013
R18759 vp_p.n7117 vp_p.n7116 0.013
R18760 vp_p.n7131 vp_p.n7130 0.013
R18761 vp_p.n7145 vp_p.n7144 0.013
R18762 vp_p.n7159 vp_p.n7158 0.013
R18763 vp_p.n7173 vp_p.n7172 0.013
R18764 vp_p.n7187 vp_p.n7186 0.013
R18765 vp_p.n24880 vp_p.n24879 0.013
R18766 vp_p.n24894 vp_p.n24893 0.013
R18767 vp_p.n24908 vp_p.n24907 0.013
R18768 vp_p.n24922 vp_p.n24921 0.013
R18769 vp_p.n24936 vp_p.n24935 0.013
R18770 vp_p.n24950 vp_p.n24949 0.013
R18771 vp_p.n24964 vp_p.n24963 0.013
R18772 vp_p.n24978 vp_p.n24977 0.013
R18773 vp_p.n24992 vp_p.n24991 0.013
R18774 vp_p.n25006 vp_p.n25005 0.013
R18775 vp_p.n25020 vp_p.n25019 0.013
R18776 vp_p.n25034 vp_p.n25033 0.013
R18777 vp_p.n25048 vp_p.n25047 0.013
R18778 vp_p.n25062 vp_p.n25061 0.013
R18779 vp_p.n25076 vp_p.n25075 0.013
R18780 vp_p.n25090 vp_p.n25089 0.013
R18781 vp_p.n25104 vp_p.n25103 0.013
R18782 vp_p.n25118 vp_p.n25117 0.013
R18783 vp_p.n25132 vp_p.n25131 0.013
R18784 vp_p.n25146 vp_p.n25145 0.013
R18785 vp_p.n25160 vp_p.n25159 0.013
R18786 vp_p.n25174 vp_p.n25173 0.013
R18787 vp_p.n25188 vp_p.n25187 0.013
R18788 vp_p.n25202 vp_p.n25201 0.013
R18789 vp_p.n25216 vp_p.n25215 0.013
R18790 vp_p.n25230 vp_p.n25229 0.013
R18791 vp_p.n25244 vp_p.n25243 0.013
R18792 vp_p.n25258 vp_p.n25257 0.013
R18793 vp_p.n25272 vp_p.n25271 0.013
R18794 vp_p.n25286 vp_p.n25285 0.013
R18795 vp_p.n25300 vp_p.n25299 0.013
R18796 vp_p.n25314 vp_p.n25313 0.013
R18797 vp_p.n25328 vp_p.n25327 0.013
R18798 vp_p.n25342 vp_p.n25341 0.013
R18799 vp_p.n25356 vp_p.n25355 0.013
R18800 vp_p.n25370 vp_p.n25369 0.013
R18801 vp_p.n25384 vp_p.n25383 0.013
R18802 vp_p.n25398 vp_p.n25397 0.013
R18803 vp_p.n25412 vp_p.n25411 0.013
R18804 vp_p.n25426 vp_p.n25425 0.013
R18805 vp_p.n25440 vp_p.n25439 0.013
R18806 vp_p.n25454 vp_p.n25453 0.013
R18807 vp_p.n25468 vp_p.n25467 0.013
R18808 vp_p.n25482 vp_p.n25481 0.013
R18809 vp_p.n25496 vp_p.n25495 0.013
R18810 vp_p.n25510 vp_p.n25509 0.013
R18811 vp_p.n25524 vp_p.n25523 0.013
R18812 vp_p.n25538 vp_p.n25537 0.013
R18813 vp_p.n25552 vp_p.n25551 0.013
R18814 vp_p.n25566 vp_p.n25565 0.013
R18815 vp_p.n25580 vp_p.n25579 0.013
R18816 vp_p.n25594 vp_p.n25593 0.013
R18817 vp_p.n25608 vp_p.n25607 0.013
R18818 vp_p.n25622 vp_p.n25621 0.013
R18819 vp_p.n25636 vp_p.n25635 0.013
R18820 vp_p.n25650 vp_p.n25649 0.013
R18821 vp_p.n25664 vp_p.n25663 0.013
R18822 vp_p.n25678 vp_p.n25677 0.013
R18823 vp_p.n25692 vp_p.n25691 0.013
R18824 vp_p.n25706 vp_p.n25705 0.013
R18825 vp_p.n25720 vp_p.n25719 0.013
R18826 vp_p.n25734 vp_p.n25733 0.013
R18827 vp_p.n25748 vp_p.n25747 0.013
R18828 vp_p.n25762 vp_p.n25761 0.013
R18829 vp_p.n25776 vp_p.n25775 0.013
R18830 vp_p.n25790 vp_p.n25789 0.013
R18831 vp_p.n25804 vp_p.n25803 0.013
R18832 vp_p.n25818 vp_p.n25817 0.013
R18833 vp_p.n25832 vp_p.n25831 0.013
R18834 vp_p.n25846 vp_p.n25845 0.013
R18835 vp_p.n25860 vp_p.n25859 0.013
R18836 vp_p.n25874 vp_p.n25873 0.013
R18837 vp_p.n25888 vp_p.n25887 0.013
R18838 vp_p.n25892 vp_p.n25891 0.013
R18839 vp_p.n7601 vp_p.n7600 0.013
R18840 vp_p.n7615 vp_p.n7614 0.013
R18841 vp_p.n7629 vp_p.n7628 0.013
R18842 vp_p.n7643 vp_p.n7642 0.013
R18843 vp_p.n7657 vp_p.n7656 0.013
R18844 vp_p.n7671 vp_p.n7670 0.013
R18845 vp_p.n7685 vp_p.n7684 0.013
R18846 vp_p.n7699 vp_p.n7698 0.013
R18847 vp_p.n7713 vp_p.n7712 0.013
R18848 vp_p.n7727 vp_p.n7726 0.013
R18849 vp_p.n7741 vp_p.n7740 0.013
R18850 vp_p.n7755 vp_p.n7754 0.013
R18851 vp_p.n7769 vp_p.n7768 0.013
R18852 vp_p.n7783 vp_p.n7782 0.013
R18853 vp_p.n7797 vp_p.n7796 0.013
R18854 vp_p.n7811 vp_p.n7810 0.013
R18855 vp_p.n7825 vp_p.n7824 0.013
R18856 vp_p.n7839 vp_p.n7838 0.013
R18857 vp_p.n7853 vp_p.n7852 0.013
R18858 vp_p.n7867 vp_p.n7866 0.013
R18859 vp_p.n7881 vp_p.n7880 0.013
R18860 vp_p.n7895 vp_p.n7894 0.013
R18861 vp_p.n7909 vp_p.n7908 0.013
R18862 vp_p.n7923 vp_p.n7922 0.013
R18863 vp_p.n7937 vp_p.n7936 0.013
R18864 vp_p.n7951 vp_p.n7950 0.013
R18865 vp_p.n7965 vp_p.n7964 0.013
R18866 vp_p.n7979 vp_p.n7978 0.013
R18867 vp_p.n7993 vp_p.n7992 0.013
R18868 vp_p.n8007 vp_p.n8006 0.013
R18869 vp_p.n8021 vp_p.n8020 0.013
R18870 vp_p.n8035 vp_p.n8034 0.013
R18871 vp_p.n8049 vp_p.n8048 0.013
R18872 vp_p.n8063 vp_p.n8062 0.013
R18873 vp_p.n8077 vp_p.n8076 0.013
R18874 vp_p.n8091 vp_p.n8090 0.013
R18875 vp_p.n8105 vp_p.n8104 0.013
R18876 vp_p.n8119 vp_p.n8118 0.013
R18877 vp_p.n8133 vp_p.n8132 0.013
R18878 vp_p.n8147 vp_p.n8146 0.013
R18879 vp_p.n8161 vp_p.n8160 0.013
R18880 vp_p.n8175 vp_p.n8174 0.013
R18881 vp_p.n8189 vp_p.n8188 0.013
R18882 vp_p.n8203 vp_p.n8202 0.013
R18883 vp_p.n8217 vp_p.n8216 0.013
R18884 vp_p.n8231 vp_p.n8230 0.013
R18885 vp_p.n8245 vp_p.n8244 0.013
R18886 vp_p.n8259 vp_p.n8258 0.013
R18887 vp_p.n8273 vp_p.n8272 0.013
R18888 vp_p.n8287 vp_p.n8286 0.013
R18889 vp_p.n8301 vp_p.n8300 0.013
R18890 vp_p.n8315 vp_p.n8314 0.013
R18891 vp_p.n8329 vp_p.n8328 0.013
R18892 vp_p.n8343 vp_p.n8342 0.013
R18893 vp_p.n8357 vp_p.n8356 0.013
R18894 vp_p.n8371 vp_p.n8370 0.013
R18895 vp_p.n8385 vp_p.n8384 0.013
R18896 vp_p.n8399 vp_p.n8398 0.013
R18897 vp_p.n8413 vp_p.n8412 0.013
R18898 vp_p.n8427 vp_p.n8426 0.013
R18899 vp_p.n8441 vp_p.n8440 0.013
R18900 vp_p.n8455 vp_p.n8454 0.013
R18901 vp_p.n8469 vp_p.n8468 0.013
R18902 vp_p.n8483 vp_p.n8482 0.013
R18903 vp_p.n8497 vp_p.n8496 0.013
R18904 vp_p.n8511 vp_p.n8510 0.013
R18905 vp_p.n8525 vp_p.n8524 0.013
R18906 vp_p.n8539 vp_p.n8538 0.013
R18907 vp_p.n8553 vp_p.n8552 0.013
R18908 vp_p.n8567 vp_p.n8566 0.013
R18909 vp_p.n8581 vp_p.n8580 0.013
R18910 vp_p.n8595 vp_p.n8594 0.013
R18911 vp_p.n8609 vp_p.n8608 0.013
R18912 vp_p.n26291 vp_p.n26290 0.013
R18913 vp_p.n26305 vp_p.n26304 0.013
R18914 vp_p.n26319 vp_p.n26318 0.013
R18915 vp_p.n26333 vp_p.n26332 0.013
R18916 vp_p.n26347 vp_p.n26346 0.013
R18917 vp_p.n26361 vp_p.n26360 0.013
R18918 vp_p.n26375 vp_p.n26374 0.013
R18919 vp_p.n26389 vp_p.n26388 0.013
R18920 vp_p.n26403 vp_p.n26402 0.013
R18921 vp_p.n26417 vp_p.n26416 0.013
R18922 vp_p.n26431 vp_p.n26430 0.013
R18923 vp_p.n26445 vp_p.n26444 0.013
R18924 vp_p.n26459 vp_p.n26458 0.013
R18925 vp_p.n26473 vp_p.n26472 0.013
R18926 vp_p.n26487 vp_p.n26486 0.013
R18927 vp_p.n26501 vp_p.n26500 0.013
R18928 vp_p.n26515 vp_p.n26514 0.013
R18929 vp_p.n26529 vp_p.n26528 0.013
R18930 vp_p.n26543 vp_p.n26542 0.013
R18931 vp_p.n26557 vp_p.n26556 0.013
R18932 vp_p.n26571 vp_p.n26570 0.013
R18933 vp_p.n26585 vp_p.n26584 0.013
R18934 vp_p.n26599 vp_p.n26598 0.013
R18935 vp_p.n26613 vp_p.n26612 0.013
R18936 vp_p.n26627 vp_p.n26626 0.013
R18937 vp_p.n26641 vp_p.n26640 0.013
R18938 vp_p.n26655 vp_p.n26654 0.013
R18939 vp_p.n26669 vp_p.n26668 0.013
R18940 vp_p.n26683 vp_p.n26682 0.013
R18941 vp_p.n26697 vp_p.n26696 0.013
R18942 vp_p.n26711 vp_p.n26710 0.013
R18943 vp_p.n26725 vp_p.n26724 0.013
R18944 vp_p.n26739 vp_p.n26738 0.013
R18945 vp_p.n26753 vp_p.n26752 0.013
R18946 vp_p.n26767 vp_p.n26766 0.013
R18947 vp_p.n26781 vp_p.n26780 0.013
R18948 vp_p.n26795 vp_p.n26794 0.013
R18949 vp_p.n26809 vp_p.n26808 0.013
R18950 vp_p.n26823 vp_p.n26822 0.013
R18951 vp_p.n26837 vp_p.n26836 0.013
R18952 vp_p.n26851 vp_p.n26850 0.013
R18953 vp_p.n26865 vp_p.n26864 0.013
R18954 vp_p.n26879 vp_p.n26878 0.013
R18955 vp_p.n26893 vp_p.n26892 0.013
R18956 vp_p.n26907 vp_p.n26906 0.013
R18957 vp_p.n26921 vp_p.n26920 0.013
R18958 vp_p.n26935 vp_p.n26934 0.013
R18959 vp_p.n26949 vp_p.n26948 0.013
R18960 vp_p.n26963 vp_p.n26962 0.013
R18961 vp_p.n26977 vp_p.n26976 0.013
R18962 vp_p.n26991 vp_p.n26990 0.013
R18963 vp_p.n27005 vp_p.n27004 0.013
R18964 vp_p.n27019 vp_p.n27018 0.013
R18965 vp_p.n27033 vp_p.n27032 0.013
R18966 vp_p.n27047 vp_p.n27046 0.013
R18967 vp_p.n27061 vp_p.n27060 0.013
R18968 vp_p.n27075 vp_p.n27074 0.013
R18969 vp_p.n27089 vp_p.n27088 0.013
R18970 vp_p.n27103 vp_p.n27102 0.013
R18971 vp_p.n27117 vp_p.n27116 0.013
R18972 vp_p.n27131 vp_p.n27130 0.013
R18973 vp_p.n27145 vp_p.n27144 0.013
R18974 vp_p.n27159 vp_p.n27158 0.013
R18975 vp_p.n27173 vp_p.n27172 0.013
R18976 vp_p.n27187 vp_p.n27186 0.013
R18977 vp_p.n27201 vp_p.n27200 0.013
R18978 vp_p.n27215 vp_p.n27214 0.013
R18979 vp_p.n27229 vp_p.n27228 0.013
R18980 vp_p.n27243 vp_p.n27242 0.013
R18981 vp_p.n27257 vp_p.n27256 0.013
R18982 vp_p.n27271 vp_p.n27270 0.013
R18983 vp_p.n27285 vp_p.n27284 0.013
R18984 vp_p.n27299 vp_p.n27298 0.013
R18985 vp_p.n27313 vp_p.n27312 0.013
R18986 vp_p.n27327 vp_p.n27326 0.013
R18987 vp_p.n12098 vp_p.n12097 0.009
R18988 vp_p.n12112 vp_p.n12111 0.009
R18989 vp_p.n12126 vp_p.n12125 0.009
R18990 vp_p.n12140 vp_p.n12139 0.009
R18991 vp_p.n12154 vp_p.n12153 0.009
R18992 vp_p.n12168 vp_p.n12167 0.009
R18993 vp_p.n12182 vp_p.n12181 0.009
R18994 vp_p.n12196 vp_p.n12195 0.009
R18995 vp_p.n12210 vp_p.n12209 0.009
R18996 vp_p.n12224 vp_p.n12223 0.009
R18997 vp_p.n12238 vp_p.n12237 0.009
R18998 vp_p.n12252 vp_p.n12251 0.009
R18999 vp_p.n12266 vp_p.n12265 0.009
R19000 vp_p.n12280 vp_p.n12279 0.009
R19001 vp_p.n12294 vp_p.n12293 0.009
R19002 vp_p.n12308 vp_p.n12307 0.009
R19003 vp_p.n12322 vp_p.n12321 0.009
R19004 vp_p.n12336 vp_p.n12335 0.009
R19005 vp_p.n12350 vp_p.n12349 0.009
R19006 vp_p.n12364 vp_p.n12363 0.009
R19007 vp_p.n12378 vp_p.n12377 0.009
R19008 vp_p.n12392 vp_p.n12391 0.009
R19009 vp_p.n12406 vp_p.n12405 0.009
R19010 vp_p.n12420 vp_p.n12419 0.009
R19011 vp_p.n12434 vp_p.n12433 0.009
R19012 vp_p.n12448 vp_p.n12447 0.009
R19013 vp_p.n12462 vp_p.n12461 0.009
R19014 vp_p.n12476 vp_p.n12475 0.009
R19015 vp_p.n12490 vp_p.n12489 0.009
R19016 vp_p.n12504 vp_p.n12503 0.009
R19017 vp_p.n12518 vp_p.n12517 0.009
R19018 vp_p.n12532 vp_p.n12531 0.009
R19019 vp_p.n12546 vp_p.n12545 0.009
R19020 vp_p.n12560 vp_p.n12559 0.009
R19021 vp_p.n12574 vp_p.n12573 0.009
R19022 vp_p.n12588 vp_p.n12587 0.009
R19023 vp_p.n12602 vp_p.n12601 0.009
R19024 vp_p.n12616 vp_p.n12615 0.009
R19025 vp_p.n12630 vp_p.n12629 0.009
R19026 vp_p.n12644 vp_p.n12643 0.009
R19027 vp_p.n12658 vp_p.n12657 0.009
R19028 vp_p.n12672 vp_p.n12671 0.009
R19029 vp_p.n12686 vp_p.n12685 0.009
R19030 vp_p.n12700 vp_p.n12699 0.009
R19031 vp_p.n12714 vp_p.n12713 0.009
R19032 vp_p.n12728 vp_p.n12727 0.009
R19033 vp_p.n12742 vp_p.n12741 0.009
R19034 vp_p.n12756 vp_p.n12755 0.009
R19035 vp_p.n12770 vp_p.n12769 0.009
R19036 vp_p.n12784 vp_p.n12783 0.009
R19037 vp_p.n12798 vp_p.n12797 0.009
R19038 vp_p.n12812 vp_p.n12811 0.009
R19039 vp_p.n12826 vp_p.n12825 0.009
R19040 vp_p.n12840 vp_p.n12839 0.009
R19041 vp_p.n12854 vp_p.n12853 0.009
R19042 vp_p.n12868 vp_p.n12867 0.009
R19043 vp_p.n12882 vp_p.n12881 0.009
R19044 vp_p.n12896 vp_p.n12895 0.009
R19045 vp_p.n12910 vp_p.n12909 0.009
R19046 vp_p.n12924 vp_p.n12923 0.009
R19047 vp_p.n12938 vp_p.n12937 0.009
R19048 vp_p.n12952 vp_p.n12951 0.009
R19049 vp_p.n12966 vp_p.n12965 0.009
R19050 vp_p.n12980 vp_p.n12979 0.009
R19051 vp_p.n12994 vp_p.n12993 0.009
R19052 vp_p.n13008 vp_p.n13007 0.009
R19053 vp_p.n14901 vp_p.n14900 0.009
R19054 vp_p.n14915 vp_p.n14914 0.009
R19055 vp_p.n14929 vp_p.n14928 0.009
R19056 vp_p.n14943 vp_p.n14942 0.009
R19057 vp_p.n14957 vp_p.n14956 0.009
R19058 vp_p.n14971 vp_p.n14970 0.009
R19059 vp_p.n14985 vp_p.n14984 0.009
R19060 vp_p.n14999 vp_p.n14998 0.009
R19061 vp_p.n15013 vp_p.n15012 0.009
R19062 vp_p.n15027 vp_p.n15026 0.009
R19063 vp_p.n15041 vp_p.n15040 0.009
R19064 vp_p.n15055 vp_p.n15054 0.009
R19065 vp_p.n15069 vp_p.n15068 0.009
R19066 vp_p.n15083 vp_p.n15082 0.009
R19067 vp_p.n15097 vp_p.n15096 0.009
R19068 vp_p.n15111 vp_p.n15110 0.009
R19069 vp_p.n15125 vp_p.n15124 0.009
R19070 vp_p.n15139 vp_p.n15138 0.009
R19071 vp_p.n15153 vp_p.n15152 0.009
R19072 vp_p.n15167 vp_p.n15166 0.009
R19073 vp_p.n15181 vp_p.n15180 0.009
R19074 vp_p.n15195 vp_p.n15194 0.009
R19075 vp_p.n15209 vp_p.n15208 0.009
R19076 vp_p.n15223 vp_p.n15222 0.009
R19077 vp_p.n15237 vp_p.n15236 0.009
R19078 vp_p.n15251 vp_p.n15250 0.009
R19079 vp_p.n15265 vp_p.n15264 0.009
R19080 vp_p.n15279 vp_p.n15278 0.009
R19081 vp_p.n15293 vp_p.n15292 0.009
R19082 vp_p.n15307 vp_p.n15306 0.009
R19083 vp_p.n15321 vp_p.n15320 0.009
R19084 vp_p.n15335 vp_p.n15334 0.009
R19085 vp_p.n15349 vp_p.n15348 0.009
R19086 vp_p.n15363 vp_p.n15362 0.009
R19087 vp_p.n15377 vp_p.n15376 0.009
R19088 vp_p.n15391 vp_p.n15390 0.009
R19089 vp_p.n15405 vp_p.n15404 0.009
R19090 vp_p.n15419 vp_p.n15418 0.009
R19091 vp_p.n15433 vp_p.n15432 0.009
R19092 vp_p.n15447 vp_p.n15446 0.009
R19093 vp_p.n15461 vp_p.n15460 0.009
R19094 vp_p.n15475 vp_p.n15474 0.009
R19095 vp_p.n15489 vp_p.n15488 0.009
R19096 vp_p.n15503 vp_p.n15502 0.009
R19097 vp_p.n15517 vp_p.n15516 0.009
R19098 vp_p.n15531 vp_p.n15530 0.009
R19099 vp_p.n15545 vp_p.n15544 0.009
R19100 vp_p.n15559 vp_p.n15558 0.009
R19101 vp_p.n15573 vp_p.n15572 0.009
R19102 vp_p.n15587 vp_p.n15586 0.009
R19103 vp_p.n15601 vp_p.n15600 0.009
R19104 vp_p.n15615 vp_p.n15614 0.009
R19105 vp_p.n15629 vp_p.n15628 0.009
R19106 vp_p.n15643 vp_p.n15642 0.009
R19107 vp_p.n15657 vp_p.n15656 0.009
R19108 vp_p.n15671 vp_p.n15670 0.009
R19109 vp_p.n15685 vp_p.n15684 0.009
R19110 vp_p.n15699 vp_p.n15698 0.009
R19111 vp_p.n15713 vp_p.n15712 0.009
R19112 vp_p.n15727 vp_p.n15726 0.009
R19113 vp_p.n15741 vp_p.n15740 0.009
R19114 vp_p.n15755 vp_p.n15754 0.009
R19115 vp_p.n15769 vp_p.n15768 0.009
R19116 vp_p.n15783 vp_p.n15782 0.009
R19117 vp_p.n15797 vp_p.n15796 0.009
R19118 vp_p.n15811 vp_p.n15810 0.009
R19119 vp_p.n10660 vp_p.n10659 0.009
R19120 vp_p.n10674 vp_p.n10673 0.009
R19121 vp_p.n10688 vp_p.n10687 0.009
R19122 vp_p.n10702 vp_p.n10701 0.009
R19123 vp_p.n10716 vp_p.n10715 0.009
R19124 vp_p.n10730 vp_p.n10729 0.009
R19125 vp_p.n10744 vp_p.n10743 0.009
R19126 vp_p.n10758 vp_p.n10757 0.009
R19127 vp_p.n10772 vp_p.n10771 0.009
R19128 vp_p.n10786 vp_p.n10785 0.009
R19129 vp_p.n10800 vp_p.n10799 0.009
R19130 vp_p.n10814 vp_p.n10813 0.009
R19131 vp_p.n10828 vp_p.n10827 0.009
R19132 vp_p.n10842 vp_p.n10841 0.009
R19133 vp_p.n10856 vp_p.n10855 0.009
R19134 vp_p.n10870 vp_p.n10869 0.009
R19135 vp_p.n10884 vp_p.n10883 0.009
R19136 vp_p.n10898 vp_p.n10897 0.009
R19137 vp_p.n10912 vp_p.n10911 0.009
R19138 vp_p.n10926 vp_p.n10925 0.009
R19139 vp_p.n10940 vp_p.n10939 0.009
R19140 vp_p.n10954 vp_p.n10953 0.009
R19141 vp_p.n10968 vp_p.n10967 0.009
R19142 vp_p.n10982 vp_p.n10981 0.009
R19143 vp_p.n10996 vp_p.n10995 0.009
R19144 vp_p.n11010 vp_p.n11009 0.009
R19145 vp_p.n11024 vp_p.n11023 0.009
R19146 vp_p.n11038 vp_p.n11037 0.009
R19147 vp_p.n11052 vp_p.n11051 0.009
R19148 vp_p.n11066 vp_p.n11065 0.009
R19149 vp_p.n11080 vp_p.n11079 0.009
R19150 vp_p.n11094 vp_p.n11093 0.009
R19151 vp_p.n11108 vp_p.n11107 0.009
R19152 vp_p.n11122 vp_p.n11121 0.009
R19153 vp_p.n11136 vp_p.n11135 0.009
R19154 vp_p.n11150 vp_p.n11149 0.009
R19155 vp_p.n11164 vp_p.n11163 0.009
R19156 vp_p.n11178 vp_p.n11177 0.009
R19157 vp_p.n11192 vp_p.n11191 0.009
R19158 vp_p.n11206 vp_p.n11205 0.009
R19159 vp_p.n11220 vp_p.n11219 0.009
R19160 vp_p.n11234 vp_p.n11233 0.009
R19161 vp_p.n11248 vp_p.n11247 0.009
R19162 vp_p.n11262 vp_p.n11261 0.009
R19163 vp_p.n11276 vp_p.n11275 0.009
R19164 vp_p.n11290 vp_p.n11289 0.009
R19165 vp_p.n11304 vp_p.n11303 0.009
R19166 vp_p.n11318 vp_p.n11317 0.009
R19167 vp_p.n11332 vp_p.n11331 0.009
R19168 vp_p.n11346 vp_p.n11345 0.009
R19169 vp_p.n11360 vp_p.n11359 0.009
R19170 vp_p.n11374 vp_p.n11373 0.009
R19171 vp_p.n11388 vp_p.n11387 0.009
R19172 vp_p.n11402 vp_p.n11401 0.009
R19173 vp_p.n11416 vp_p.n11415 0.009
R19174 vp_p.n11430 vp_p.n11429 0.009
R19175 vp_p.n11444 vp_p.n11443 0.009
R19176 vp_p.n11458 vp_p.n11457 0.009
R19177 vp_p.n11472 vp_p.n11471 0.009
R19178 vp_p.n11486 vp_p.n11485 0.009
R19179 vp_p.n11500 vp_p.n11499 0.009
R19180 vp_p.n11514 vp_p.n11513 0.009
R19181 vp_p.n11528 vp_p.n11527 0.009
R19182 vp_p.n11542 vp_p.n11541 0.009
R19183 vp_p.n11556 vp_p.n11555 0.009
R19184 vp_p.n11570 vp_p.n11569 0.009
R19185 vp_p.n11584 vp_p.n11583 0.009
R19186 vp_p.n16329 vp_p.n16328 0.009
R19187 vp_p.n16343 vp_p.n16342 0.009
R19188 vp_p.n16357 vp_p.n16356 0.009
R19189 vp_p.n16371 vp_p.n16370 0.009
R19190 vp_p.n16385 vp_p.n16384 0.009
R19191 vp_p.n16399 vp_p.n16398 0.009
R19192 vp_p.n16413 vp_p.n16412 0.009
R19193 vp_p.n16427 vp_p.n16426 0.009
R19194 vp_p.n16441 vp_p.n16440 0.009
R19195 vp_p.n16455 vp_p.n16454 0.009
R19196 vp_p.n16469 vp_p.n16468 0.009
R19197 vp_p.n16483 vp_p.n16482 0.009
R19198 vp_p.n16497 vp_p.n16496 0.009
R19199 vp_p.n16511 vp_p.n16510 0.009
R19200 vp_p.n16525 vp_p.n16524 0.009
R19201 vp_p.n16539 vp_p.n16538 0.009
R19202 vp_p.n16553 vp_p.n16552 0.009
R19203 vp_p.n16567 vp_p.n16566 0.009
R19204 vp_p.n16581 vp_p.n16580 0.009
R19205 vp_p.n16595 vp_p.n16594 0.009
R19206 vp_p.n16609 vp_p.n16608 0.009
R19207 vp_p.n16623 vp_p.n16622 0.009
R19208 vp_p.n16637 vp_p.n16636 0.009
R19209 vp_p.n16651 vp_p.n16650 0.009
R19210 vp_p.n16665 vp_p.n16664 0.009
R19211 vp_p.n16679 vp_p.n16678 0.009
R19212 vp_p.n16693 vp_p.n16692 0.009
R19213 vp_p.n16707 vp_p.n16706 0.009
R19214 vp_p.n16721 vp_p.n16720 0.009
R19215 vp_p.n16735 vp_p.n16734 0.009
R19216 vp_p.n16749 vp_p.n16748 0.009
R19217 vp_p.n16763 vp_p.n16762 0.009
R19218 vp_p.n16777 vp_p.n16776 0.009
R19219 vp_p.n16791 vp_p.n16790 0.009
R19220 vp_p.n16805 vp_p.n16804 0.009
R19221 vp_p.n16819 vp_p.n16818 0.009
R19222 vp_p.n16833 vp_p.n16832 0.009
R19223 vp_p.n16847 vp_p.n16846 0.009
R19224 vp_p.n16861 vp_p.n16860 0.009
R19225 vp_p.n16875 vp_p.n16874 0.009
R19226 vp_p.n16889 vp_p.n16888 0.009
R19227 vp_p.n16903 vp_p.n16902 0.009
R19228 vp_p.n16917 vp_p.n16916 0.009
R19229 vp_p.n16931 vp_p.n16930 0.009
R19230 vp_p.n16945 vp_p.n16944 0.009
R19231 vp_p.n16959 vp_p.n16958 0.009
R19232 vp_p.n16973 vp_p.n16972 0.009
R19233 vp_p.n16987 vp_p.n16986 0.009
R19234 vp_p.n17001 vp_p.n17000 0.009
R19235 vp_p.n17015 vp_p.n17014 0.009
R19236 vp_p.n17029 vp_p.n17028 0.009
R19237 vp_p.n17043 vp_p.n17042 0.009
R19238 vp_p.n17057 vp_p.n17056 0.009
R19239 vp_p.n17071 vp_p.n17070 0.009
R19240 vp_p.n17085 vp_p.n17084 0.009
R19241 vp_p.n17099 vp_p.n17098 0.009
R19242 vp_p.n17113 vp_p.n17112 0.009
R19243 vp_p.n17127 vp_p.n17126 0.009
R19244 vp_p.n17141 vp_p.n17140 0.009
R19245 vp_p.n17155 vp_p.n17154 0.009
R19246 vp_p.n17169 vp_p.n17168 0.009
R19247 vp_p.n17183 vp_p.n17182 0.009
R19248 vp_p.n17197 vp_p.n17196 0.009
R19249 vp_p.n17211 vp_p.n17210 0.009
R19250 vp_p.n17225 vp_p.n17224 0.009
R19251 vp_p.n17239 vp_p.n17238 0.009
R19252 vp_p.n17253 vp_p.n17252 0.009
R19253 vp_p.n9223 vp_p.n9222 0.009
R19254 vp_p.n9237 vp_p.n9236 0.009
R19255 vp_p.n9251 vp_p.n9250 0.009
R19256 vp_p.n9265 vp_p.n9264 0.009
R19257 vp_p.n9279 vp_p.n9278 0.009
R19258 vp_p.n9293 vp_p.n9292 0.009
R19259 vp_p.n9307 vp_p.n9306 0.009
R19260 vp_p.n9321 vp_p.n9320 0.009
R19261 vp_p.n9335 vp_p.n9334 0.009
R19262 vp_p.n9349 vp_p.n9348 0.009
R19263 vp_p.n9363 vp_p.n9362 0.009
R19264 vp_p.n9377 vp_p.n9376 0.009
R19265 vp_p.n9391 vp_p.n9390 0.009
R19266 vp_p.n9405 vp_p.n9404 0.009
R19267 vp_p.n9419 vp_p.n9418 0.009
R19268 vp_p.n9433 vp_p.n9432 0.009
R19269 vp_p.n9447 vp_p.n9446 0.009
R19270 vp_p.n9461 vp_p.n9460 0.009
R19271 vp_p.n9475 vp_p.n9474 0.009
R19272 vp_p.n9489 vp_p.n9488 0.009
R19273 vp_p.n9503 vp_p.n9502 0.009
R19274 vp_p.n9517 vp_p.n9516 0.009
R19275 vp_p.n9531 vp_p.n9530 0.009
R19276 vp_p.n9545 vp_p.n9544 0.009
R19277 vp_p.n9559 vp_p.n9558 0.009
R19278 vp_p.n9573 vp_p.n9572 0.009
R19279 vp_p.n9587 vp_p.n9586 0.009
R19280 vp_p.n9601 vp_p.n9600 0.009
R19281 vp_p.n9615 vp_p.n9614 0.009
R19282 vp_p.n9629 vp_p.n9628 0.009
R19283 vp_p.n9643 vp_p.n9642 0.009
R19284 vp_p.n9657 vp_p.n9656 0.009
R19285 vp_p.n9671 vp_p.n9670 0.009
R19286 vp_p.n9685 vp_p.n9684 0.009
R19287 vp_p.n9699 vp_p.n9698 0.009
R19288 vp_p.n9713 vp_p.n9712 0.009
R19289 vp_p.n9727 vp_p.n9726 0.009
R19290 vp_p.n9741 vp_p.n9740 0.009
R19291 vp_p.n9755 vp_p.n9754 0.009
R19292 vp_p.n9769 vp_p.n9768 0.009
R19293 vp_p.n9783 vp_p.n9782 0.009
R19294 vp_p.n9797 vp_p.n9796 0.009
R19295 vp_p.n9811 vp_p.n9810 0.009
R19296 vp_p.n9825 vp_p.n9824 0.009
R19297 vp_p.n9839 vp_p.n9838 0.009
R19298 vp_p.n9853 vp_p.n9852 0.009
R19299 vp_p.n9867 vp_p.n9866 0.009
R19300 vp_p.n9881 vp_p.n9880 0.009
R19301 vp_p.n9895 vp_p.n9894 0.009
R19302 vp_p.n9909 vp_p.n9908 0.009
R19303 vp_p.n9923 vp_p.n9922 0.009
R19304 vp_p.n9937 vp_p.n9936 0.009
R19305 vp_p.n9951 vp_p.n9950 0.009
R19306 vp_p.n9965 vp_p.n9964 0.009
R19307 vp_p.n9979 vp_p.n9978 0.009
R19308 vp_p.n9993 vp_p.n9992 0.009
R19309 vp_p.n10007 vp_p.n10006 0.009
R19310 vp_p.n10021 vp_p.n10020 0.009
R19311 vp_p.n10035 vp_p.n10034 0.009
R19312 vp_p.n10049 vp_p.n10048 0.009
R19313 vp_p.n10063 vp_p.n10062 0.009
R19314 vp_p.n10077 vp_p.n10076 0.009
R19315 vp_p.n10091 vp_p.n10090 0.009
R19316 vp_p.n10105 vp_p.n10104 0.009
R19317 vp_p.n10119 vp_p.n10118 0.009
R19318 vp_p.n10133 vp_p.n10132 0.009
R19319 vp_p.n10147 vp_p.n10146 0.009
R19320 vp_p.n10161 vp_p.n10160 0.009
R19321 vp_p.n17756 vp_p.n17755 0.009
R19322 vp_p.n17770 vp_p.n17769 0.009
R19323 vp_p.n17784 vp_p.n17783 0.009
R19324 vp_p.n17798 vp_p.n17797 0.009
R19325 vp_p.n17812 vp_p.n17811 0.009
R19326 vp_p.n17826 vp_p.n17825 0.009
R19327 vp_p.n17840 vp_p.n17839 0.009
R19328 vp_p.n17854 vp_p.n17853 0.009
R19329 vp_p.n17868 vp_p.n17867 0.009
R19330 vp_p.n17882 vp_p.n17881 0.009
R19331 vp_p.n17896 vp_p.n17895 0.009
R19332 vp_p.n17910 vp_p.n17909 0.009
R19333 vp_p.n17924 vp_p.n17923 0.009
R19334 vp_p.n17938 vp_p.n17937 0.009
R19335 vp_p.n17952 vp_p.n17951 0.009
R19336 vp_p.n17966 vp_p.n17965 0.009
R19337 vp_p.n17980 vp_p.n17979 0.009
R19338 vp_p.n17994 vp_p.n17993 0.009
R19339 vp_p.n18008 vp_p.n18007 0.009
R19340 vp_p.n18022 vp_p.n18021 0.009
R19341 vp_p.n18036 vp_p.n18035 0.009
R19342 vp_p.n18050 vp_p.n18049 0.009
R19343 vp_p.n18064 vp_p.n18063 0.009
R19344 vp_p.n18078 vp_p.n18077 0.009
R19345 vp_p.n18092 vp_p.n18091 0.009
R19346 vp_p.n18106 vp_p.n18105 0.009
R19347 vp_p.n18120 vp_p.n18119 0.009
R19348 vp_p.n18134 vp_p.n18133 0.009
R19349 vp_p.n18148 vp_p.n18147 0.009
R19350 vp_p.n18162 vp_p.n18161 0.009
R19351 vp_p.n18176 vp_p.n18175 0.009
R19352 vp_p.n18190 vp_p.n18189 0.009
R19353 vp_p.n18204 vp_p.n18203 0.009
R19354 vp_p.n18218 vp_p.n18217 0.009
R19355 vp_p.n18232 vp_p.n18231 0.009
R19356 vp_p.n18246 vp_p.n18245 0.009
R19357 vp_p.n18260 vp_p.n18259 0.009
R19358 vp_p.n18274 vp_p.n18273 0.009
R19359 vp_p.n18288 vp_p.n18287 0.009
R19360 vp_p.n18302 vp_p.n18301 0.009
R19361 vp_p.n18316 vp_p.n18315 0.009
R19362 vp_p.n18330 vp_p.n18329 0.009
R19363 vp_p.n18344 vp_p.n18343 0.009
R19364 vp_p.n18358 vp_p.n18357 0.009
R19365 vp_p.n18372 vp_p.n18371 0.009
R19366 vp_p.n18386 vp_p.n18385 0.009
R19367 vp_p.n18400 vp_p.n18399 0.009
R19368 vp_p.n18414 vp_p.n18413 0.009
R19369 vp_p.n18428 vp_p.n18427 0.009
R19370 vp_p.n18442 vp_p.n18441 0.009
R19371 vp_p.n18456 vp_p.n18455 0.009
R19372 vp_p.n18470 vp_p.n18469 0.009
R19373 vp_p.n18484 vp_p.n18483 0.009
R19374 vp_p.n18498 vp_p.n18497 0.009
R19375 vp_p.n18512 vp_p.n18511 0.009
R19376 vp_p.n18526 vp_p.n18525 0.009
R19377 vp_p.n18540 vp_p.n18539 0.009
R19378 vp_p.n18554 vp_p.n18553 0.009
R19379 vp_p.n18568 vp_p.n18567 0.009
R19380 vp_p.n18582 vp_p.n18581 0.009
R19381 vp_p.n18596 vp_p.n18595 0.009
R19382 vp_p.n18610 vp_p.n18609 0.009
R19383 vp_p.n18624 vp_p.n18623 0.009
R19384 vp_p.n18638 vp_p.n18637 0.009
R19385 vp_p.n18652 vp_p.n18651 0.009
R19386 vp_p.n18666 vp_p.n18665 0.009
R19387 vp_p.n18680 vp_p.n18679 0.009
R19388 vp_p.n18694 vp_p.n18693 0.009
R19389 vp_p.n477 vp_p.n476 0.009
R19390 vp_p.n491 vp_p.n490 0.009
R19391 vp_p.n505 vp_p.n504 0.009
R19392 vp_p.n519 vp_p.n518 0.009
R19393 vp_p.n533 vp_p.n532 0.009
R19394 vp_p.n547 vp_p.n546 0.009
R19395 vp_p.n561 vp_p.n560 0.009
R19396 vp_p.n575 vp_p.n574 0.009
R19397 vp_p.n589 vp_p.n588 0.009
R19398 vp_p.n603 vp_p.n602 0.009
R19399 vp_p.n617 vp_p.n616 0.009
R19400 vp_p.n631 vp_p.n630 0.009
R19401 vp_p.n645 vp_p.n644 0.009
R19402 vp_p.n659 vp_p.n658 0.009
R19403 vp_p.n673 vp_p.n672 0.009
R19404 vp_p.n687 vp_p.n686 0.009
R19405 vp_p.n701 vp_p.n700 0.009
R19406 vp_p.n715 vp_p.n714 0.009
R19407 vp_p.n729 vp_p.n728 0.009
R19408 vp_p.n743 vp_p.n742 0.009
R19409 vp_p.n757 vp_p.n756 0.009
R19410 vp_p.n771 vp_p.n770 0.009
R19411 vp_p.n785 vp_p.n784 0.009
R19412 vp_p.n799 vp_p.n798 0.009
R19413 vp_p.n813 vp_p.n812 0.009
R19414 vp_p.n827 vp_p.n826 0.009
R19415 vp_p.n841 vp_p.n840 0.009
R19416 vp_p.n855 vp_p.n854 0.009
R19417 vp_p.n869 vp_p.n868 0.009
R19418 vp_p.n883 vp_p.n882 0.009
R19419 vp_p.n897 vp_p.n896 0.009
R19420 vp_p.n911 vp_p.n910 0.009
R19421 vp_p.n925 vp_p.n924 0.009
R19422 vp_p.n939 vp_p.n938 0.009
R19423 vp_p.n953 vp_p.n952 0.009
R19424 vp_p.n967 vp_p.n966 0.009
R19425 vp_p.n981 vp_p.n980 0.009
R19426 vp_p.n995 vp_p.n994 0.009
R19427 vp_p.n1009 vp_p.n1008 0.009
R19428 vp_p.n1023 vp_p.n1022 0.009
R19429 vp_p.n1037 vp_p.n1036 0.009
R19430 vp_p.n1051 vp_p.n1050 0.009
R19431 vp_p.n1065 vp_p.n1064 0.009
R19432 vp_p.n1079 vp_p.n1078 0.009
R19433 vp_p.n1093 vp_p.n1092 0.009
R19434 vp_p.n1107 vp_p.n1106 0.009
R19435 vp_p.n1121 vp_p.n1120 0.009
R19436 vp_p.n1135 vp_p.n1134 0.009
R19437 vp_p.n1149 vp_p.n1148 0.009
R19438 vp_p.n1163 vp_p.n1162 0.009
R19439 vp_p.n1177 vp_p.n1176 0.009
R19440 vp_p.n1191 vp_p.n1190 0.009
R19441 vp_p.n1205 vp_p.n1204 0.009
R19442 vp_p.n1219 vp_p.n1218 0.009
R19443 vp_p.n1233 vp_p.n1232 0.009
R19444 vp_p.n1247 vp_p.n1246 0.009
R19445 vp_p.n1261 vp_p.n1260 0.009
R19446 vp_p.n1275 vp_p.n1274 0.009
R19447 vp_p.n1289 vp_p.n1288 0.009
R19448 vp_p.n1303 vp_p.n1302 0.009
R19449 vp_p.n1317 vp_p.n1316 0.009
R19450 vp_p.n1331 vp_p.n1330 0.009
R19451 vp_p.n1345 vp_p.n1344 0.009
R19452 vp_p.n1359 vp_p.n1358 0.009
R19453 vp_p.n1373 vp_p.n1372 0.009
R19454 vp_p.n1387 vp_p.n1386 0.009
R19455 vp_p.n1401 vp_p.n1400 0.009
R19456 vp_p.n1415 vp_p.n1414 0.009
R19457 vp_p.n1429 vp_p.n1428 0.009
R19458 vp_p.n19182 vp_p.n19181 0.009
R19459 vp_p.n19196 vp_p.n19195 0.009
R19460 vp_p.n19210 vp_p.n19209 0.009
R19461 vp_p.n19224 vp_p.n19223 0.009
R19462 vp_p.n19238 vp_p.n19237 0.009
R19463 vp_p.n19252 vp_p.n19251 0.009
R19464 vp_p.n19266 vp_p.n19265 0.009
R19465 vp_p.n19280 vp_p.n19279 0.009
R19466 vp_p.n19294 vp_p.n19293 0.009
R19467 vp_p.n19308 vp_p.n19307 0.009
R19468 vp_p.n19322 vp_p.n19321 0.009
R19469 vp_p.n19336 vp_p.n19335 0.009
R19470 vp_p.n19350 vp_p.n19349 0.009
R19471 vp_p.n19364 vp_p.n19363 0.009
R19472 vp_p.n19378 vp_p.n19377 0.009
R19473 vp_p.n19392 vp_p.n19391 0.009
R19474 vp_p.n19406 vp_p.n19405 0.009
R19475 vp_p.n19420 vp_p.n19419 0.009
R19476 vp_p.n19434 vp_p.n19433 0.009
R19477 vp_p.n19448 vp_p.n19447 0.009
R19478 vp_p.n19462 vp_p.n19461 0.009
R19479 vp_p.n19476 vp_p.n19475 0.009
R19480 vp_p.n19490 vp_p.n19489 0.009
R19481 vp_p.n19504 vp_p.n19503 0.009
R19482 vp_p.n19518 vp_p.n19517 0.009
R19483 vp_p.n19532 vp_p.n19531 0.009
R19484 vp_p.n19546 vp_p.n19545 0.009
R19485 vp_p.n19560 vp_p.n19559 0.009
R19486 vp_p.n19574 vp_p.n19573 0.009
R19487 vp_p.n19588 vp_p.n19587 0.009
R19488 vp_p.n19602 vp_p.n19601 0.009
R19489 vp_p.n19616 vp_p.n19615 0.009
R19490 vp_p.n19630 vp_p.n19629 0.009
R19491 vp_p.n19644 vp_p.n19643 0.009
R19492 vp_p.n19658 vp_p.n19657 0.009
R19493 vp_p.n19672 vp_p.n19671 0.009
R19494 vp_p.n19686 vp_p.n19685 0.009
R19495 vp_p.n19700 vp_p.n19699 0.009
R19496 vp_p.n19714 vp_p.n19713 0.009
R19497 vp_p.n19728 vp_p.n19727 0.009
R19498 vp_p.n19742 vp_p.n19741 0.009
R19499 vp_p.n19756 vp_p.n19755 0.009
R19500 vp_p.n19770 vp_p.n19769 0.009
R19501 vp_p.n19784 vp_p.n19783 0.009
R19502 vp_p.n19798 vp_p.n19797 0.009
R19503 vp_p.n19812 vp_p.n19811 0.009
R19504 vp_p.n19826 vp_p.n19825 0.009
R19505 vp_p.n19840 vp_p.n19839 0.009
R19506 vp_p.n19854 vp_p.n19853 0.009
R19507 vp_p.n19868 vp_p.n19867 0.009
R19508 vp_p.n19882 vp_p.n19881 0.009
R19509 vp_p.n19896 vp_p.n19895 0.009
R19510 vp_p.n19910 vp_p.n19909 0.009
R19511 vp_p.n19924 vp_p.n19923 0.009
R19512 vp_p.n19938 vp_p.n19937 0.009
R19513 vp_p.n19952 vp_p.n19951 0.009
R19514 vp_p.n19966 vp_p.n19965 0.009
R19515 vp_p.n19980 vp_p.n19979 0.009
R19516 vp_p.n19994 vp_p.n19993 0.009
R19517 vp_p.n20008 vp_p.n20007 0.009
R19518 vp_p.n20022 vp_p.n20021 0.009
R19519 vp_p.n20036 vp_p.n20035 0.009
R19520 vp_p.n20050 vp_p.n20049 0.009
R19521 vp_p.n20064 vp_p.n20063 0.009
R19522 vp_p.n20078 vp_p.n20077 0.009
R19523 vp_p.n20092 vp_p.n20091 0.009
R19524 vp_p.n20106 vp_p.n20105 0.009
R19525 vp_p.n20120 vp_p.n20119 0.009
R19526 vp_p.n20134 vp_p.n20133 0.009
R19527 vp_p.n1903 vp_p.n1902 0.009
R19528 vp_p.n1917 vp_p.n1916 0.009
R19529 vp_p.n1931 vp_p.n1930 0.009
R19530 vp_p.n1945 vp_p.n1944 0.009
R19531 vp_p.n1959 vp_p.n1958 0.009
R19532 vp_p.n1973 vp_p.n1972 0.009
R19533 vp_p.n1987 vp_p.n1986 0.009
R19534 vp_p.n2001 vp_p.n2000 0.009
R19535 vp_p.n2015 vp_p.n2014 0.009
R19536 vp_p.n2029 vp_p.n2028 0.009
R19537 vp_p.n2043 vp_p.n2042 0.009
R19538 vp_p.n2057 vp_p.n2056 0.009
R19539 vp_p.n2071 vp_p.n2070 0.009
R19540 vp_p.n2085 vp_p.n2084 0.009
R19541 vp_p.n2099 vp_p.n2098 0.009
R19542 vp_p.n2113 vp_p.n2112 0.009
R19543 vp_p.n2127 vp_p.n2126 0.009
R19544 vp_p.n2141 vp_p.n2140 0.009
R19545 vp_p.n2155 vp_p.n2154 0.009
R19546 vp_p.n2169 vp_p.n2168 0.009
R19547 vp_p.n2183 vp_p.n2182 0.009
R19548 vp_p.n2197 vp_p.n2196 0.009
R19549 vp_p.n2211 vp_p.n2210 0.009
R19550 vp_p.n2225 vp_p.n2224 0.009
R19551 vp_p.n2239 vp_p.n2238 0.009
R19552 vp_p.n2253 vp_p.n2252 0.009
R19553 vp_p.n2267 vp_p.n2266 0.009
R19554 vp_p.n2281 vp_p.n2280 0.009
R19555 vp_p.n2295 vp_p.n2294 0.009
R19556 vp_p.n2309 vp_p.n2308 0.009
R19557 vp_p.n2323 vp_p.n2322 0.009
R19558 vp_p.n2337 vp_p.n2336 0.009
R19559 vp_p.n2351 vp_p.n2350 0.009
R19560 vp_p.n2365 vp_p.n2364 0.009
R19561 vp_p.n2379 vp_p.n2378 0.009
R19562 vp_p.n2393 vp_p.n2392 0.009
R19563 vp_p.n2407 vp_p.n2406 0.009
R19564 vp_p.n2421 vp_p.n2420 0.009
R19565 vp_p.n2435 vp_p.n2434 0.009
R19566 vp_p.n2449 vp_p.n2448 0.009
R19567 vp_p.n2463 vp_p.n2462 0.009
R19568 vp_p.n2477 vp_p.n2476 0.009
R19569 vp_p.n2491 vp_p.n2490 0.009
R19570 vp_p.n2505 vp_p.n2504 0.009
R19571 vp_p.n2519 vp_p.n2518 0.009
R19572 vp_p.n2533 vp_p.n2532 0.009
R19573 vp_p.n2547 vp_p.n2546 0.009
R19574 vp_p.n2561 vp_p.n2560 0.009
R19575 vp_p.n2575 vp_p.n2574 0.009
R19576 vp_p.n2589 vp_p.n2588 0.009
R19577 vp_p.n2603 vp_p.n2602 0.009
R19578 vp_p.n2617 vp_p.n2616 0.009
R19579 vp_p.n2631 vp_p.n2630 0.009
R19580 vp_p.n2645 vp_p.n2644 0.009
R19581 vp_p.n2659 vp_p.n2658 0.009
R19582 vp_p.n2673 vp_p.n2672 0.009
R19583 vp_p.n2687 vp_p.n2686 0.009
R19584 vp_p.n2701 vp_p.n2700 0.009
R19585 vp_p.n2715 vp_p.n2714 0.009
R19586 vp_p.n2729 vp_p.n2728 0.009
R19587 vp_p.n2743 vp_p.n2742 0.009
R19588 vp_p.n2757 vp_p.n2756 0.009
R19589 vp_p.n2771 vp_p.n2770 0.009
R19590 vp_p.n2785 vp_p.n2784 0.009
R19591 vp_p.n2799 vp_p.n2798 0.009
R19592 vp_p.n2813 vp_p.n2812 0.009
R19593 vp_p.n2827 vp_p.n2826 0.009
R19594 vp_p.n2841 vp_p.n2840 0.009
R19595 vp_p.n2855 vp_p.n2854 0.009
R19596 vp_p.n2869 vp_p.n2868 0.009
R19597 vp_p.n20607 vp_p.n20606 0.009
R19598 vp_p.n20621 vp_p.n20620 0.009
R19599 vp_p.n20635 vp_p.n20634 0.009
R19600 vp_p.n20649 vp_p.n20648 0.009
R19601 vp_p.n20663 vp_p.n20662 0.009
R19602 vp_p.n20677 vp_p.n20676 0.009
R19603 vp_p.n20691 vp_p.n20690 0.009
R19604 vp_p.n20705 vp_p.n20704 0.009
R19605 vp_p.n20719 vp_p.n20718 0.009
R19606 vp_p.n20733 vp_p.n20732 0.009
R19607 vp_p.n20747 vp_p.n20746 0.009
R19608 vp_p.n20761 vp_p.n20760 0.009
R19609 vp_p.n20775 vp_p.n20774 0.009
R19610 vp_p.n20789 vp_p.n20788 0.009
R19611 vp_p.n20803 vp_p.n20802 0.009
R19612 vp_p.n20817 vp_p.n20816 0.009
R19613 vp_p.n20831 vp_p.n20830 0.009
R19614 vp_p.n20845 vp_p.n20844 0.009
R19615 vp_p.n20859 vp_p.n20858 0.009
R19616 vp_p.n20873 vp_p.n20872 0.009
R19617 vp_p.n20887 vp_p.n20886 0.009
R19618 vp_p.n20901 vp_p.n20900 0.009
R19619 vp_p.n20915 vp_p.n20914 0.009
R19620 vp_p.n20929 vp_p.n20928 0.009
R19621 vp_p.n20943 vp_p.n20942 0.009
R19622 vp_p.n20957 vp_p.n20956 0.009
R19623 vp_p.n20971 vp_p.n20970 0.009
R19624 vp_p.n20985 vp_p.n20984 0.009
R19625 vp_p.n20999 vp_p.n20998 0.009
R19626 vp_p.n21013 vp_p.n21012 0.009
R19627 vp_p.n21027 vp_p.n21026 0.009
R19628 vp_p.n21041 vp_p.n21040 0.009
R19629 vp_p.n21055 vp_p.n21054 0.009
R19630 vp_p.n21069 vp_p.n21068 0.009
R19631 vp_p.n21083 vp_p.n21082 0.009
R19632 vp_p.n21097 vp_p.n21096 0.009
R19633 vp_p.n21111 vp_p.n21110 0.009
R19634 vp_p.n21125 vp_p.n21124 0.009
R19635 vp_p.n21139 vp_p.n21138 0.009
R19636 vp_p.n21153 vp_p.n21152 0.009
R19637 vp_p.n21167 vp_p.n21166 0.009
R19638 vp_p.n21181 vp_p.n21180 0.009
R19639 vp_p.n21195 vp_p.n21194 0.009
R19640 vp_p.n21209 vp_p.n21208 0.009
R19641 vp_p.n21223 vp_p.n21222 0.009
R19642 vp_p.n21237 vp_p.n21236 0.009
R19643 vp_p.n21251 vp_p.n21250 0.009
R19644 vp_p.n21265 vp_p.n21264 0.009
R19645 vp_p.n21279 vp_p.n21278 0.009
R19646 vp_p.n21293 vp_p.n21292 0.009
R19647 vp_p.n21307 vp_p.n21306 0.009
R19648 vp_p.n21321 vp_p.n21320 0.009
R19649 vp_p.n21335 vp_p.n21334 0.009
R19650 vp_p.n21349 vp_p.n21348 0.009
R19651 vp_p.n21363 vp_p.n21362 0.009
R19652 vp_p.n21377 vp_p.n21376 0.009
R19653 vp_p.n21391 vp_p.n21390 0.009
R19654 vp_p.n21405 vp_p.n21404 0.009
R19655 vp_p.n21419 vp_p.n21418 0.009
R19656 vp_p.n21433 vp_p.n21432 0.009
R19657 vp_p.n21447 vp_p.n21446 0.009
R19658 vp_p.n21461 vp_p.n21460 0.009
R19659 vp_p.n21475 vp_p.n21474 0.009
R19660 vp_p.n21489 vp_p.n21488 0.009
R19661 vp_p.n21503 vp_p.n21502 0.009
R19662 vp_p.n21517 vp_p.n21516 0.009
R19663 vp_p.n21531 vp_p.n21530 0.009
R19664 vp_p.n21545 vp_p.n21544 0.009
R19665 vp_p.n21559 vp_p.n21558 0.009
R19666 vp_p.n21573 vp_p.n21572 0.009
R19667 vp_p.n3328 vp_p.n3327 0.009
R19668 vp_p.n3342 vp_p.n3341 0.009
R19669 vp_p.n3356 vp_p.n3355 0.009
R19670 vp_p.n3370 vp_p.n3369 0.009
R19671 vp_p.n3384 vp_p.n3383 0.009
R19672 vp_p.n3398 vp_p.n3397 0.009
R19673 vp_p.n3412 vp_p.n3411 0.009
R19674 vp_p.n3426 vp_p.n3425 0.009
R19675 vp_p.n3440 vp_p.n3439 0.009
R19676 vp_p.n3454 vp_p.n3453 0.009
R19677 vp_p.n3468 vp_p.n3467 0.009
R19678 vp_p.n3482 vp_p.n3481 0.009
R19679 vp_p.n3496 vp_p.n3495 0.009
R19680 vp_p.n3510 vp_p.n3509 0.009
R19681 vp_p.n3524 vp_p.n3523 0.009
R19682 vp_p.n3538 vp_p.n3537 0.009
R19683 vp_p.n3552 vp_p.n3551 0.009
R19684 vp_p.n3566 vp_p.n3565 0.009
R19685 vp_p.n3580 vp_p.n3579 0.009
R19686 vp_p.n3594 vp_p.n3593 0.009
R19687 vp_p.n3608 vp_p.n3607 0.009
R19688 vp_p.n3622 vp_p.n3621 0.009
R19689 vp_p.n3636 vp_p.n3635 0.009
R19690 vp_p.n3650 vp_p.n3649 0.009
R19691 vp_p.n3664 vp_p.n3663 0.009
R19692 vp_p.n3678 vp_p.n3677 0.009
R19693 vp_p.n3692 vp_p.n3691 0.009
R19694 vp_p.n3706 vp_p.n3705 0.009
R19695 vp_p.n3720 vp_p.n3719 0.009
R19696 vp_p.n3734 vp_p.n3733 0.009
R19697 vp_p.n3748 vp_p.n3747 0.009
R19698 vp_p.n3762 vp_p.n3761 0.009
R19699 vp_p.n3776 vp_p.n3775 0.009
R19700 vp_p.n3790 vp_p.n3789 0.009
R19701 vp_p.n3804 vp_p.n3803 0.009
R19702 vp_p.n3818 vp_p.n3817 0.009
R19703 vp_p.n3832 vp_p.n3831 0.009
R19704 vp_p.n3846 vp_p.n3845 0.009
R19705 vp_p.n3860 vp_p.n3859 0.009
R19706 vp_p.n3874 vp_p.n3873 0.009
R19707 vp_p.n3888 vp_p.n3887 0.009
R19708 vp_p.n3902 vp_p.n3901 0.009
R19709 vp_p.n3916 vp_p.n3915 0.009
R19710 vp_p.n3930 vp_p.n3929 0.009
R19711 vp_p.n3944 vp_p.n3943 0.009
R19712 vp_p.n3958 vp_p.n3957 0.009
R19713 vp_p.n3972 vp_p.n3971 0.009
R19714 vp_p.n3986 vp_p.n3985 0.009
R19715 vp_p.n4000 vp_p.n3999 0.009
R19716 vp_p.n4014 vp_p.n4013 0.009
R19717 vp_p.n4028 vp_p.n4027 0.009
R19718 vp_p.n4042 vp_p.n4041 0.009
R19719 vp_p.n4056 vp_p.n4055 0.009
R19720 vp_p.n4070 vp_p.n4069 0.009
R19721 vp_p.n4084 vp_p.n4083 0.009
R19722 vp_p.n4098 vp_p.n4097 0.009
R19723 vp_p.n4112 vp_p.n4111 0.009
R19724 vp_p.n4126 vp_p.n4125 0.009
R19725 vp_p.n4140 vp_p.n4139 0.009
R19726 vp_p.n4154 vp_p.n4153 0.009
R19727 vp_p.n4168 vp_p.n4167 0.009
R19728 vp_p.n4182 vp_p.n4181 0.009
R19729 vp_p.n4196 vp_p.n4195 0.009
R19730 vp_p.n4210 vp_p.n4209 0.009
R19731 vp_p.n4224 vp_p.n4223 0.009
R19732 vp_p.n4238 vp_p.n4237 0.009
R19733 vp_p.n4252 vp_p.n4251 0.009
R19734 vp_p.n4266 vp_p.n4265 0.009
R19735 vp_p.n4280 vp_p.n4279 0.009
R19736 vp_p.n4294 vp_p.n4293 0.009
R19737 vp_p.n4308 vp_p.n4307 0.009
R19738 vp_p.n22031 vp_p.n22030 0.009
R19739 vp_p.n22045 vp_p.n22044 0.009
R19740 vp_p.n22059 vp_p.n22058 0.009
R19741 vp_p.n22073 vp_p.n22072 0.009
R19742 vp_p.n22087 vp_p.n22086 0.009
R19743 vp_p.n22101 vp_p.n22100 0.009
R19744 vp_p.n22115 vp_p.n22114 0.009
R19745 vp_p.n22129 vp_p.n22128 0.009
R19746 vp_p.n22143 vp_p.n22142 0.009
R19747 vp_p.n22157 vp_p.n22156 0.009
R19748 vp_p.n22171 vp_p.n22170 0.009
R19749 vp_p.n22185 vp_p.n22184 0.009
R19750 vp_p.n22199 vp_p.n22198 0.009
R19751 vp_p.n22213 vp_p.n22212 0.009
R19752 vp_p.n22227 vp_p.n22226 0.009
R19753 vp_p.n22241 vp_p.n22240 0.009
R19754 vp_p.n22255 vp_p.n22254 0.009
R19755 vp_p.n22269 vp_p.n22268 0.009
R19756 vp_p.n22283 vp_p.n22282 0.009
R19757 vp_p.n22297 vp_p.n22296 0.009
R19758 vp_p.n22311 vp_p.n22310 0.009
R19759 vp_p.n22325 vp_p.n22324 0.009
R19760 vp_p.n22339 vp_p.n22338 0.009
R19761 vp_p.n22353 vp_p.n22352 0.009
R19762 vp_p.n22367 vp_p.n22366 0.009
R19763 vp_p.n22381 vp_p.n22380 0.009
R19764 vp_p.n22395 vp_p.n22394 0.009
R19765 vp_p.n22409 vp_p.n22408 0.009
R19766 vp_p.n22423 vp_p.n22422 0.009
R19767 vp_p.n22437 vp_p.n22436 0.009
R19768 vp_p.n22451 vp_p.n22450 0.009
R19769 vp_p.n22465 vp_p.n22464 0.009
R19770 vp_p.n22479 vp_p.n22478 0.009
R19771 vp_p.n22493 vp_p.n22492 0.009
R19772 vp_p.n22507 vp_p.n22506 0.009
R19773 vp_p.n22521 vp_p.n22520 0.009
R19774 vp_p.n22535 vp_p.n22534 0.009
R19775 vp_p.n22549 vp_p.n22548 0.009
R19776 vp_p.n22563 vp_p.n22562 0.009
R19777 vp_p.n22577 vp_p.n22576 0.009
R19778 vp_p.n22591 vp_p.n22590 0.009
R19779 vp_p.n22605 vp_p.n22604 0.009
R19780 vp_p.n22619 vp_p.n22618 0.009
R19781 vp_p.n22633 vp_p.n22632 0.009
R19782 vp_p.n22647 vp_p.n22646 0.009
R19783 vp_p.n22661 vp_p.n22660 0.009
R19784 vp_p.n22675 vp_p.n22674 0.009
R19785 vp_p.n22689 vp_p.n22688 0.009
R19786 vp_p.n22703 vp_p.n22702 0.009
R19787 vp_p.n22717 vp_p.n22716 0.009
R19788 vp_p.n22731 vp_p.n22730 0.009
R19789 vp_p.n22745 vp_p.n22744 0.009
R19790 vp_p.n22759 vp_p.n22758 0.009
R19791 vp_p.n22773 vp_p.n22772 0.009
R19792 vp_p.n22787 vp_p.n22786 0.009
R19793 vp_p.n22801 vp_p.n22800 0.009
R19794 vp_p.n22815 vp_p.n22814 0.009
R19795 vp_p.n22829 vp_p.n22828 0.009
R19796 vp_p.n22843 vp_p.n22842 0.009
R19797 vp_p.n22857 vp_p.n22856 0.009
R19798 vp_p.n22871 vp_p.n22870 0.009
R19799 vp_p.n22885 vp_p.n22884 0.009
R19800 vp_p.n22899 vp_p.n22898 0.009
R19801 vp_p.n22913 vp_p.n22912 0.009
R19802 vp_p.n22927 vp_p.n22926 0.009
R19803 vp_p.n22941 vp_p.n22940 0.009
R19804 vp_p.n22955 vp_p.n22954 0.009
R19805 vp_p.n22969 vp_p.n22968 0.009
R19806 vp_p.n22983 vp_p.n22982 0.009
R19807 vp_p.n22997 vp_p.n22996 0.009
R19808 vp_p.n23011 vp_p.n23010 0.009
R19809 vp_p.n4752 vp_p.n4751 0.009
R19810 vp_p.n4766 vp_p.n4765 0.009
R19811 vp_p.n4780 vp_p.n4779 0.009
R19812 vp_p.n4794 vp_p.n4793 0.009
R19813 vp_p.n4808 vp_p.n4807 0.009
R19814 vp_p.n4822 vp_p.n4821 0.009
R19815 vp_p.n4836 vp_p.n4835 0.009
R19816 vp_p.n4850 vp_p.n4849 0.009
R19817 vp_p.n4864 vp_p.n4863 0.009
R19818 vp_p.n4878 vp_p.n4877 0.009
R19819 vp_p.n4892 vp_p.n4891 0.009
R19820 vp_p.n4906 vp_p.n4905 0.009
R19821 vp_p.n4920 vp_p.n4919 0.009
R19822 vp_p.n4934 vp_p.n4933 0.009
R19823 vp_p.n4948 vp_p.n4947 0.009
R19824 vp_p.n4962 vp_p.n4961 0.009
R19825 vp_p.n4976 vp_p.n4975 0.009
R19826 vp_p.n4990 vp_p.n4989 0.009
R19827 vp_p.n5004 vp_p.n5003 0.009
R19828 vp_p.n5018 vp_p.n5017 0.009
R19829 vp_p.n5032 vp_p.n5031 0.009
R19830 vp_p.n5046 vp_p.n5045 0.009
R19831 vp_p.n5060 vp_p.n5059 0.009
R19832 vp_p.n5074 vp_p.n5073 0.009
R19833 vp_p.n5088 vp_p.n5087 0.009
R19834 vp_p.n5102 vp_p.n5101 0.009
R19835 vp_p.n5116 vp_p.n5115 0.009
R19836 vp_p.n5130 vp_p.n5129 0.009
R19837 vp_p.n5144 vp_p.n5143 0.009
R19838 vp_p.n5158 vp_p.n5157 0.009
R19839 vp_p.n5172 vp_p.n5171 0.009
R19840 vp_p.n5186 vp_p.n5185 0.009
R19841 vp_p.n5200 vp_p.n5199 0.009
R19842 vp_p.n5214 vp_p.n5213 0.009
R19843 vp_p.n5228 vp_p.n5227 0.009
R19844 vp_p.n5242 vp_p.n5241 0.009
R19845 vp_p.n5256 vp_p.n5255 0.009
R19846 vp_p.n5270 vp_p.n5269 0.009
R19847 vp_p.n5284 vp_p.n5283 0.009
R19848 vp_p.n5298 vp_p.n5297 0.009
R19849 vp_p.n5312 vp_p.n5311 0.009
R19850 vp_p.n5326 vp_p.n5325 0.009
R19851 vp_p.n5340 vp_p.n5339 0.009
R19852 vp_p.n5354 vp_p.n5353 0.009
R19853 vp_p.n5368 vp_p.n5367 0.009
R19854 vp_p.n5382 vp_p.n5381 0.009
R19855 vp_p.n5396 vp_p.n5395 0.009
R19856 vp_p.n5410 vp_p.n5409 0.009
R19857 vp_p.n5424 vp_p.n5423 0.009
R19858 vp_p.n5438 vp_p.n5437 0.009
R19859 vp_p.n5452 vp_p.n5451 0.009
R19860 vp_p.n5466 vp_p.n5465 0.009
R19861 vp_p.n5480 vp_p.n5479 0.009
R19862 vp_p.n5494 vp_p.n5493 0.009
R19863 vp_p.n5508 vp_p.n5507 0.009
R19864 vp_p.n5522 vp_p.n5521 0.009
R19865 vp_p.n5536 vp_p.n5535 0.009
R19866 vp_p.n5550 vp_p.n5549 0.009
R19867 vp_p.n5564 vp_p.n5563 0.009
R19868 vp_p.n5578 vp_p.n5577 0.009
R19869 vp_p.n5592 vp_p.n5591 0.009
R19870 vp_p.n5606 vp_p.n5605 0.009
R19871 vp_p.n5620 vp_p.n5619 0.009
R19872 vp_p.n5634 vp_p.n5633 0.009
R19873 vp_p.n5648 vp_p.n5647 0.009
R19874 vp_p.n5662 vp_p.n5661 0.009
R19875 vp_p.n5676 vp_p.n5675 0.009
R19876 vp_p.n5690 vp_p.n5689 0.009
R19877 vp_p.n5704 vp_p.n5703 0.009
R19878 vp_p.n5718 vp_p.n5717 0.009
R19879 vp_p.n5732 vp_p.n5731 0.009
R19880 vp_p.n5746 vp_p.n5745 0.009
R19881 vp_p.n23454 vp_p.n23453 0.009
R19882 vp_p.n23468 vp_p.n23467 0.009
R19883 vp_p.n23482 vp_p.n23481 0.009
R19884 vp_p.n23496 vp_p.n23495 0.009
R19885 vp_p.n23510 vp_p.n23509 0.009
R19886 vp_p.n23524 vp_p.n23523 0.009
R19887 vp_p.n23538 vp_p.n23537 0.009
R19888 vp_p.n23552 vp_p.n23551 0.009
R19889 vp_p.n23566 vp_p.n23565 0.009
R19890 vp_p.n23580 vp_p.n23579 0.009
R19891 vp_p.n23594 vp_p.n23593 0.009
R19892 vp_p.n23608 vp_p.n23607 0.009
R19893 vp_p.n23622 vp_p.n23621 0.009
R19894 vp_p.n23636 vp_p.n23635 0.009
R19895 vp_p.n23650 vp_p.n23649 0.009
R19896 vp_p.n23664 vp_p.n23663 0.009
R19897 vp_p.n23678 vp_p.n23677 0.009
R19898 vp_p.n23692 vp_p.n23691 0.009
R19899 vp_p.n23706 vp_p.n23705 0.009
R19900 vp_p.n23720 vp_p.n23719 0.009
R19901 vp_p.n23734 vp_p.n23733 0.009
R19902 vp_p.n23748 vp_p.n23747 0.009
R19903 vp_p.n23762 vp_p.n23761 0.009
R19904 vp_p.n23776 vp_p.n23775 0.009
R19905 vp_p.n23790 vp_p.n23789 0.009
R19906 vp_p.n23804 vp_p.n23803 0.009
R19907 vp_p.n23818 vp_p.n23817 0.009
R19908 vp_p.n23832 vp_p.n23831 0.009
R19909 vp_p.n23846 vp_p.n23845 0.009
R19910 vp_p.n23860 vp_p.n23859 0.009
R19911 vp_p.n23874 vp_p.n23873 0.009
R19912 vp_p.n23888 vp_p.n23887 0.009
R19913 vp_p.n23902 vp_p.n23901 0.009
R19914 vp_p.n23916 vp_p.n23915 0.009
R19915 vp_p.n23930 vp_p.n23929 0.009
R19916 vp_p.n23944 vp_p.n23943 0.009
R19917 vp_p.n23958 vp_p.n23957 0.009
R19918 vp_p.n23972 vp_p.n23971 0.009
R19919 vp_p.n23986 vp_p.n23985 0.009
R19920 vp_p.n24000 vp_p.n23999 0.009
R19921 vp_p.n24014 vp_p.n24013 0.009
R19922 vp_p.n24028 vp_p.n24027 0.009
R19923 vp_p.n24042 vp_p.n24041 0.009
R19924 vp_p.n24056 vp_p.n24055 0.009
R19925 vp_p.n24070 vp_p.n24069 0.009
R19926 vp_p.n24084 vp_p.n24083 0.009
R19927 vp_p.n24098 vp_p.n24097 0.009
R19928 vp_p.n24112 vp_p.n24111 0.009
R19929 vp_p.n24126 vp_p.n24125 0.009
R19930 vp_p.n24140 vp_p.n24139 0.009
R19931 vp_p.n24154 vp_p.n24153 0.009
R19932 vp_p.n24168 vp_p.n24167 0.009
R19933 vp_p.n24182 vp_p.n24181 0.009
R19934 vp_p.n24196 vp_p.n24195 0.009
R19935 vp_p.n24210 vp_p.n24209 0.009
R19936 vp_p.n24224 vp_p.n24223 0.009
R19937 vp_p.n24238 vp_p.n24237 0.009
R19938 vp_p.n24252 vp_p.n24251 0.009
R19939 vp_p.n24266 vp_p.n24265 0.009
R19940 vp_p.n24280 vp_p.n24279 0.009
R19941 vp_p.n24294 vp_p.n24293 0.009
R19942 vp_p.n24308 vp_p.n24307 0.009
R19943 vp_p.n24322 vp_p.n24321 0.009
R19944 vp_p.n24336 vp_p.n24335 0.009
R19945 vp_p.n24350 vp_p.n24349 0.009
R19946 vp_p.n24364 vp_p.n24363 0.009
R19947 vp_p.n24378 vp_p.n24377 0.009
R19948 vp_p.n24392 vp_p.n24391 0.009
R19949 vp_p.n24406 vp_p.n24405 0.009
R19950 vp_p.n24420 vp_p.n24419 0.009
R19951 vp_p.n24434 vp_p.n24433 0.009
R19952 vp_p.n24448 vp_p.n24447 0.009
R19953 vp_p.n6175 vp_p.n6174 0.009
R19954 vp_p.n6189 vp_p.n6188 0.009
R19955 vp_p.n6203 vp_p.n6202 0.009
R19956 vp_p.n6217 vp_p.n6216 0.009
R19957 vp_p.n6231 vp_p.n6230 0.009
R19958 vp_p.n6245 vp_p.n6244 0.009
R19959 vp_p.n6259 vp_p.n6258 0.009
R19960 vp_p.n6273 vp_p.n6272 0.009
R19961 vp_p.n6287 vp_p.n6286 0.009
R19962 vp_p.n6301 vp_p.n6300 0.009
R19963 vp_p.n6315 vp_p.n6314 0.009
R19964 vp_p.n6329 vp_p.n6328 0.009
R19965 vp_p.n6343 vp_p.n6342 0.009
R19966 vp_p.n6357 vp_p.n6356 0.009
R19967 vp_p.n6371 vp_p.n6370 0.009
R19968 vp_p.n6385 vp_p.n6384 0.009
R19969 vp_p.n6399 vp_p.n6398 0.009
R19970 vp_p.n6413 vp_p.n6412 0.009
R19971 vp_p.n6427 vp_p.n6426 0.009
R19972 vp_p.n6441 vp_p.n6440 0.009
R19973 vp_p.n6455 vp_p.n6454 0.009
R19974 vp_p.n6469 vp_p.n6468 0.009
R19975 vp_p.n6483 vp_p.n6482 0.009
R19976 vp_p.n6497 vp_p.n6496 0.009
R19977 vp_p.n6511 vp_p.n6510 0.009
R19978 vp_p.n6525 vp_p.n6524 0.009
R19979 vp_p.n6539 vp_p.n6538 0.009
R19980 vp_p.n6553 vp_p.n6552 0.009
R19981 vp_p.n6567 vp_p.n6566 0.009
R19982 vp_p.n6581 vp_p.n6580 0.009
R19983 vp_p.n6595 vp_p.n6594 0.009
R19984 vp_p.n6609 vp_p.n6608 0.009
R19985 vp_p.n6623 vp_p.n6622 0.009
R19986 vp_p.n6637 vp_p.n6636 0.009
R19987 vp_p.n6651 vp_p.n6650 0.009
R19988 vp_p.n6665 vp_p.n6664 0.009
R19989 vp_p.n6679 vp_p.n6678 0.009
R19990 vp_p.n6693 vp_p.n6692 0.009
R19991 vp_p.n6707 vp_p.n6706 0.009
R19992 vp_p.n6721 vp_p.n6720 0.009
R19993 vp_p.n6735 vp_p.n6734 0.009
R19994 vp_p.n6749 vp_p.n6748 0.009
R19995 vp_p.n6763 vp_p.n6762 0.009
R19996 vp_p.n6777 vp_p.n6776 0.009
R19997 vp_p.n6791 vp_p.n6790 0.009
R19998 vp_p.n6805 vp_p.n6804 0.009
R19999 vp_p.n6819 vp_p.n6818 0.009
R20000 vp_p.n6833 vp_p.n6832 0.009
R20001 vp_p.n6847 vp_p.n6846 0.009
R20002 vp_p.n6861 vp_p.n6860 0.009
R20003 vp_p.n6875 vp_p.n6874 0.009
R20004 vp_p.n6889 vp_p.n6888 0.009
R20005 vp_p.n6903 vp_p.n6902 0.009
R20006 vp_p.n6917 vp_p.n6916 0.009
R20007 vp_p.n6931 vp_p.n6930 0.009
R20008 vp_p.n6945 vp_p.n6944 0.009
R20009 vp_p.n6959 vp_p.n6958 0.009
R20010 vp_p.n6973 vp_p.n6972 0.009
R20011 vp_p.n6987 vp_p.n6986 0.009
R20012 vp_p.n7001 vp_p.n7000 0.009
R20013 vp_p.n7015 vp_p.n7014 0.009
R20014 vp_p.n7029 vp_p.n7028 0.009
R20015 vp_p.n7043 vp_p.n7042 0.009
R20016 vp_p.n7057 vp_p.n7056 0.009
R20017 vp_p.n7071 vp_p.n7070 0.009
R20018 vp_p.n7085 vp_p.n7084 0.009
R20019 vp_p.n7099 vp_p.n7098 0.009
R20020 vp_p.n7113 vp_p.n7112 0.009
R20021 vp_p.n7127 vp_p.n7126 0.009
R20022 vp_p.n7141 vp_p.n7140 0.009
R20023 vp_p.n7155 vp_p.n7154 0.009
R20024 vp_p.n7169 vp_p.n7168 0.009
R20025 vp_p.n7183 vp_p.n7182 0.009
R20026 vp_p.n24876 vp_p.n24875 0.009
R20027 vp_p.n24890 vp_p.n24889 0.009
R20028 vp_p.n24904 vp_p.n24903 0.009
R20029 vp_p.n24918 vp_p.n24917 0.009
R20030 vp_p.n24932 vp_p.n24931 0.009
R20031 vp_p.n24946 vp_p.n24945 0.009
R20032 vp_p.n24960 vp_p.n24959 0.009
R20033 vp_p.n24974 vp_p.n24973 0.009
R20034 vp_p.n24988 vp_p.n24987 0.009
R20035 vp_p.n25002 vp_p.n25001 0.009
R20036 vp_p.n25016 vp_p.n25015 0.009
R20037 vp_p.n25030 vp_p.n25029 0.009
R20038 vp_p.n25044 vp_p.n25043 0.009
R20039 vp_p.n25058 vp_p.n25057 0.009
R20040 vp_p.n25072 vp_p.n25071 0.009
R20041 vp_p.n25086 vp_p.n25085 0.009
R20042 vp_p.n25100 vp_p.n25099 0.009
R20043 vp_p.n25114 vp_p.n25113 0.009
R20044 vp_p.n25128 vp_p.n25127 0.009
R20045 vp_p.n25142 vp_p.n25141 0.009
R20046 vp_p.n25156 vp_p.n25155 0.009
R20047 vp_p.n25170 vp_p.n25169 0.009
R20048 vp_p.n25184 vp_p.n25183 0.009
R20049 vp_p.n25198 vp_p.n25197 0.009
R20050 vp_p.n25212 vp_p.n25211 0.009
R20051 vp_p.n25226 vp_p.n25225 0.009
R20052 vp_p.n25240 vp_p.n25239 0.009
R20053 vp_p.n25254 vp_p.n25253 0.009
R20054 vp_p.n25268 vp_p.n25267 0.009
R20055 vp_p.n25282 vp_p.n25281 0.009
R20056 vp_p.n25296 vp_p.n25295 0.009
R20057 vp_p.n25310 vp_p.n25309 0.009
R20058 vp_p.n25324 vp_p.n25323 0.009
R20059 vp_p.n25338 vp_p.n25337 0.009
R20060 vp_p.n25352 vp_p.n25351 0.009
R20061 vp_p.n25366 vp_p.n25365 0.009
R20062 vp_p.n25380 vp_p.n25379 0.009
R20063 vp_p.n25394 vp_p.n25393 0.009
R20064 vp_p.n25408 vp_p.n25407 0.009
R20065 vp_p.n25422 vp_p.n25421 0.009
R20066 vp_p.n25436 vp_p.n25435 0.009
R20067 vp_p.n25450 vp_p.n25449 0.009
R20068 vp_p.n25464 vp_p.n25463 0.009
R20069 vp_p.n25478 vp_p.n25477 0.009
R20070 vp_p.n25492 vp_p.n25491 0.009
R20071 vp_p.n25506 vp_p.n25505 0.009
R20072 vp_p.n25520 vp_p.n25519 0.009
R20073 vp_p.n25534 vp_p.n25533 0.009
R20074 vp_p.n25548 vp_p.n25547 0.009
R20075 vp_p.n25562 vp_p.n25561 0.009
R20076 vp_p.n25576 vp_p.n25575 0.009
R20077 vp_p.n25590 vp_p.n25589 0.009
R20078 vp_p.n25604 vp_p.n25603 0.009
R20079 vp_p.n25618 vp_p.n25617 0.009
R20080 vp_p.n25632 vp_p.n25631 0.009
R20081 vp_p.n25646 vp_p.n25645 0.009
R20082 vp_p.n25660 vp_p.n25659 0.009
R20083 vp_p.n25674 vp_p.n25673 0.009
R20084 vp_p.n25688 vp_p.n25687 0.009
R20085 vp_p.n25702 vp_p.n25701 0.009
R20086 vp_p.n25716 vp_p.n25715 0.009
R20087 vp_p.n25730 vp_p.n25729 0.009
R20088 vp_p.n25744 vp_p.n25743 0.009
R20089 vp_p.n25758 vp_p.n25757 0.009
R20090 vp_p.n25772 vp_p.n25771 0.009
R20091 vp_p.n25786 vp_p.n25785 0.009
R20092 vp_p.n25800 vp_p.n25799 0.009
R20093 vp_p.n25814 vp_p.n25813 0.009
R20094 vp_p.n25828 vp_p.n25827 0.009
R20095 vp_p.n25842 vp_p.n25841 0.009
R20096 vp_p.n25856 vp_p.n25855 0.009
R20097 vp_p.n25870 vp_p.n25869 0.009
R20098 vp_p.n25884 vp_p.n25883 0.009
R20099 vp_p.n7597 vp_p.n7596 0.009
R20100 vp_p.n7611 vp_p.n7610 0.009
R20101 vp_p.n7625 vp_p.n7624 0.009
R20102 vp_p.n7639 vp_p.n7638 0.009
R20103 vp_p.n7653 vp_p.n7652 0.009
R20104 vp_p.n7667 vp_p.n7666 0.009
R20105 vp_p.n7681 vp_p.n7680 0.009
R20106 vp_p.n7695 vp_p.n7694 0.009
R20107 vp_p.n7709 vp_p.n7708 0.009
R20108 vp_p.n7723 vp_p.n7722 0.009
R20109 vp_p.n7737 vp_p.n7736 0.009
R20110 vp_p.n7751 vp_p.n7750 0.009
R20111 vp_p.n7765 vp_p.n7764 0.009
R20112 vp_p.n7779 vp_p.n7778 0.009
R20113 vp_p.n7793 vp_p.n7792 0.009
R20114 vp_p.n7807 vp_p.n7806 0.009
R20115 vp_p.n7821 vp_p.n7820 0.009
R20116 vp_p.n7835 vp_p.n7834 0.009
R20117 vp_p.n7849 vp_p.n7848 0.009
R20118 vp_p.n7863 vp_p.n7862 0.009
R20119 vp_p.n7877 vp_p.n7876 0.009
R20120 vp_p.n7891 vp_p.n7890 0.009
R20121 vp_p.n7905 vp_p.n7904 0.009
R20122 vp_p.n7919 vp_p.n7918 0.009
R20123 vp_p.n7933 vp_p.n7932 0.009
R20124 vp_p.n7947 vp_p.n7946 0.009
R20125 vp_p.n7961 vp_p.n7960 0.009
R20126 vp_p.n7975 vp_p.n7974 0.009
R20127 vp_p.n7989 vp_p.n7988 0.009
R20128 vp_p.n8003 vp_p.n8002 0.009
R20129 vp_p.n8017 vp_p.n8016 0.009
R20130 vp_p.n8031 vp_p.n8030 0.009
R20131 vp_p.n8045 vp_p.n8044 0.009
R20132 vp_p.n8059 vp_p.n8058 0.009
R20133 vp_p.n8073 vp_p.n8072 0.009
R20134 vp_p.n8087 vp_p.n8086 0.009
R20135 vp_p.n8101 vp_p.n8100 0.009
R20136 vp_p.n8115 vp_p.n8114 0.009
R20137 vp_p.n8129 vp_p.n8128 0.009
R20138 vp_p.n8143 vp_p.n8142 0.009
R20139 vp_p.n8157 vp_p.n8156 0.009
R20140 vp_p.n8171 vp_p.n8170 0.009
R20141 vp_p.n8185 vp_p.n8184 0.009
R20142 vp_p.n8199 vp_p.n8198 0.009
R20143 vp_p.n8213 vp_p.n8212 0.009
R20144 vp_p.n8227 vp_p.n8226 0.009
R20145 vp_p.n8241 vp_p.n8240 0.009
R20146 vp_p.n8255 vp_p.n8254 0.009
R20147 vp_p.n8269 vp_p.n8268 0.009
R20148 vp_p.n8283 vp_p.n8282 0.009
R20149 vp_p.n8297 vp_p.n8296 0.009
R20150 vp_p.n8311 vp_p.n8310 0.009
R20151 vp_p.n8325 vp_p.n8324 0.009
R20152 vp_p.n8339 vp_p.n8338 0.009
R20153 vp_p.n8353 vp_p.n8352 0.009
R20154 vp_p.n8367 vp_p.n8366 0.009
R20155 vp_p.n8381 vp_p.n8380 0.009
R20156 vp_p.n8395 vp_p.n8394 0.009
R20157 vp_p.n8409 vp_p.n8408 0.009
R20158 vp_p.n8423 vp_p.n8422 0.009
R20159 vp_p.n8437 vp_p.n8436 0.009
R20160 vp_p.n8451 vp_p.n8450 0.009
R20161 vp_p.n8465 vp_p.n8464 0.009
R20162 vp_p.n8479 vp_p.n8478 0.009
R20163 vp_p.n8493 vp_p.n8492 0.009
R20164 vp_p.n8507 vp_p.n8506 0.009
R20165 vp_p.n8521 vp_p.n8520 0.009
R20166 vp_p.n8535 vp_p.n8534 0.009
R20167 vp_p.n8549 vp_p.n8548 0.009
R20168 vp_p.n8563 vp_p.n8562 0.009
R20169 vp_p.n8577 vp_p.n8576 0.009
R20170 vp_p.n8591 vp_p.n8590 0.009
R20171 vp_p.n8605 vp_p.n8604 0.009
R20172 vp_p.n8619 vp_p.n8618 0.009
R20173 vp_p.n26301 vp_p.n26300 0.009
R20174 vp_p.n26315 vp_p.n26314 0.009
R20175 vp_p.n26329 vp_p.n26328 0.009
R20176 vp_p.n26343 vp_p.n26342 0.009
R20177 vp_p.n26357 vp_p.n26356 0.009
R20178 vp_p.n26371 vp_p.n26370 0.009
R20179 vp_p.n26385 vp_p.n26384 0.009
R20180 vp_p.n26399 vp_p.n26398 0.009
R20181 vp_p.n26413 vp_p.n26412 0.009
R20182 vp_p.n26427 vp_p.n26426 0.009
R20183 vp_p.n26441 vp_p.n26440 0.009
R20184 vp_p.n26455 vp_p.n26454 0.009
R20185 vp_p.n26469 vp_p.n26468 0.009
R20186 vp_p.n26483 vp_p.n26482 0.009
R20187 vp_p.n26497 vp_p.n26496 0.009
R20188 vp_p.n26511 vp_p.n26510 0.009
R20189 vp_p.n26525 vp_p.n26524 0.009
R20190 vp_p.n26539 vp_p.n26538 0.009
R20191 vp_p.n26553 vp_p.n26552 0.009
R20192 vp_p.n26567 vp_p.n26566 0.009
R20193 vp_p.n26581 vp_p.n26580 0.009
R20194 vp_p.n26595 vp_p.n26594 0.009
R20195 vp_p.n26609 vp_p.n26608 0.009
R20196 vp_p.n26623 vp_p.n26622 0.009
R20197 vp_p.n26637 vp_p.n26636 0.009
R20198 vp_p.n26651 vp_p.n26650 0.009
R20199 vp_p.n26665 vp_p.n26664 0.009
R20200 vp_p.n26679 vp_p.n26678 0.009
R20201 vp_p.n26693 vp_p.n26692 0.009
R20202 vp_p.n26707 vp_p.n26706 0.009
R20203 vp_p.n26721 vp_p.n26720 0.009
R20204 vp_p.n26735 vp_p.n26734 0.009
R20205 vp_p.n26749 vp_p.n26748 0.009
R20206 vp_p.n26763 vp_p.n26762 0.009
R20207 vp_p.n26777 vp_p.n26776 0.009
R20208 vp_p.n26791 vp_p.n26790 0.009
R20209 vp_p.n26805 vp_p.n26804 0.009
R20210 vp_p.n26819 vp_p.n26818 0.009
R20211 vp_p.n26833 vp_p.n26832 0.009
R20212 vp_p.n26847 vp_p.n26846 0.009
R20213 vp_p.n26861 vp_p.n26860 0.009
R20214 vp_p.n26875 vp_p.n26874 0.009
R20215 vp_p.n26889 vp_p.n26888 0.009
R20216 vp_p.n26903 vp_p.n26902 0.009
R20217 vp_p.n26917 vp_p.n26916 0.009
R20218 vp_p.n26931 vp_p.n26930 0.009
R20219 vp_p.n26945 vp_p.n26944 0.009
R20220 vp_p.n26959 vp_p.n26958 0.009
R20221 vp_p.n26973 vp_p.n26972 0.009
R20222 vp_p.n26987 vp_p.n26986 0.009
R20223 vp_p.n27001 vp_p.n27000 0.009
R20224 vp_p.n27015 vp_p.n27014 0.009
R20225 vp_p.n27029 vp_p.n27028 0.009
R20226 vp_p.n27043 vp_p.n27042 0.009
R20227 vp_p.n27057 vp_p.n27056 0.009
R20228 vp_p.n27071 vp_p.n27070 0.009
R20229 vp_p.n27085 vp_p.n27084 0.009
R20230 vp_p.n27099 vp_p.n27098 0.009
R20231 vp_p.n27113 vp_p.n27112 0.009
R20232 vp_p.n27127 vp_p.n27126 0.009
R20233 vp_p.n27141 vp_p.n27140 0.009
R20234 vp_p.n27155 vp_p.n27154 0.009
R20235 vp_p.n27169 vp_p.n27168 0.009
R20236 vp_p.n27183 vp_p.n27182 0.009
R20237 vp_p.n27197 vp_p.n27196 0.009
R20238 vp_p.n27211 vp_p.n27210 0.009
R20239 vp_p.n27225 vp_p.n27224 0.009
R20240 vp_p.n27239 vp_p.n27238 0.009
R20241 vp_p.n27253 vp_p.n27252 0.009
R20242 vp_p.n27267 vp_p.n27266 0.009
R20243 vp_p.n27281 vp_p.n27280 0.009
R20244 vp_p.n27295 vp_p.n27294 0.009
R20245 vp_p.n27309 vp_p.n27308 0.009
R20246 vp_p.n27323 vp_p.n27322 0.009
R20247 vp_p.n7576 vp_p.n7575 0.007
R20248 vp_p.n24860 vp_p.n24859 0.007
R20249 vp_p.n24865 vp_p.n24864 0.007
R20250 vp_p.n6159 vp_p.n6158 0.007
R20251 vp_p.n6164 vp_p.n6163 0.007
R20252 vp_p.n23438 vp_p.n23437 0.007
R20253 vp_p.n23443 vp_p.n23442 0.007
R20254 vp_p.n4736 vp_p.n4735 0.007
R20255 vp_p.n4741 vp_p.n4740 0.007
R20256 vp_p.n22015 vp_p.n22014 0.007
R20257 vp_p.n22020 vp_p.n22019 0.007
R20258 vp_p.n3312 vp_p.n3311 0.007
R20259 vp_p.n3317 vp_p.n3316 0.007
R20260 vp_p.n20591 vp_p.n20590 0.007
R20261 vp_p.n20596 vp_p.n20595 0.007
R20262 vp_p.n1887 vp_p.n1886 0.007
R20263 vp_p.n1892 vp_p.n1891 0.007
R20264 vp_p.n19166 vp_p.n19165 0.007
R20265 vp_p.n19171 vp_p.n19170 0.007
R20266 vp_p.n461 vp_p.n460 0.007
R20267 vp_p.n466 vp_p.n465 0.007
R20268 vp_p.n17740 vp_p.n17739 0.007
R20269 vp_p.n17745 vp_p.n17744 0.007
R20270 vp_p.n9207 vp_p.n9206 0.007
R20271 vp_p.n9212 vp_p.n9211 0.007
R20272 vp_p.n16313 vp_p.n16312 0.007
R20273 vp_p.n16318 vp_p.n16317 0.007
R20274 vp_p.n10644 vp_p.n10643 0.007
R20275 vp_p.n10649 vp_p.n10648 0.007
R20276 vp_p.n14885 vp_p.n14884 0.007
R20277 vp_p.n14890 vp_p.n14889 0.007
R20278 vp_p.n12082 vp_p.n12081 0.007
R20279 vp_p.n12087 vp_p.n12086 0.007
R20280 vp_p.n13846 vp_p.n13845 0.007
R20281 vp_p.n13851 vp_p.n13850 0.007
R20282 vp_p.n14390 vp_p.n14389 0.007
R20283 vp_p.n14395 vp_p.n14394 0.007
R20284 vp_p.n14400 vp_p.n14399 0.007
R20285 vp_p.n14405 vp_p.n14404 0.007
R20286 vp_p.n14410 vp_p.n14409 0.007
R20287 vp_p.n14415 vp_p.n14414 0.007
R20288 vp_p.n14420 vp_p.n14419 0.007
R20289 vp_p.n14425 vp_p.n14424 0.007
R20290 vp_p.n14430 vp_p.n14429 0.007
R20291 vp_p.n14435 vp_p.n14434 0.007
R20292 vp_p.n14440 vp_p.n14439 0.007
R20293 vp_p.n14445 vp_p.n14444 0.007
R20294 vp_p.n14450 vp_p.n14449 0.007
R20295 vp_p.n14455 vp_p.n14454 0.007
R20296 vp_p.n14460 vp_p.n14459 0.007
R20297 vp_p.n14465 vp_p.n14464 0.007
R20298 vp_p.n14385 vp_p.n14384 0.007
R20299 vp_p.n13026 vp_p.n13025 0.007
R20300 vp_p.n13031 vp_p.n13030 0.007
R20301 vp_p.n13036 vp_p.n13035 0.007
R20302 vp_p.n13041 vp_p.n13040 0.007
R20303 vp_p.n13046 vp_p.n13045 0.007
R20304 vp_p.n13051 vp_p.n13050 0.007
R20305 vp_p.n13056 vp_p.n13055 0.007
R20306 vp_p.n13061 vp_p.n13060 0.007
R20307 vp_p.n13066 vp_p.n13065 0.007
R20308 vp_p.n13071 vp_p.n13070 0.007
R20309 vp_p.n13076 vp_p.n13075 0.007
R20310 vp_p.n13081 vp_p.n13080 0.007
R20311 vp_p.n13086 vp_p.n13085 0.007
R20312 vp_p.n13091 vp_p.n13090 0.007
R20313 vp_p.n13096 vp_p.n13095 0.007
R20314 vp_p.n13021 vp_p.n13020 0.007
R20315 vp_p.n15833 vp_p.n15832 0.007
R20316 vp_p.n15838 vp_p.n15837 0.007
R20317 vp_p.n15843 vp_p.n15842 0.007
R20318 vp_p.n15848 vp_p.n15847 0.007
R20319 vp_p.n15853 vp_p.n15852 0.007
R20320 vp_p.n15858 vp_p.n15857 0.007
R20321 vp_p.n15863 vp_p.n15862 0.007
R20322 vp_p.n15868 vp_p.n15867 0.007
R20323 vp_p.n15873 vp_p.n15872 0.007
R20324 vp_p.n15878 vp_p.n15877 0.007
R20325 vp_p.n15883 vp_p.n15882 0.007
R20326 vp_p.n15888 vp_p.n15887 0.007
R20327 vp_p.n15893 vp_p.n15892 0.007
R20328 vp_p.n15898 vp_p.n15897 0.007
R20329 vp_p.n15828 vp_p.n15827 0.007
R20330 vp_p.n11602 vp_p.n11601 0.007
R20331 vp_p.n11607 vp_p.n11606 0.007
R20332 vp_p.n11612 vp_p.n11611 0.007
R20333 vp_p.n11617 vp_p.n11616 0.007
R20334 vp_p.n11622 vp_p.n11621 0.007
R20335 vp_p.n11627 vp_p.n11626 0.007
R20336 vp_p.n11632 vp_p.n11631 0.007
R20337 vp_p.n11637 vp_p.n11636 0.007
R20338 vp_p.n11642 vp_p.n11641 0.007
R20339 vp_p.n11647 vp_p.n11646 0.007
R20340 vp_p.n11652 vp_p.n11651 0.007
R20341 vp_p.n11657 vp_p.n11656 0.007
R20342 vp_p.n11662 vp_p.n11661 0.007
R20343 vp_p.n11597 vp_p.n11596 0.007
R20344 vp_p.n17275 vp_p.n17274 0.007
R20345 vp_p.n17280 vp_p.n17279 0.007
R20346 vp_p.n17285 vp_p.n17284 0.007
R20347 vp_p.n17290 vp_p.n17289 0.007
R20348 vp_p.n17295 vp_p.n17294 0.007
R20349 vp_p.n17300 vp_p.n17299 0.007
R20350 vp_p.n17305 vp_p.n17304 0.007
R20351 vp_p.n17310 vp_p.n17309 0.007
R20352 vp_p.n17315 vp_p.n17314 0.007
R20353 vp_p.n17320 vp_p.n17319 0.007
R20354 vp_p.n17325 vp_p.n17324 0.007
R20355 vp_p.n17330 vp_p.n17329 0.007
R20356 vp_p.n17270 vp_p.n17269 0.007
R20357 vp_p.n10179 vp_p.n10178 0.007
R20358 vp_p.n10184 vp_p.n10183 0.007
R20359 vp_p.n10189 vp_p.n10188 0.007
R20360 vp_p.n10194 vp_p.n10193 0.007
R20361 vp_p.n10199 vp_p.n10198 0.007
R20362 vp_p.n10204 vp_p.n10203 0.007
R20363 vp_p.n10209 vp_p.n10208 0.007
R20364 vp_p.n10214 vp_p.n10213 0.007
R20365 vp_p.n10219 vp_p.n10218 0.007
R20366 vp_p.n10224 vp_p.n10223 0.007
R20367 vp_p.n10229 vp_p.n10228 0.007
R20368 vp_p.n10174 vp_p.n10173 0.007
R20369 vp_p.n18716 vp_p.n18715 0.007
R20370 vp_p.n18721 vp_p.n18720 0.007
R20371 vp_p.n18726 vp_p.n18725 0.007
R20372 vp_p.n18731 vp_p.n18730 0.007
R20373 vp_p.n18736 vp_p.n18735 0.007
R20374 vp_p.n18741 vp_p.n18740 0.007
R20375 vp_p.n18746 vp_p.n18745 0.007
R20376 vp_p.n18751 vp_p.n18750 0.007
R20377 vp_p.n18756 vp_p.n18755 0.007
R20378 vp_p.n18761 vp_p.n18760 0.007
R20379 vp_p.n18711 vp_p.n18710 0.007
R20380 vp_p.n1447 vp_p.n1446 0.007
R20381 vp_p.n1452 vp_p.n1451 0.007
R20382 vp_p.n1457 vp_p.n1456 0.007
R20383 vp_p.n1462 vp_p.n1461 0.007
R20384 vp_p.n1467 vp_p.n1466 0.007
R20385 vp_p.n1472 vp_p.n1471 0.007
R20386 vp_p.n1477 vp_p.n1476 0.007
R20387 vp_p.n1482 vp_p.n1481 0.007
R20388 vp_p.n1487 vp_p.n1486 0.007
R20389 vp_p.n1442 vp_p.n1441 0.007
R20390 vp_p.n20156 vp_p.n20155 0.007
R20391 vp_p.n20161 vp_p.n20160 0.007
R20392 vp_p.n20166 vp_p.n20165 0.007
R20393 vp_p.n20171 vp_p.n20170 0.007
R20394 vp_p.n20176 vp_p.n20175 0.007
R20395 vp_p.n20181 vp_p.n20180 0.007
R20396 vp_p.n20186 vp_p.n20185 0.007
R20397 vp_p.n20191 vp_p.n20190 0.007
R20398 vp_p.n20151 vp_p.n20150 0.007
R20399 vp_p.n2887 vp_p.n2886 0.007
R20400 vp_p.n2892 vp_p.n2891 0.007
R20401 vp_p.n2897 vp_p.n2896 0.007
R20402 vp_p.n2902 vp_p.n2901 0.007
R20403 vp_p.n2907 vp_p.n2906 0.007
R20404 vp_p.n2912 vp_p.n2911 0.007
R20405 vp_p.n2917 vp_p.n2916 0.007
R20406 vp_p.n2882 vp_p.n2881 0.007
R20407 vp_p.n21595 vp_p.n21594 0.007
R20408 vp_p.n21600 vp_p.n21599 0.007
R20409 vp_p.n21605 vp_p.n21604 0.007
R20410 vp_p.n21610 vp_p.n21609 0.007
R20411 vp_p.n21615 vp_p.n21614 0.007
R20412 vp_p.n21620 vp_p.n21619 0.007
R20413 vp_p.n21590 vp_p.n21589 0.007
R20414 vp_p.n4326 vp_p.n4325 0.007
R20415 vp_p.n4331 vp_p.n4330 0.007
R20416 vp_p.n4336 vp_p.n4335 0.007
R20417 vp_p.n4341 vp_p.n4340 0.007
R20418 vp_p.n4346 vp_p.n4345 0.007
R20419 vp_p.n4321 vp_p.n4320 0.007
R20420 vp_p.n23033 vp_p.n23032 0.007
R20421 vp_p.n23038 vp_p.n23037 0.007
R20422 vp_p.n23043 vp_p.n23042 0.007
R20423 vp_p.n23048 vp_p.n23047 0.007
R20424 vp_p.n23028 vp_p.n23027 0.007
R20425 vp_p.n5764 vp_p.n5763 0.007
R20426 vp_p.n5769 vp_p.n5768 0.007
R20427 vp_p.n5774 vp_p.n5773 0.007
R20428 vp_p.n5759 vp_p.n5758 0.007
R20429 vp_p.n24470 vp_p.n24469 0.007
R20430 vp_p.n24475 vp_p.n24474 0.007
R20431 vp_p.n24465 vp_p.n24464 0.007
R20432 vp_p.n7201 vp_p.n7200 0.007
R20433 vp_p.n7196 vp_p.n7195 0.007
R20434 vp_p.n25901 vp_p.n25900 0.007
R20435 vp_p.n7586 vp_p.n7585 0.007
R20436 vp_p.n8629 vp_p.n8628 0.007
R20437 vp_p.n8628 vp_p.n8627 0.007
R20438 vp_p.n26287 vp_p.n26286 0.007
R20439 vp_p.n26286 vp_p.n26285 0.007
R20440 vp_p.n13847 vp_p.n13846 0.007
R20441 vp_p.n13852 vp_p.n13851 0.007
R20442 vp_p.n14386 vp_p.n14385 0.007
R20443 vp_p.n14391 vp_p.n14390 0.007
R20444 vp_p.n14396 vp_p.n14395 0.007
R20445 vp_p.n14401 vp_p.n14400 0.007
R20446 vp_p.n14406 vp_p.n14405 0.007
R20447 vp_p.n14411 vp_p.n14410 0.007
R20448 vp_p.n14416 vp_p.n14415 0.007
R20449 vp_p.n14421 vp_p.n14420 0.007
R20450 vp_p.n14426 vp_p.n14425 0.007
R20451 vp_p.n14431 vp_p.n14430 0.007
R20452 vp_p.n14436 vp_p.n14435 0.007
R20453 vp_p.n14441 vp_p.n14440 0.007
R20454 vp_p.n14446 vp_p.n14445 0.007
R20455 vp_p.n14451 vp_p.n14450 0.007
R20456 vp_p.n14456 vp_p.n14455 0.007
R20457 vp_p.n14461 vp_p.n14460 0.007
R20458 vp_p.n14466 vp_p.n14465 0.007
R20459 vp_p.n12083 vp_p.n12082 0.007
R20460 vp_p.n12088 vp_p.n12087 0.007
R20461 vp_p.n13022 vp_p.n13021 0.007
R20462 vp_p.n13027 vp_p.n13026 0.007
R20463 vp_p.n13032 vp_p.n13031 0.007
R20464 vp_p.n13037 vp_p.n13036 0.007
R20465 vp_p.n13042 vp_p.n13041 0.007
R20466 vp_p.n13047 vp_p.n13046 0.007
R20467 vp_p.n13052 vp_p.n13051 0.007
R20468 vp_p.n13057 vp_p.n13056 0.007
R20469 vp_p.n13062 vp_p.n13061 0.007
R20470 vp_p.n13067 vp_p.n13066 0.007
R20471 vp_p.n13072 vp_p.n13071 0.007
R20472 vp_p.n13077 vp_p.n13076 0.007
R20473 vp_p.n13082 vp_p.n13081 0.007
R20474 vp_p.n13087 vp_p.n13086 0.007
R20475 vp_p.n13092 vp_p.n13091 0.007
R20476 vp_p.n13097 vp_p.n13096 0.007
R20477 vp_p.n14886 vp_p.n14885 0.007
R20478 vp_p.n14891 vp_p.n14890 0.007
R20479 vp_p.n15829 vp_p.n15828 0.007
R20480 vp_p.n15834 vp_p.n15833 0.007
R20481 vp_p.n15839 vp_p.n15838 0.007
R20482 vp_p.n15844 vp_p.n15843 0.007
R20483 vp_p.n15849 vp_p.n15848 0.007
R20484 vp_p.n15854 vp_p.n15853 0.007
R20485 vp_p.n15859 vp_p.n15858 0.007
R20486 vp_p.n15864 vp_p.n15863 0.007
R20487 vp_p.n15869 vp_p.n15868 0.007
R20488 vp_p.n15874 vp_p.n15873 0.007
R20489 vp_p.n15879 vp_p.n15878 0.007
R20490 vp_p.n15884 vp_p.n15883 0.007
R20491 vp_p.n15889 vp_p.n15888 0.007
R20492 vp_p.n15894 vp_p.n15893 0.007
R20493 vp_p.n15899 vp_p.n15898 0.007
R20494 vp_p.n10645 vp_p.n10644 0.007
R20495 vp_p.n10650 vp_p.n10649 0.007
R20496 vp_p.n11598 vp_p.n11597 0.007
R20497 vp_p.n11603 vp_p.n11602 0.007
R20498 vp_p.n11608 vp_p.n11607 0.007
R20499 vp_p.n11613 vp_p.n11612 0.007
R20500 vp_p.n11618 vp_p.n11617 0.007
R20501 vp_p.n11623 vp_p.n11622 0.007
R20502 vp_p.n11628 vp_p.n11627 0.007
R20503 vp_p.n11633 vp_p.n11632 0.007
R20504 vp_p.n11638 vp_p.n11637 0.007
R20505 vp_p.n11643 vp_p.n11642 0.007
R20506 vp_p.n11648 vp_p.n11647 0.007
R20507 vp_p.n11653 vp_p.n11652 0.007
R20508 vp_p.n11658 vp_p.n11657 0.007
R20509 vp_p.n11663 vp_p.n11662 0.007
R20510 vp_p.n16314 vp_p.n16313 0.007
R20511 vp_p.n16319 vp_p.n16318 0.007
R20512 vp_p.n17271 vp_p.n17270 0.007
R20513 vp_p.n17276 vp_p.n17275 0.007
R20514 vp_p.n17281 vp_p.n17280 0.007
R20515 vp_p.n17286 vp_p.n17285 0.007
R20516 vp_p.n17291 vp_p.n17290 0.007
R20517 vp_p.n17296 vp_p.n17295 0.007
R20518 vp_p.n17301 vp_p.n17300 0.007
R20519 vp_p.n17306 vp_p.n17305 0.007
R20520 vp_p.n17311 vp_p.n17310 0.007
R20521 vp_p.n17316 vp_p.n17315 0.007
R20522 vp_p.n17321 vp_p.n17320 0.007
R20523 vp_p.n17326 vp_p.n17325 0.007
R20524 vp_p.n17331 vp_p.n17330 0.007
R20525 vp_p.n9208 vp_p.n9207 0.007
R20526 vp_p.n9213 vp_p.n9212 0.007
R20527 vp_p.n10175 vp_p.n10174 0.007
R20528 vp_p.n10180 vp_p.n10179 0.007
R20529 vp_p.n10185 vp_p.n10184 0.007
R20530 vp_p.n10190 vp_p.n10189 0.007
R20531 vp_p.n10195 vp_p.n10194 0.007
R20532 vp_p.n10200 vp_p.n10199 0.007
R20533 vp_p.n10205 vp_p.n10204 0.007
R20534 vp_p.n10210 vp_p.n10209 0.007
R20535 vp_p.n10215 vp_p.n10214 0.007
R20536 vp_p.n10220 vp_p.n10219 0.007
R20537 vp_p.n10225 vp_p.n10224 0.007
R20538 vp_p.n10230 vp_p.n10229 0.007
R20539 vp_p.n17741 vp_p.n17740 0.007
R20540 vp_p.n17746 vp_p.n17745 0.007
R20541 vp_p.n18712 vp_p.n18711 0.007
R20542 vp_p.n18717 vp_p.n18716 0.007
R20543 vp_p.n18722 vp_p.n18721 0.007
R20544 vp_p.n18727 vp_p.n18726 0.007
R20545 vp_p.n18732 vp_p.n18731 0.007
R20546 vp_p.n18737 vp_p.n18736 0.007
R20547 vp_p.n18742 vp_p.n18741 0.007
R20548 vp_p.n18747 vp_p.n18746 0.007
R20549 vp_p.n18752 vp_p.n18751 0.007
R20550 vp_p.n18757 vp_p.n18756 0.007
R20551 vp_p.n18762 vp_p.n18761 0.007
R20552 vp_p.n462 vp_p.n461 0.007
R20553 vp_p.n467 vp_p.n466 0.007
R20554 vp_p.n1443 vp_p.n1442 0.007
R20555 vp_p.n1448 vp_p.n1447 0.007
R20556 vp_p.n1453 vp_p.n1452 0.007
R20557 vp_p.n1458 vp_p.n1457 0.007
R20558 vp_p.n1463 vp_p.n1462 0.007
R20559 vp_p.n1468 vp_p.n1467 0.007
R20560 vp_p.n1473 vp_p.n1472 0.007
R20561 vp_p.n1478 vp_p.n1477 0.007
R20562 vp_p.n1483 vp_p.n1482 0.007
R20563 vp_p.n1488 vp_p.n1487 0.007
R20564 vp_p.n19167 vp_p.n19166 0.007
R20565 vp_p.n19172 vp_p.n19171 0.007
R20566 vp_p.n20152 vp_p.n20151 0.007
R20567 vp_p.n20157 vp_p.n20156 0.007
R20568 vp_p.n20162 vp_p.n20161 0.007
R20569 vp_p.n20167 vp_p.n20166 0.007
R20570 vp_p.n20172 vp_p.n20171 0.007
R20571 vp_p.n20177 vp_p.n20176 0.007
R20572 vp_p.n20182 vp_p.n20181 0.007
R20573 vp_p.n20187 vp_p.n20186 0.007
R20574 vp_p.n20192 vp_p.n20191 0.007
R20575 vp_p.n1888 vp_p.n1887 0.007
R20576 vp_p.n1893 vp_p.n1892 0.007
R20577 vp_p.n2883 vp_p.n2882 0.007
R20578 vp_p.n2888 vp_p.n2887 0.007
R20579 vp_p.n2893 vp_p.n2892 0.007
R20580 vp_p.n2898 vp_p.n2897 0.007
R20581 vp_p.n2903 vp_p.n2902 0.007
R20582 vp_p.n2908 vp_p.n2907 0.007
R20583 vp_p.n2913 vp_p.n2912 0.007
R20584 vp_p.n2918 vp_p.n2917 0.007
R20585 vp_p.n20592 vp_p.n20591 0.007
R20586 vp_p.n20597 vp_p.n20596 0.007
R20587 vp_p.n21591 vp_p.n21590 0.007
R20588 vp_p.n21596 vp_p.n21595 0.007
R20589 vp_p.n21601 vp_p.n21600 0.007
R20590 vp_p.n21606 vp_p.n21605 0.007
R20591 vp_p.n21611 vp_p.n21610 0.007
R20592 vp_p.n21616 vp_p.n21615 0.007
R20593 vp_p.n21621 vp_p.n21620 0.007
R20594 vp_p.n3313 vp_p.n3312 0.007
R20595 vp_p.n3318 vp_p.n3317 0.007
R20596 vp_p.n4322 vp_p.n4321 0.007
R20597 vp_p.n4327 vp_p.n4326 0.007
R20598 vp_p.n4332 vp_p.n4331 0.007
R20599 vp_p.n4337 vp_p.n4336 0.007
R20600 vp_p.n4342 vp_p.n4341 0.007
R20601 vp_p.n4347 vp_p.n4346 0.007
R20602 vp_p.n22016 vp_p.n22015 0.007
R20603 vp_p.n22021 vp_p.n22020 0.007
R20604 vp_p.n23029 vp_p.n23028 0.007
R20605 vp_p.n23034 vp_p.n23033 0.007
R20606 vp_p.n23039 vp_p.n23038 0.007
R20607 vp_p.n23044 vp_p.n23043 0.007
R20608 vp_p.n23049 vp_p.n23048 0.007
R20609 vp_p.n4737 vp_p.n4736 0.007
R20610 vp_p.n4742 vp_p.n4741 0.007
R20611 vp_p.n5760 vp_p.n5759 0.007
R20612 vp_p.n5765 vp_p.n5764 0.007
R20613 vp_p.n5770 vp_p.n5769 0.007
R20614 vp_p.n5775 vp_p.n5774 0.007
R20615 vp_p.n23439 vp_p.n23438 0.007
R20616 vp_p.n23444 vp_p.n23443 0.007
R20617 vp_p.n24466 vp_p.n24465 0.007
R20618 vp_p.n24471 vp_p.n24470 0.007
R20619 vp_p.n24476 vp_p.n24475 0.007
R20620 vp_p.n6160 vp_p.n6159 0.007
R20621 vp_p.n6165 vp_p.n6164 0.007
R20622 vp_p.n7197 vp_p.n7196 0.007
R20623 vp_p.n7202 vp_p.n7201 0.007
R20624 vp_p.n24861 vp_p.n24860 0.007
R20625 vp_p.n24866 vp_p.n24865 0.007
R20626 vp_p.n25902 vp_p.n25901 0.007
R20627 vp_p.n7577 vp_p.n7576 0.007
R20628 vp_p.n7587 vp_p.n7586 0.007
R20629 vp_p.n8627 vp_p.n8621 0.007
R20630 vp_p.n13844 vp_p.n13843 0.006
R20631 vp_p.n13849 vp_p.n13848 0.006
R20632 vp_p.n13854 vp_p.n13853 0.006
R20633 vp_p.n13858 vp_p.n13857 0.006
R20634 vp_p.n13862 vp_p.n13861 0.006
R20635 vp_p.n13866 vp_p.n13865 0.006
R20636 vp_p.n13870 vp_p.n13869 0.006
R20637 vp_p.n13874 vp_p.n13873 0.006
R20638 vp_p.n13878 vp_p.n13877 0.006
R20639 vp_p.n13882 vp_p.n13881 0.006
R20640 vp_p.n13886 vp_p.n13885 0.006
R20641 vp_p.n13890 vp_p.n13889 0.006
R20642 vp_p.n13894 vp_p.n13893 0.006
R20643 vp_p.n13898 vp_p.n13897 0.006
R20644 vp_p.n13902 vp_p.n13901 0.006
R20645 vp_p.n13906 vp_p.n13905 0.006
R20646 vp_p.n13910 vp_p.n13909 0.006
R20647 vp_p.n13914 vp_p.n13913 0.006
R20648 vp_p.n13918 vp_p.n13917 0.006
R20649 vp_p.n13922 vp_p.n13921 0.006
R20650 vp_p.n13926 vp_p.n13925 0.006
R20651 vp_p.n13930 vp_p.n13929 0.006
R20652 vp_p.n13934 vp_p.n13933 0.006
R20653 vp_p.n13938 vp_p.n13937 0.006
R20654 vp_p.n13942 vp_p.n13941 0.006
R20655 vp_p.n13946 vp_p.n13945 0.006
R20656 vp_p.n13950 vp_p.n13949 0.006
R20657 vp_p.n13954 vp_p.n13953 0.006
R20658 vp_p.n13958 vp_p.n13957 0.006
R20659 vp_p.n13962 vp_p.n13961 0.006
R20660 vp_p.n13966 vp_p.n13965 0.006
R20661 vp_p.n13970 vp_p.n13969 0.006
R20662 vp_p.n13974 vp_p.n13973 0.006
R20663 vp_p.n13978 vp_p.n13977 0.006
R20664 vp_p.n13982 vp_p.n13981 0.006
R20665 vp_p.n13986 vp_p.n13985 0.006
R20666 vp_p.n13990 vp_p.n13989 0.006
R20667 vp_p.n13994 vp_p.n13993 0.006
R20668 vp_p.n13998 vp_p.n13997 0.006
R20669 vp_p.n14002 vp_p.n14001 0.006
R20670 vp_p.n14006 vp_p.n14005 0.006
R20671 vp_p.n14010 vp_p.n14009 0.006
R20672 vp_p.n14014 vp_p.n14013 0.006
R20673 vp_p.n14018 vp_p.n14017 0.006
R20674 vp_p.n14022 vp_p.n14021 0.006
R20675 vp_p.n14026 vp_p.n14025 0.006
R20676 vp_p.n14030 vp_p.n14029 0.006
R20677 vp_p.n14034 vp_p.n14033 0.006
R20678 vp_p.n14038 vp_p.n14037 0.006
R20679 vp_p.n14042 vp_p.n14041 0.006
R20680 vp_p.n14046 vp_p.n14045 0.006
R20681 vp_p.n14050 vp_p.n14049 0.006
R20682 vp_p.n14054 vp_p.n14053 0.006
R20683 vp_p.n14058 vp_p.n14057 0.006
R20684 vp_p.n14062 vp_p.n14061 0.006
R20685 vp_p.n14066 vp_p.n14065 0.006
R20686 vp_p.n14070 vp_p.n14069 0.006
R20687 vp_p.n14074 vp_p.n14073 0.006
R20688 vp_p.n14078 vp_p.n14077 0.006
R20689 vp_p.n14082 vp_p.n14081 0.006
R20690 vp_p.n14086 vp_p.n14085 0.006
R20691 vp_p.n14090 vp_p.n14089 0.006
R20692 vp_p.n14094 vp_p.n14093 0.006
R20693 vp_p.n14098 vp_p.n14097 0.006
R20694 vp_p.n14102 vp_p.n14101 0.006
R20695 vp_p.n14106 vp_p.n14105 0.006
R20696 vp_p.n14110 vp_p.n14109 0.006
R20697 vp_p.n14114 vp_p.n14113 0.006
R20698 vp_p.n14118 vp_p.n14117 0.006
R20699 vp_p.n14122 vp_p.n14121 0.006
R20700 vp_p.n14126 vp_p.n14125 0.006
R20701 vp_p.n14130 vp_p.n14129 0.006
R20702 vp_p.n14134 vp_p.n14133 0.006
R20703 vp_p.n14138 vp_p.n14137 0.006
R20704 vp_p.n14142 vp_p.n14141 0.006
R20705 vp_p.n14146 vp_p.n14145 0.006
R20706 vp_p.n14150 vp_p.n14149 0.006
R20707 vp_p.n14154 vp_p.n14153 0.006
R20708 vp_p.n14158 vp_p.n14157 0.006
R20709 vp_p.n14162 vp_p.n14161 0.006
R20710 vp_p.n14166 vp_p.n14165 0.006
R20711 vp_p.n14170 vp_p.n14169 0.006
R20712 vp_p.n14174 vp_p.n14173 0.006
R20713 vp_p.n14178 vp_p.n14177 0.006
R20714 vp_p.n14182 vp_p.n14181 0.006
R20715 vp_p.n14186 vp_p.n14185 0.006
R20716 vp_p.n14190 vp_p.n14189 0.006
R20717 vp_p.n14194 vp_p.n14193 0.006
R20718 vp_p.n14198 vp_p.n14197 0.006
R20719 vp_p.n14202 vp_p.n14201 0.006
R20720 vp_p.n14206 vp_p.n14205 0.006
R20721 vp_p.n14210 vp_p.n14209 0.006
R20722 vp_p.n14214 vp_p.n14213 0.006
R20723 vp_p.n14218 vp_p.n14217 0.006
R20724 vp_p.n14222 vp_p.n14221 0.006
R20725 vp_p.n14226 vp_p.n14225 0.006
R20726 vp_p.n14230 vp_p.n14229 0.006
R20727 vp_p.n14234 vp_p.n14233 0.006
R20728 vp_p.n14238 vp_p.n14237 0.006
R20729 vp_p.n14242 vp_p.n14241 0.006
R20730 vp_p.n14246 vp_p.n14245 0.006
R20731 vp_p.n14250 vp_p.n14249 0.006
R20732 vp_p.n14254 vp_p.n14253 0.006
R20733 vp_p.n14258 vp_p.n14257 0.006
R20734 vp_p.n14262 vp_p.n14261 0.006
R20735 vp_p.n14266 vp_p.n14265 0.006
R20736 vp_p.n14270 vp_p.n14269 0.006
R20737 vp_p.n14274 vp_p.n14273 0.006
R20738 vp_p.n14278 vp_p.n14277 0.006
R20739 vp_p.n14282 vp_p.n14281 0.006
R20740 vp_p.n14286 vp_p.n14285 0.006
R20741 vp_p.n14290 vp_p.n14289 0.006
R20742 vp_p.n14294 vp_p.n14293 0.006
R20743 vp_p.n14298 vp_p.n14297 0.006
R20744 vp_p.n14302 vp_p.n14301 0.006
R20745 vp_p.n14306 vp_p.n14305 0.006
R20746 vp_p.n14310 vp_p.n14309 0.006
R20747 vp_p.n14314 vp_p.n14313 0.006
R20748 vp_p.n14318 vp_p.n14317 0.006
R20749 vp_p.n14322 vp_p.n14321 0.006
R20750 vp_p.n14326 vp_p.n14325 0.006
R20751 vp_p.n14330 vp_p.n14329 0.006
R20752 vp_p.n14334 vp_p.n14333 0.006
R20753 vp_p.n14338 vp_p.n14337 0.006
R20754 vp_p.n14342 vp_p.n14341 0.006
R20755 vp_p.n14346 vp_p.n14345 0.006
R20756 vp_p.n14350 vp_p.n14349 0.006
R20757 vp_p.n14354 vp_p.n14353 0.006
R20758 vp_p.n14358 vp_p.n14357 0.006
R20759 vp_p.n14362 vp_p.n14361 0.006
R20760 vp_p.n14366 vp_p.n14365 0.006
R20761 vp_p.n14370 vp_p.n14369 0.006
R20762 vp_p.n14374 vp_p.n14373 0.006
R20763 vp_p.n14384 vp_p.n14378 0.006
R20764 vp_p.n14388 vp_p.n14387 0.006
R20765 vp_p.n14393 vp_p.n14392 0.006
R20766 vp_p.n14398 vp_p.n14397 0.006
R20767 vp_p.n14403 vp_p.n14402 0.006
R20768 vp_p.n14408 vp_p.n14407 0.006
R20769 vp_p.n14413 vp_p.n14412 0.006
R20770 vp_p.n14418 vp_p.n14417 0.006
R20771 vp_p.n14423 vp_p.n14422 0.006
R20772 vp_p.n14428 vp_p.n14427 0.006
R20773 vp_p.n14433 vp_p.n14432 0.006
R20774 vp_p.n14438 vp_p.n14437 0.006
R20775 vp_p.n14443 vp_p.n14442 0.006
R20776 vp_p.n14448 vp_p.n14447 0.006
R20777 vp_p.n14453 vp_p.n14452 0.006
R20778 vp_p.n14458 vp_p.n14457 0.006
R20779 vp_p.n14463 vp_p.n14462 0.006
R20780 vp_p.n14375 vp_p.n14374 0.006
R20781 vp_p.n14371 vp_p.n14370 0.006
R20782 vp_p.n14367 vp_p.n14366 0.006
R20783 vp_p.n14363 vp_p.n14362 0.006
R20784 vp_p.n14359 vp_p.n14358 0.006
R20785 vp_p.n14355 vp_p.n14354 0.006
R20786 vp_p.n14351 vp_p.n14350 0.006
R20787 vp_p.n14347 vp_p.n14346 0.006
R20788 vp_p.n14343 vp_p.n14342 0.006
R20789 vp_p.n14339 vp_p.n14338 0.006
R20790 vp_p.n14335 vp_p.n14334 0.006
R20791 vp_p.n14331 vp_p.n14330 0.006
R20792 vp_p.n14327 vp_p.n14326 0.006
R20793 vp_p.n14323 vp_p.n14322 0.006
R20794 vp_p.n14319 vp_p.n14318 0.006
R20795 vp_p.n14315 vp_p.n14314 0.006
R20796 vp_p.n14311 vp_p.n14310 0.006
R20797 vp_p.n14307 vp_p.n14306 0.006
R20798 vp_p.n14303 vp_p.n14302 0.006
R20799 vp_p.n14299 vp_p.n14298 0.006
R20800 vp_p.n14295 vp_p.n14294 0.006
R20801 vp_p.n14291 vp_p.n14290 0.006
R20802 vp_p.n14287 vp_p.n14286 0.006
R20803 vp_p.n14283 vp_p.n14282 0.006
R20804 vp_p.n14279 vp_p.n14278 0.006
R20805 vp_p.n14275 vp_p.n14274 0.006
R20806 vp_p.n14271 vp_p.n14270 0.006
R20807 vp_p.n14267 vp_p.n14266 0.006
R20808 vp_p.n14263 vp_p.n14262 0.006
R20809 vp_p.n14259 vp_p.n14258 0.006
R20810 vp_p.n14255 vp_p.n14254 0.006
R20811 vp_p.n14251 vp_p.n14250 0.006
R20812 vp_p.n14247 vp_p.n14246 0.006
R20813 vp_p.n14243 vp_p.n14242 0.006
R20814 vp_p.n14239 vp_p.n14238 0.006
R20815 vp_p.n14235 vp_p.n14234 0.006
R20816 vp_p.n14231 vp_p.n14230 0.006
R20817 vp_p.n14227 vp_p.n14226 0.006
R20818 vp_p.n14223 vp_p.n14222 0.006
R20819 vp_p.n14219 vp_p.n14218 0.006
R20820 vp_p.n14215 vp_p.n14214 0.006
R20821 vp_p.n14211 vp_p.n14210 0.006
R20822 vp_p.n14207 vp_p.n14206 0.006
R20823 vp_p.n14203 vp_p.n14202 0.006
R20824 vp_p.n14199 vp_p.n14198 0.006
R20825 vp_p.n14195 vp_p.n14194 0.006
R20826 vp_p.n14191 vp_p.n14190 0.006
R20827 vp_p.n14187 vp_p.n14186 0.006
R20828 vp_p.n14183 vp_p.n14182 0.006
R20829 vp_p.n14179 vp_p.n14178 0.006
R20830 vp_p.n14175 vp_p.n14174 0.006
R20831 vp_p.n14171 vp_p.n14170 0.006
R20832 vp_p.n14167 vp_p.n14166 0.006
R20833 vp_p.n14163 vp_p.n14162 0.006
R20834 vp_p.n14159 vp_p.n14158 0.006
R20835 vp_p.n14155 vp_p.n14154 0.006
R20836 vp_p.n14151 vp_p.n14150 0.006
R20837 vp_p.n14147 vp_p.n14146 0.006
R20838 vp_p.n14143 vp_p.n14142 0.006
R20839 vp_p.n14139 vp_p.n14138 0.006
R20840 vp_p.n14135 vp_p.n14134 0.006
R20841 vp_p.n14131 vp_p.n14130 0.006
R20842 vp_p.n14127 vp_p.n14126 0.006
R20843 vp_p.n14123 vp_p.n14122 0.006
R20844 vp_p.n14119 vp_p.n14118 0.006
R20845 vp_p.n14115 vp_p.n14114 0.006
R20846 vp_p.n14111 vp_p.n14110 0.006
R20847 vp_p.n14107 vp_p.n14106 0.006
R20848 vp_p.n14103 vp_p.n14102 0.006
R20849 vp_p.n14099 vp_p.n14098 0.006
R20850 vp_p.n14095 vp_p.n14094 0.006
R20851 vp_p.n14091 vp_p.n14090 0.006
R20852 vp_p.n14087 vp_p.n14086 0.006
R20853 vp_p.n14083 vp_p.n14082 0.006
R20854 vp_p.n14079 vp_p.n14078 0.006
R20855 vp_p.n14075 vp_p.n14074 0.006
R20856 vp_p.n14071 vp_p.n14070 0.006
R20857 vp_p.n14067 vp_p.n14066 0.006
R20858 vp_p.n14063 vp_p.n14062 0.006
R20859 vp_p.n14059 vp_p.n14058 0.006
R20860 vp_p.n14055 vp_p.n14054 0.006
R20861 vp_p.n14051 vp_p.n14050 0.006
R20862 vp_p.n14047 vp_p.n14046 0.006
R20863 vp_p.n14043 vp_p.n14042 0.006
R20864 vp_p.n14039 vp_p.n14038 0.006
R20865 vp_p.n14035 vp_p.n14034 0.006
R20866 vp_p.n14031 vp_p.n14030 0.006
R20867 vp_p.n14027 vp_p.n14026 0.006
R20868 vp_p.n14023 vp_p.n14022 0.006
R20869 vp_p.n14019 vp_p.n14018 0.006
R20870 vp_p.n14015 vp_p.n14014 0.006
R20871 vp_p.n14011 vp_p.n14010 0.006
R20872 vp_p.n14007 vp_p.n14006 0.006
R20873 vp_p.n14003 vp_p.n14002 0.006
R20874 vp_p.n13999 vp_p.n13998 0.006
R20875 vp_p.n13995 vp_p.n13994 0.006
R20876 vp_p.n13991 vp_p.n13990 0.006
R20877 vp_p.n13987 vp_p.n13986 0.006
R20878 vp_p.n13983 vp_p.n13982 0.006
R20879 vp_p.n13979 vp_p.n13978 0.006
R20880 vp_p.n13975 vp_p.n13974 0.006
R20881 vp_p.n13971 vp_p.n13970 0.006
R20882 vp_p.n13967 vp_p.n13966 0.006
R20883 vp_p.n13963 vp_p.n13962 0.006
R20884 vp_p.n13959 vp_p.n13958 0.006
R20885 vp_p.n13955 vp_p.n13954 0.006
R20886 vp_p.n13951 vp_p.n13950 0.006
R20887 vp_p.n13947 vp_p.n13946 0.006
R20888 vp_p.n13943 vp_p.n13942 0.006
R20889 vp_p.n13939 vp_p.n13938 0.006
R20890 vp_p.n13935 vp_p.n13934 0.006
R20891 vp_p.n13931 vp_p.n13930 0.006
R20892 vp_p.n13927 vp_p.n13926 0.006
R20893 vp_p.n13923 vp_p.n13922 0.006
R20894 vp_p.n13919 vp_p.n13918 0.006
R20895 vp_p.n13915 vp_p.n13914 0.006
R20896 vp_p.n13911 vp_p.n13910 0.006
R20897 vp_p.n13907 vp_p.n13906 0.006
R20898 vp_p.n13903 vp_p.n13902 0.006
R20899 vp_p.n13899 vp_p.n13898 0.006
R20900 vp_p.n13895 vp_p.n13894 0.006
R20901 vp_p.n13891 vp_p.n13890 0.006
R20902 vp_p.n13887 vp_p.n13886 0.006
R20903 vp_p.n13883 vp_p.n13882 0.006
R20904 vp_p.n13879 vp_p.n13878 0.006
R20905 vp_p.n13875 vp_p.n13874 0.006
R20906 vp_p.n13871 vp_p.n13870 0.006
R20907 vp_p.n13867 vp_p.n13866 0.006
R20908 vp_p.n13863 vp_p.n13862 0.006
R20909 vp_p.n13859 vp_p.n13858 0.006
R20910 vp_p.n13855 vp_p.n13854 0.006
R20911 vp_p.n14378 vp_p.n14377 0.006
R20912 vp_p.n12080 vp_p.n12079 0.006
R20913 vp_p.n12085 vp_p.n12084 0.006
R20914 vp_p.n12096 vp_p.n12090 0.006
R20915 vp_p.n12100 vp_p.n12099 0.006
R20916 vp_p.n12110 vp_p.n12104 0.006
R20917 vp_p.n12114 vp_p.n12113 0.006
R20918 vp_p.n12124 vp_p.n12118 0.006
R20919 vp_p.n12128 vp_p.n12127 0.006
R20920 vp_p.n12138 vp_p.n12132 0.006
R20921 vp_p.n12142 vp_p.n12141 0.006
R20922 vp_p.n12152 vp_p.n12146 0.006
R20923 vp_p.n12156 vp_p.n12155 0.006
R20924 vp_p.n12166 vp_p.n12160 0.006
R20925 vp_p.n12170 vp_p.n12169 0.006
R20926 vp_p.n12180 vp_p.n12174 0.006
R20927 vp_p.n12184 vp_p.n12183 0.006
R20928 vp_p.n12194 vp_p.n12188 0.006
R20929 vp_p.n12198 vp_p.n12197 0.006
R20930 vp_p.n12208 vp_p.n12202 0.006
R20931 vp_p.n12212 vp_p.n12211 0.006
R20932 vp_p.n12222 vp_p.n12216 0.006
R20933 vp_p.n12226 vp_p.n12225 0.006
R20934 vp_p.n12236 vp_p.n12230 0.006
R20935 vp_p.n12240 vp_p.n12239 0.006
R20936 vp_p.n12250 vp_p.n12244 0.006
R20937 vp_p.n12254 vp_p.n12253 0.006
R20938 vp_p.n12264 vp_p.n12258 0.006
R20939 vp_p.n12268 vp_p.n12267 0.006
R20940 vp_p.n12278 vp_p.n12272 0.006
R20941 vp_p.n12282 vp_p.n12281 0.006
R20942 vp_p.n12292 vp_p.n12286 0.006
R20943 vp_p.n12296 vp_p.n12295 0.006
R20944 vp_p.n12306 vp_p.n12300 0.006
R20945 vp_p.n12310 vp_p.n12309 0.006
R20946 vp_p.n12320 vp_p.n12314 0.006
R20947 vp_p.n12324 vp_p.n12323 0.006
R20948 vp_p.n12334 vp_p.n12328 0.006
R20949 vp_p.n12338 vp_p.n12337 0.006
R20950 vp_p.n12348 vp_p.n12342 0.006
R20951 vp_p.n12352 vp_p.n12351 0.006
R20952 vp_p.n12362 vp_p.n12356 0.006
R20953 vp_p.n12366 vp_p.n12365 0.006
R20954 vp_p.n12376 vp_p.n12370 0.006
R20955 vp_p.n12380 vp_p.n12379 0.006
R20956 vp_p.n12390 vp_p.n12384 0.006
R20957 vp_p.n12394 vp_p.n12393 0.006
R20958 vp_p.n12404 vp_p.n12398 0.006
R20959 vp_p.n12408 vp_p.n12407 0.006
R20960 vp_p.n12418 vp_p.n12412 0.006
R20961 vp_p.n12422 vp_p.n12421 0.006
R20962 vp_p.n12432 vp_p.n12426 0.006
R20963 vp_p.n12436 vp_p.n12435 0.006
R20964 vp_p.n12446 vp_p.n12440 0.006
R20965 vp_p.n12450 vp_p.n12449 0.006
R20966 vp_p.n12460 vp_p.n12454 0.006
R20967 vp_p.n12464 vp_p.n12463 0.006
R20968 vp_p.n12474 vp_p.n12468 0.006
R20969 vp_p.n12478 vp_p.n12477 0.006
R20970 vp_p.n12488 vp_p.n12482 0.006
R20971 vp_p.n12492 vp_p.n12491 0.006
R20972 vp_p.n12502 vp_p.n12496 0.006
R20973 vp_p.n12506 vp_p.n12505 0.006
R20974 vp_p.n12516 vp_p.n12510 0.006
R20975 vp_p.n12520 vp_p.n12519 0.006
R20976 vp_p.n12530 vp_p.n12524 0.006
R20977 vp_p.n12534 vp_p.n12533 0.006
R20978 vp_p.n12544 vp_p.n12538 0.006
R20979 vp_p.n12548 vp_p.n12547 0.006
R20980 vp_p.n12558 vp_p.n12552 0.006
R20981 vp_p.n12562 vp_p.n12561 0.006
R20982 vp_p.n12572 vp_p.n12566 0.006
R20983 vp_p.n12576 vp_p.n12575 0.006
R20984 vp_p.n12586 vp_p.n12580 0.006
R20985 vp_p.n12590 vp_p.n12589 0.006
R20986 vp_p.n12600 vp_p.n12594 0.006
R20987 vp_p.n12604 vp_p.n12603 0.006
R20988 vp_p.n12614 vp_p.n12608 0.006
R20989 vp_p.n12618 vp_p.n12617 0.006
R20990 vp_p.n12628 vp_p.n12622 0.006
R20991 vp_p.n12632 vp_p.n12631 0.006
R20992 vp_p.n12642 vp_p.n12636 0.006
R20993 vp_p.n12646 vp_p.n12645 0.006
R20994 vp_p.n12656 vp_p.n12650 0.006
R20995 vp_p.n12660 vp_p.n12659 0.006
R20996 vp_p.n12670 vp_p.n12664 0.006
R20997 vp_p.n12674 vp_p.n12673 0.006
R20998 vp_p.n12684 vp_p.n12678 0.006
R20999 vp_p.n12688 vp_p.n12687 0.006
R21000 vp_p.n12698 vp_p.n12692 0.006
R21001 vp_p.n12702 vp_p.n12701 0.006
R21002 vp_p.n12712 vp_p.n12706 0.006
R21003 vp_p.n12716 vp_p.n12715 0.006
R21004 vp_p.n12726 vp_p.n12720 0.006
R21005 vp_p.n12730 vp_p.n12729 0.006
R21006 vp_p.n12740 vp_p.n12734 0.006
R21007 vp_p.n12744 vp_p.n12743 0.006
R21008 vp_p.n12754 vp_p.n12748 0.006
R21009 vp_p.n12758 vp_p.n12757 0.006
R21010 vp_p.n12768 vp_p.n12762 0.006
R21011 vp_p.n12772 vp_p.n12771 0.006
R21012 vp_p.n12782 vp_p.n12776 0.006
R21013 vp_p.n12786 vp_p.n12785 0.006
R21014 vp_p.n12796 vp_p.n12790 0.006
R21015 vp_p.n12800 vp_p.n12799 0.006
R21016 vp_p.n12810 vp_p.n12804 0.006
R21017 vp_p.n12814 vp_p.n12813 0.006
R21018 vp_p.n12824 vp_p.n12818 0.006
R21019 vp_p.n12828 vp_p.n12827 0.006
R21020 vp_p.n12838 vp_p.n12832 0.006
R21021 vp_p.n12842 vp_p.n12841 0.006
R21022 vp_p.n12852 vp_p.n12846 0.006
R21023 vp_p.n12856 vp_p.n12855 0.006
R21024 vp_p.n12866 vp_p.n12860 0.006
R21025 vp_p.n12870 vp_p.n12869 0.006
R21026 vp_p.n12880 vp_p.n12874 0.006
R21027 vp_p.n12884 vp_p.n12883 0.006
R21028 vp_p.n12894 vp_p.n12888 0.006
R21029 vp_p.n12898 vp_p.n12897 0.006
R21030 vp_p.n12908 vp_p.n12902 0.006
R21031 vp_p.n12912 vp_p.n12911 0.006
R21032 vp_p.n12922 vp_p.n12916 0.006
R21033 vp_p.n12926 vp_p.n12925 0.006
R21034 vp_p.n12936 vp_p.n12930 0.006
R21035 vp_p.n12940 vp_p.n12939 0.006
R21036 vp_p.n12950 vp_p.n12944 0.006
R21037 vp_p.n12954 vp_p.n12953 0.006
R21038 vp_p.n12964 vp_p.n12958 0.006
R21039 vp_p.n12968 vp_p.n12967 0.006
R21040 vp_p.n12978 vp_p.n12972 0.006
R21041 vp_p.n12982 vp_p.n12981 0.006
R21042 vp_p.n12992 vp_p.n12986 0.006
R21043 vp_p.n12996 vp_p.n12995 0.006
R21044 vp_p.n13006 vp_p.n13000 0.006
R21045 vp_p.n13010 vp_p.n13009 0.006
R21046 vp_p.n13020 vp_p.n13014 0.006
R21047 vp_p.n13024 vp_p.n13023 0.006
R21048 vp_p.n13029 vp_p.n13028 0.006
R21049 vp_p.n13034 vp_p.n13033 0.006
R21050 vp_p.n13039 vp_p.n13038 0.006
R21051 vp_p.n13044 vp_p.n13043 0.006
R21052 vp_p.n13049 vp_p.n13048 0.006
R21053 vp_p.n13054 vp_p.n13053 0.006
R21054 vp_p.n13059 vp_p.n13058 0.006
R21055 vp_p.n13064 vp_p.n13063 0.006
R21056 vp_p.n13069 vp_p.n13068 0.006
R21057 vp_p.n13074 vp_p.n13073 0.006
R21058 vp_p.n13079 vp_p.n13078 0.006
R21059 vp_p.n13084 vp_p.n13083 0.006
R21060 vp_p.n13089 vp_p.n13088 0.006
R21061 vp_p.n13094 vp_p.n13093 0.006
R21062 vp_p.n13011 vp_p.n13010 0.006
R21063 vp_p.n13000 vp_p.n12999 0.006
R21064 vp_p.n12997 vp_p.n12996 0.006
R21065 vp_p.n12986 vp_p.n12985 0.006
R21066 vp_p.n12983 vp_p.n12982 0.006
R21067 vp_p.n12972 vp_p.n12971 0.006
R21068 vp_p.n12969 vp_p.n12968 0.006
R21069 vp_p.n12958 vp_p.n12957 0.006
R21070 vp_p.n12955 vp_p.n12954 0.006
R21071 vp_p.n12944 vp_p.n12943 0.006
R21072 vp_p.n12941 vp_p.n12940 0.006
R21073 vp_p.n12930 vp_p.n12929 0.006
R21074 vp_p.n12927 vp_p.n12926 0.006
R21075 vp_p.n12916 vp_p.n12915 0.006
R21076 vp_p.n12913 vp_p.n12912 0.006
R21077 vp_p.n12902 vp_p.n12901 0.006
R21078 vp_p.n12899 vp_p.n12898 0.006
R21079 vp_p.n12888 vp_p.n12887 0.006
R21080 vp_p.n12885 vp_p.n12884 0.006
R21081 vp_p.n12874 vp_p.n12873 0.006
R21082 vp_p.n12871 vp_p.n12870 0.006
R21083 vp_p.n12860 vp_p.n12859 0.006
R21084 vp_p.n12857 vp_p.n12856 0.006
R21085 vp_p.n12846 vp_p.n12845 0.006
R21086 vp_p.n12843 vp_p.n12842 0.006
R21087 vp_p.n12832 vp_p.n12831 0.006
R21088 vp_p.n12829 vp_p.n12828 0.006
R21089 vp_p.n12818 vp_p.n12817 0.006
R21090 vp_p.n12815 vp_p.n12814 0.006
R21091 vp_p.n12804 vp_p.n12803 0.006
R21092 vp_p.n12801 vp_p.n12800 0.006
R21093 vp_p.n12790 vp_p.n12789 0.006
R21094 vp_p.n12787 vp_p.n12786 0.006
R21095 vp_p.n12776 vp_p.n12775 0.006
R21096 vp_p.n12773 vp_p.n12772 0.006
R21097 vp_p.n12762 vp_p.n12761 0.006
R21098 vp_p.n12759 vp_p.n12758 0.006
R21099 vp_p.n12748 vp_p.n12747 0.006
R21100 vp_p.n12745 vp_p.n12744 0.006
R21101 vp_p.n12734 vp_p.n12733 0.006
R21102 vp_p.n12731 vp_p.n12730 0.006
R21103 vp_p.n12720 vp_p.n12719 0.006
R21104 vp_p.n12717 vp_p.n12716 0.006
R21105 vp_p.n12706 vp_p.n12705 0.006
R21106 vp_p.n12703 vp_p.n12702 0.006
R21107 vp_p.n12692 vp_p.n12691 0.006
R21108 vp_p.n12689 vp_p.n12688 0.006
R21109 vp_p.n12678 vp_p.n12677 0.006
R21110 vp_p.n12675 vp_p.n12674 0.006
R21111 vp_p.n12664 vp_p.n12663 0.006
R21112 vp_p.n12661 vp_p.n12660 0.006
R21113 vp_p.n12650 vp_p.n12649 0.006
R21114 vp_p.n12647 vp_p.n12646 0.006
R21115 vp_p.n12636 vp_p.n12635 0.006
R21116 vp_p.n12633 vp_p.n12632 0.006
R21117 vp_p.n12622 vp_p.n12621 0.006
R21118 vp_p.n12619 vp_p.n12618 0.006
R21119 vp_p.n12608 vp_p.n12607 0.006
R21120 vp_p.n12605 vp_p.n12604 0.006
R21121 vp_p.n12594 vp_p.n12593 0.006
R21122 vp_p.n12591 vp_p.n12590 0.006
R21123 vp_p.n12580 vp_p.n12579 0.006
R21124 vp_p.n12577 vp_p.n12576 0.006
R21125 vp_p.n12566 vp_p.n12565 0.006
R21126 vp_p.n12563 vp_p.n12562 0.006
R21127 vp_p.n12552 vp_p.n12551 0.006
R21128 vp_p.n12549 vp_p.n12548 0.006
R21129 vp_p.n12538 vp_p.n12537 0.006
R21130 vp_p.n12535 vp_p.n12534 0.006
R21131 vp_p.n12524 vp_p.n12523 0.006
R21132 vp_p.n12521 vp_p.n12520 0.006
R21133 vp_p.n12510 vp_p.n12509 0.006
R21134 vp_p.n12507 vp_p.n12506 0.006
R21135 vp_p.n12496 vp_p.n12495 0.006
R21136 vp_p.n12493 vp_p.n12492 0.006
R21137 vp_p.n12482 vp_p.n12481 0.006
R21138 vp_p.n12479 vp_p.n12478 0.006
R21139 vp_p.n12468 vp_p.n12467 0.006
R21140 vp_p.n12465 vp_p.n12464 0.006
R21141 vp_p.n12454 vp_p.n12453 0.006
R21142 vp_p.n12451 vp_p.n12450 0.006
R21143 vp_p.n12440 vp_p.n12439 0.006
R21144 vp_p.n12437 vp_p.n12436 0.006
R21145 vp_p.n12426 vp_p.n12425 0.006
R21146 vp_p.n12423 vp_p.n12422 0.006
R21147 vp_p.n12412 vp_p.n12411 0.006
R21148 vp_p.n12409 vp_p.n12408 0.006
R21149 vp_p.n12398 vp_p.n12397 0.006
R21150 vp_p.n12395 vp_p.n12394 0.006
R21151 vp_p.n12384 vp_p.n12383 0.006
R21152 vp_p.n12381 vp_p.n12380 0.006
R21153 vp_p.n12370 vp_p.n12369 0.006
R21154 vp_p.n12367 vp_p.n12366 0.006
R21155 vp_p.n12356 vp_p.n12355 0.006
R21156 vp_p.n12353 vp_p.n12352 0.006
R21157 vp_p.n12342 vp_p.n12341 0.006
R21158 vp_p.n12339 vp_p.n12338 0.006
R21159 vp_p.n12328 vp_p.n12327 0.006
R21160 vp_p.n12325 vp_p.n12324 0.006
R21161 vp_p.n12314 vp_p.n12313 0.006
R21162 vp_p.n12311 vp_p.n12310 0.006
R21163 vp_p.n12300 vp_p.n12299 0.006
R21164 vp_p.n12297 vp_p.n12296 0.006
R21165 vp_p.n12286 vp_p.n12285 0.006
R21166 vp_p.n12283 vp_p.n12282 0.006
R21167 vp_p.n12272 vp_p.n12271 0.006
R21168 vp_p.n12269 vp_p.n12268 0.006
R21169 vp_p.n12258 vp_p.n12257 0.006
R21170 vp_p.n12255 vp_p.n12254 0.006
R21171 vp_p.n12244 vp_p.n12243 0.006
R21172 vp_p.n12241 vp_p.n12240 0.006
R21173 vp_p.n12230 vp_p.n12229 0.006
R21174 vp_p.n12227 vp_p.n12226 0.006
R21175 vp_p.n12216 vp_p.n12215 0.006
R21176 vp_p.n12213 vp_p.n12212 0.006
R21177 vp_p.n12202 vp_p.n12201 0.006
R21178 vp_p.n12199 vp_p.n12198 0.006
R21179 vp_p.n12188 vp_p.n12187 0.006
R21180 vp_p.n12185 vp_p.n12184 0.006
R21181 vp_p.n12174 vp_p.n12173 0.006
R21182 vp_p.n12171 vp_p.n12170 0.006
R21183 vp_p.n12160 vp_p.n12159 0.006
R21184 vp_p.n12157 vp_p.n12156 0.006
R21185 vp_p.n12146 vp_p.n12145 0.006
R21186 vp_p.n12143 vp_p.n12142 0.006
R21187 vp_p.n12132 vp_p.n12131 0.006
R21188 vp_p.n12129 vp_p.n12128 0.006
R21189 vp_p.n12118 vp_p.n12117 0.006
R21190 vp_p.n12115 vp_p.n12114 0.006
R21191 vp_p.n12104 vp_p.n12103 0.006
R21192 vp_p.n12101 vp_p.n12100 0.006
R21193 vp_p.n12090 vp_p.n12089 0.006
R21194 vp_p.n13014 vp_p.n13013 0.006
R21195 vp_p.n14389 vp_p.n14388 0.006
R21196 vp_p.n14883 vp_p.n14882 0.006
R21197 vp_p.n14888 vp_p.n14887 0.006
R21198 vp_p.n14899 vp_p.n14893 0.006
R21199 vp_p.n14903 vp_p.n14902 0.006
R21200 vp_p.n14913 vp_p.n14907 0.006
R21201 vp_p.n14917 vp_p.n14916 0.006
R21202 vp_p.n14927 vp_p.n14921 0.006
R21203 vp_p.n14931 vp_p.n14930 0.006
R21204 vp_p.n14941 vp_p.n14935 0.006
R21205 vp_p.n14945 vp_p.n14944 0.006
R21206 vp_p.n14955 vp_p.n14949 0.006
R21207 vp_p.n14959 vp_p.n14958 0.006
R21208 vp_p.n14969 vp_p.n14963 0.006
R21209 vp_p.n14973 vp_p.n14972 0.006
R21210 vp_p.n14983 vp_p.n14977 0.006
R21211 vp_p.n14987 vp_p.n14986 0.006
R21212 vp_p.n14997 vp_p.n14991 0.006
R21213 vp_p.n15001 vp_p.n15000 0.006
R21214 vp_p.n15011 vp_p.n15005 0.006
R21215 vp_p.n15015 vp_p.n15014 0.006
R21216 vp_p.n15025 vp_p.n15019 0.006
R21217 vp_p.n15029 vp_p.n15028 0.006
R21218 vp_p.n15039 vp_p.n15033 0.006
R21219 vp_p.n15043 vp_p.n15042 0.006
R21220 vp_p.n15053 vp_p.n15047 0.006
R21221 vp_p.n15057 vp_p.n15056 0.006
R21222 vp_p.n15067 vp_p.n15061 0.006
R21223 vp_p.n15071 vp_p.n15070 0.006
R21224 vp_p.n15081 vp_p.n15075 0.006
R21225 vp_p.n15085 vp_p.n15084 0.006
R21226 vp_p.n15095 vp_p.n15089 0.006
R21227 vp_p.n15099 vp_p.n15098 0.006
R21228 vp_p.n15109 vp_p.n15103 0.006
R21229 vp_p.n15113 vp_p.n15112 0.006
R21230 vp_p.n15123 vp_p.n15117 0.006
R21231 vp_p.n15127 vp_p.n15126 0.006
R21232 vp_p.n15137 vp_p.n15131 0.006
R21233 vp_p.n15141 vp_p.n15140 0.006
R21234 vp_p.n15151 vp_p.n15145 0.006
R21235 vp_p.n15155 vp_p.n15154 0.006
R21236 vp_p.n15165 vp_p.n15159 0.006
R21237 vp_p.n15169 vp_p.n15168 0.006
R21238 vp_p.n15179 vp_p.n15173 0.006
R21239 vp_p.n15183 vp_p.n15182 0.006
R21240 vp_p.n15193 vp_p.n15187 0.006
R21241 vp_p.n15197 vp_p.n15196 0.006
R21242 vp_p.n15207 vp_p.n15201 0.006
R21243 vp_p.n15211 vp_p.n15210 0.006
R21244 vp_p.n15221 vp_p.n15215 0.006
R21245 vp_p.n15225 vp_p.n15224 0.006
R21246 vp_p.n15235 vp_p.n15229 0.006
R21247 vp_p.n15239 vp_p.n15238 0.006
R21248 vp_p.n15249 vp_p.n15243 0.006
R21249 vp_p.n15253 vp_p.n15252 0.006
R21250 vp_p.n15263 vp_p.n15257 0.006
R21251 vp_p.n15267 vp_p.n15266 0.006
R21252 vp_p.n15277 vp_p.n15271 0.006
R21253 vp_p.n15281 vp_p.n15280 0.006
R21254 vp_p.n15291 vp_p.n15285 0.006
R21255 vp_p.n15295 vp_p.n15294 0.006
R21256 vp_p.n15305 vp_p.n15299 0.006
R21257 vp_p.n15309 vp_p.n15308 0.006
R21258 vp_p.n15319 vp_p.n15313 0.006
R21259 vp_p.n15323 vp_p.n15322 0.006
R21260 vp_p.n15333 vp_p.n15327 0.006
R21261 vp_p.n15337 vp_p.n15336 0.006
R21262 vp_p.n15347 vp_p.n15341 0.006
R21263 vp_p.n15351 vp_p.n15350 0.006
R21264 vp_p.n15361 vp_p.n15355 0.006
R21265 vp_p.n15365 vp_p.n15364 0.006
R21266 vp_p.n15375 vp_p.n15369 0.006
R21267 vp_p.n15379 vp_p.n15378 0.006
R21268 vp_p.n15389 vp_p.n15383 0.006
R21269 vp_p.n15393 vp_p.n15392 0.006
R21270 vp_p.n15403 vp_p.n15397 0.006
R21271 vp_p.n15407 vp_p.n15406 0.006
R21272 vp_p.n15417 vp_p.n15411 0.006
R21273 vp_p.n15421 vp_p.n15420 0.006
R21274 vp_p.n15431 vp_p.n15425 0.006
R21275 vp_p.n15435 vp_p.n15434 0.006
R21276 vp_p.n15445 vp_p.n15439 0.006
R21277 vp_p.n15449 vp_p.n15448 0.006
R21278 vp_p.n15459 vp_p.n15453 0.006
R21279 vp_p.n15463 vp_p.n15462 0.006
R21280 vp_p.n15473 vp_p.n15467 0.006
R21281 vp_p.n15477 vp_p.n15476 0.006
R21282 vp_p.n15487 vp_p.n15481 0.006
R21283 vp_p.n15491 vp_p.n15490 0.006
R21284 vp_p.n15501 vp_p.n15495 0.006
R21285 vp_p.n15505 vp_p.n15504 0.006
R21286 vp_p.n15515 vp_p.n15509 0.006
R21287 vp_p.n15519 vp_p.n15518 0.006
R21288 vp_p.n15529 vp_p.n15523 0.006
R21289 vp_p.n15533 vp_p.n15532 0.006
R21290 vp_p.n15543 vp_p.n15537 0.006
R21291 vp_p.n15547 vp_p.n15546 0.006
R21292 vp_p.n15557 vp_p.n15551 0.006
R21293 vp_p.n15561 vp_p.n15560 0.006
R21294 vp_p.n15571 vp_p.n15565 0.006
R21295 vp_p.n15575 vp_p.n15574 0.006
R21296 vp_p.n15585 vp_p.n15579 0.006
R21297 vp_p.n15589 vp_p.n15588 0.006
R21298 vp_p.n15599 vp_p.n15593 0.006
R21299 vp_p.n15603 vp_p.n15602 0.006
R21300 vp_p.n15613 vp_p.n15607 0.006
R21301 vp_p.n15617 vp_p.n15616 0.006
R21302 vp_p.n15627 vp_p.n15621 0.006
R21303 vp_p.n15631 vp_p.n15630 0.006
R21304 vp_p.n15641 vp_p.n15635 0.006
R21305 vp_p.n15645 vp_p.n15644 0.006
R21306 vp_p.n15655 vp_p.n15649 0.006
R21307 vp_p.n15659 vp_p.n15658 0.006
R21308 vp_p.n15669 vp_p.n15663 0.006
R21309 vp_p.n15673 vp_p.n15672 0.006
R21310 vp_p.n15683 vp_p.n15677 0.006
R21311 vp_p.n15687 vp_p.n15686 0.006
R21312 vp_p.n15697 vp_p.n15691 0.006
R21313 vp_p.n15701 vp_p.n15700 0.006
R21314 vp_p.n15711 vp_p.n15705 0.006
R21315 vp_p.n15715 vp_p.n15714 0.006
R21316 vp_p.n15725 vp_p.n15719 0.006
R21317 vp_p.n15729 vp_p.n15728 0.006
R21318 vp_p.n15739 vp_p.n15733 0.006
R21319 vp_p.n15743 vp_p.n15742 0.006
R21320 vp_p.n15753 vp_p.n15747 0.006
R21321 vp_p.n15757 vp_p.n15756 0.006
R21322 vp_p.n15767 vp_p.n15761 0.006
R21323 vp_p.n15771 vp_p.n15770 0.006
R21324 vp_p.n15781 vp_p.n15775 0.006
R21325 vp_p.n15785 vp_p.n15784 0.006
R21326 vp_p.n15795 vp_p.n15789 0.006
R21327 vp_p.n15799 vp_p.n15798 0.006
R21328 vp_p.n15809 vp_p.n15803 0.006
R21329 vp_p.n15813 vp_p.n15812 0.006
R21330 vp_p.n15817 vp_p.n15816 0.006
R21331 vp_p.n15827 vp_p.n15821 0.006
R21332 vp_p.n15831 vp_p.n15830 0.006
R21333 vp_p.n15836 vp_p.n15835 0.006
R21334 vp_p.n15841 vp_p.n15840 0.006
R21335 vp_p.n15846 vp_p.n15845 0.006
R21336 vp_p.n15851 vp_p.n15850 0.006
R21337 vp_p.n15856 vp_p.n15855 0.006
R21338 vp_p.n15861 vp_p.n15860 0.006
R21339 vp_p.n15866 vp_p.n15865 0.006
R21340 vp_p.n15871 vp_p.n15870 0.006
R21341 vp_p.n15876 vp_p.n15875 0.006
R21342 vp_p.n15881 vp_p.n15880 0.006
R21343 vp_p.n15886 vp_p.n15885 0.006
R21344 vp_p.n15891 vp_p.n15890 0.006
R21345 vp_p.n15896 vp_p.n15895 0.006
R21346 vp_p.n15818 vp_p.n15817 0.006
R21347 vp_p.n15814 vp_p.n15813 0.006
R21348 vp_p.n15803 vp_p.n15802 0.006
R21349 vp_p.n15800 vp_p.n15799 0.006
R21350 vp_p.n15789 vp_p.n15788 0.006
R21351 vp_p.n15786 vp_p.n15785 0.006
R21352 vp_p.n15775 vp_p.n15774 0.006
R21353 vp_p.n15772 vp_p.n15771 0.006
R21354 vp_p.n15761 vp_p.n15760 0.006
R21355 vp_p.n15758 vp_p.n15757 0.006
R21356 vp_p.n15747 vp_p.n15746 0.006
R21357 vp_p.n15744 vp_p.n15743 0.006
R21358 vp_p.n15733 vp_p.n15732 0.006
R21359 vp_p.n15730 vp_p.n15729 0.006
R21360 vp_p.n15719 vp_p.n15718 0.006
R21361 vp_p.n15716 vp_p.n15715 0.006
R21362 vp_p.n15705 vp_p.n15704 0.006
R21363 vp_p.n15702 vp_p.n15701 0.006
R21364 vp_p.n15691 vp_p.n15690 0.006
R21365 vp_p.n15688 vp_p.n15687 0.006
R21366 vp_p.n15677 vp_p.n15676 0.006
R21367 vp_p.n15674 vp_p.n15673 0.006
R21368 vp_p.n15663 vp_p.n15662 0.006
R21369 vp_p.n15660 vp_p.n15659 0.006
R21370 vp_p.n15649 vp_p.n15648 0.006
R21371 vp_p.n15646 vp_p.n15645 0.006
R21372 vp_p.n15635 vp_p.n15634 0.006
R21373 vp_p.n15632 vp_p.n15631 0.006
R21374 vp_p.n15621 vp_p.n15620 0.006
R21375 vp_p.n15618 vp_p.n15617 0.006
R21376 vp_p.n15607 vp_p.n15606 0.006
R21377 vp_p.n15604 vp_p.n15603 0.006
R21378 vp_p.n15593 vp_p.n15592 0.006
R21379 vp_p.n15590 vp_p.n15589 0.006
R21380 vp_p.n15579 vp_p.n15578 0.006
R21381 vp_p.n15576 vp_p.n15575 0.006
R21382 vp_p.n15565 vp_p.n15564 0.006
R21383 vp_p.n15562 vp_p.n15561 0.006
R21384 vp_p.n15551 vp_p.n15550 0.006
R21385 vp_p.n15548 vp_p.n15547 0.006
R21386 vp_p.n15537 vp_p.n15536 0.006
R21387 vp_p.n15534 vp_p.n15533 0.006
R21388 vp_p.n15523 vp_p.n15522 0.006
R21389 vp_p.n15520 vp_p.n15519 0.006
R21390 vp_p.n15509 vp_p.n15508 0.006
R21391 vp_p.n15506 vp_p.n15505 0.006
R21392 vp_p.n15495 vp_p.n15494 0.006
R21393 vp_p.n15492 vp_p.n15491 0.006
R21394 vp_p.n15481 vp_p.n15480 0.006
R21395 vp_p.n15478 vp_p.n15477 0.006
R21396 vp_p.n15467 vp_p.n15466 0.006
R21397 vp_p.n15464 vp_p.n15463 0.006
R21398 vp_p.n15453 vp_p.n15452 0.006
R21399 vp_p.n15450 vp_p.n15449 0.006
R21400 vp_p.n15439 vp_p.n15438 0.006
R21401 vp_p.n15436 vp_p.n15435 0.006
R21402 vp_p.n15425 vp_p.n15424 0.006
R21403 vp_p.n15422 vp_p.n15421 0.006
R21404 vp_p.n15411 vp_p.n15410 0.006
R21405 vp_p.n15408 vp_p.n15407 0.006
R21406 vp_p.n15397 vp_p.n15396 0.006
R21407 vp_p.n15394 vp_p.n15393 0.006
R21408 vp_p.n15383 vp_p.n15382 0.006
R21409 vp_p.n15380 vp_p.n15379 0.006
R21410 vp_p.n15369 vp_p.n15368 0.006
R21411 vp_p.n15366 vp_p.n15365 0.006
R21412 vp_p.n15355 vp_p.n15354 0.006
R21413 vp_p.n15352 vp_p.n15351 0.006
R21414 vp_p.n15341 vp_p.n15340 0.006
R21415 vp_p.n15338 vp_p.n15337 0.006
R21416 vp_p.n15327 vp_p.n15326 0.006
R21417 vp_p.n15324 vp_p.n15323 0.006
R21418 vp_p.n15313 vp_p.n15312 0.006
R21419 vp_p.n15310 vp_p.n15309 0.006
R21420 vp_p.n15299 vp_p.n15298 0.006
R21421 vp_p.n15296 vp_p.n15295 0.006
R21422 vp_p.n15285 vp_p.n15284 0.006
R21423 vp_p.n15282 vp_p.n15281 0.006
R21424 vp_p.n15271 vp_p.n15270 0.006
R21425 vp_p.n15268 vp_p.n15267 0.006
R21426 vp_p.n15257 vp_p.n15256 0.006
R21427 vp_p.n15254 vp_p.n15253 0.006
R21428 vp_p.n15243 vp_p.n15242 0.006
R21429 vp_p.n15240 vp_p.n15239 0.006
R21430 vp_p.n15229 vp_p.n15228 0.006
R21431 vp_p.n15226 vp_p.n15225 0.006
R21432 vp_p.n15215 vp_p.n15214 0.006
R21433 vp_p.n15212 vp_p.n15211 0.006
R21434 vp_p.n15201 vp_p.n15200 0.006
R21435 vp_p.n15198 vp_p.n15197 0.006
R21436 vp_p.n15187 vp_p.n15186 0.006
R21437 vp_p.n15184 vp_p.n15183 0.006
R21438 vp_p.n15173 vp_p.n15172 0.006
R21439 vp_p.n15170 vp_p.n15169 0.006
R21440 vp_p.n15159 vp_p.n15158 0.006
R21441 vp_p.n15156 vp_p.n15155 0.006
R21442 vp_p.n15145 vp_p.n15144 0.006
R21443 vp_p.n15142 vp_p.n15141 0.006
R21444 vp_p.n15131 vp_p.n15130 0.006
R21445 vp_p.n15128 vp_p.n15127 0.006
R21446 vp_p.n15117 vp_p.n15116 0.006
R21447 vp_p.n15114 vp_p.n15113 0.006
R21448 vp_p.n15103 vp_p.n15102 0.006
R21449 vp_p.n15100 vp_p.n15099 0.006
R21450 vp_p.n15089 vp_p.n15088 0.006
R21451 vp_p.n15086 vp_p.n15085 0.006
R21452 vp_p.n15075 vp_p.n15074 0.006
R21453 vp_p.n15072 vp_p.n15071 0.006
R21454 vp_p.n15061 vp_p.n15060 0.006
R21455 vp_p.n15058 vp_p.n15057 0.006
R21456 vp_p.n15047 vp_p.n15046 0.006
R21457 vp_p.n15044 vp_p.n15043 0.006
R21458 vp_p.n15033 vp_p.n15032 0.006
R21459 vp_p.n15030 vp_p.n15029 0.006
R21460 vp_p.n15019 vp_p.n15018 0.006
R21461 vp_p.n15016 vp_p.n15015 0.006
R21462 vp_p.n15005 vp_p.n15004 0.006
R21463 vp_p.n15002 vp_p.n15001 0.006
R21464 vp_p.n14991 vp_p.n14990 0.006
R21465 vp_p.n14988 vp_p.n14987 0.006
R21466 vp_p.n14977 vp_p.n14976 0.006
R21467 vp_p.n14974 vp_p.n14973 0.006
R21468 vp_p.n14963 vp_p.n14962 0.006
R21469 vp_p.n14960 vp_p.n14959 0.006
R21470 vp_p.n14949 vp_p.n14948 0.006
R21471 vp_p.n14946 vp_p.n14945 0.006
R21472 vp_p.n14935 vp_p.n14934 0.006
R21473 vp_p.n14932 vp_p.n14931 0.006
R21474 vp_p.n14921 vp_p.n14920 0.006
R21475 vp_p.n14918 vp_p.n14917 0.006
R21476 vp_p.n14907 vp_p.n14906 0.006
R21477 vp_p.n14904 vp_p.n14903 0.006
R21478 vp_p.n14893 vp_p.n14892 0.006
R21479 vp_p.n15821 vp_p.n15820 0.006
R21480 vp_p.n14394 vp_p.n14393 0.006
R21481 vp_p.n13025 vp_p.n13024 0.006
R21482 vp_p.n10642 vp_p.n10641 0.006
R21483 vp_p.n10647 vp_p.n10646 0.006
R21484 vp_p.n10658 vp_p.n10652 0.006
R21485 vp_p.n10662 vp_p.n10661 0.006
R21486 vp_p.n10672 vp_p.n10666 0.006
R21487 vp_p.n10676 vp_p.n10675 0.006
R21488 vp_p.n10686 vp_p.n10680 0.006
R21489 vp_p.n10690 vp_p.n10689 0.006
R21490 vp_p.n10700 vp_p.n10694 0.006
R21491 vp_p.n10704 vp_p.n10703 0.006
R21492 vp_p.n10714 vp_p.n10708 0.006
R21493 vp_p.n10718 vp_p.n10717 0.006
R21494 vp_p.n10728 vp_p.n10722 0.006
R21495 vp_p.n10732 vp_p.n10731 0.006
R21496 vp_p.n10742 vp_p.n10736 0.006
R21497 vp_p.n10746 vp_p.n10745 0.006
R21498 vp_p.n10756 vp_p.n10750 0.006
R21499 vp_p.n10760 vp_p.n10759 0.006
R21500 vp_p.n10770 vp_p.n10764 0.006
R21501 vp_p.n10774 vp_p.n10773 0.006
R21502 vp_p.n10784 vp_p.n10778 0.006
R21503 vp_p.n10788 vp_p.n10787 0.006
R21504 vp_p.n10798 vp_p.n10792 0.006
R21505 vp_p.n10802 vp_p.n10801 0.006
R21506 vp_p.n10812 vp_p.n10806 0.006
R21507 vp_p.n10816 vp_p.n10815 0.006
R21508 vp_p.n10826 vp_p.n10820 0.006
R21509 vp_p.n10830 vp_p.n10829 0.006
R21510 vp_p.n10840 vp_p.n10834 0.006
R21511 vp_p.n10844 vp_p.n10843 0.006
R21512 vp_p.n10854 vp_p.n10848 0.006
R21513 vp_p.n10858 vp_p.n10857 0.006
R21514 vp_p.n10868 vp_p.n10862 0.006
R21515 vp_p.n10872 vp_p.n10871 0.006
R21516 vp_p.n10882 vp_p.n10876 0.006
R21517 vp_p.n10886 vp_p.n10885 0.006
R21518 vp_p.n10896 vp_p.n10890 0.006
R21519 vp_p.n10900 vp_p.n10899 0.006
R21520 vp_p.n10910 vp_p.n10904 0.006
R21521 vp_p.n10914 vp_p.n10913 0.006
R21522 vp_p.n10924 vp_p.n10918 0.006
R21523 vp_p.n10928 vp_p.n10927 0.006
R21524 vp_p.n10938 vp_p.n10932 0.006
R21525 vp_p.n10942 vp_p.n10941 0.006
R21526 vp_p.n10952 vp_p.n10946 0.006
R21527 vp_p.n10956 vp_p.n10955 0.006
R21528 vp_p.n10966 vp_p.n10960 0.006
R21529 vp_p.n10970 vp_p.n10969 0.006
R21530 vp_p.n10980 vp_p.n10974 0.006
R21531 vp_p.n10984 vp_p.n10983 0.006
R21532 vp_p.n10994 vp_p.n10988 0.006
R21533 vp_p.n10998 vp_p.n10997 0.006
R21534 vp_p.n11008 vp_p.n11002 0.006
R21535 vp_p.n11012 vp_p.n11011 0.006
R21536 vp_p.n11022 vp_p.n11016 0.006
R21537 vp_p.n11026 vp_p.n11025 0.006
R21538 vp_p.n11036 vp_p.n11030 0.006
R21539 vp_p.n11040 vp_p.n11039 0.006
R21540 vp_p.n11050 vp_p.n11044 0.006
R21541 vp_p.n11054 vp_p.n11053 0.006
R21542 vp_p.n11064 vp_p.n11058 0.006
R21543 vp_p.n11068 vp_p.n11067 0.006
R21544 vp_p.n11078 vp_p.n11072 0.006
R21545 vp_p.n11082 vp_p.n11081 0.006
R21546 vp_p.n11092 vp_p.n11086 0.006
R21547 vp_p.n11096 vp_p.n11095 0.006
R21548 vp_p.n11106 vp_p.n11100 0.006
R21549 vp_p.n11110 vp_p.n11109 0.006
R21550 vp_p.n11120 vp_p.n11114 0.006
R21551 vp_p.n11124 vp_p.n11123 0.006
R21552 vp_p.n11134 vp_p.n11128 0.006
R21553 vp_p.n11138 vp_p.n11137 0.006
R21554 vp_p.n11148 vp_p.n11142 0.006
R21555 vp_p.n11152 vp_p.n11151 0.006
R21556 vp_p.n11162 vp_p.n11156 0.006
R21557 vp_p.n11166 vp_p.n11165 0.006
R21558 vp_p.n11176 vp_p.n11170 0.006
R21559 vp_p.n11180 vp_p.n11179 0.006
R21560 vp_p.n11190 vp_p.n11184 0.006
R21561 vp_p.n11194 vp_p.n11193 0.006
R21562 vp_p.n11204 vp_p.n11198 0.006
R21563 vp_p.n11208 vp_p.n11207 0.006
R21564 vp_p.n11218 vp_p.n11212 0.006
R21565 vp_p.n11222 vp_p.n11221 0.006
R21566 vp_p.n11232 vp_p.n11226 0.006
R21567 vp_p.n11236 vp_p.n11235 0.006
R21568 vp_p.n11246 vp_p.n11240 0.006
R21569 vp_p.n11250 vp_p.n11249 0.006
R21570 vp_p.n11260 vp_p.n11254 0.006
R21571 vp_p.n11264 vp_p.n11263 0.006
R21572 vp_p.n11274 vp_p.n11268 0.006
R21573 vp_p.n11278 vp_p.n11277 0.006
R21574 vp_p.n11288 vp_p.n11282 0.006
R21575 vp_p.n11292 vp_p.n11291 0.006
R21576 vp_p.n11302 vp_p.n11296 0.006
R21577 vp_p.n11306 vp_p.n11305 0.006
R21578 vp_p.n11316 vp_p.n11310 0.006
R21579 vp_p.n11320 vp_p.n11319 0.006
R21580 vp_p.n11330 vp_p.n11324 0.006
R21581 vp_p.n11334 vp_p.n11333 0.006
R21582 vp_p.n11344 vp_p.n11338 0.006
R21583 vp_p.n11348 vp_p.n11347 0.006
R21584 vp_p.n11358 vp_p.n11352 0.006
R21585 vp_p.n11362 vp_p.n11361 0.006
R21586 vp_p.n11372 vp_p.n11366 0.006
R21587 vp_p.n11376 vp_p.n11375 0.006
R21588 vp_p.n11386 vp_p.n11380 0.006
R21589 vp_p.n11390 vp_p.n11389 0.006
R21590 vp_p.n11400 vp_p.n11394 0.006
R21591 vp_p.n11404 vp_p.n11403 0.006
R21592 vp_p.n11414 vp_p.n11408 0.006
R21593 vp_p.n11418 vp_p.n11417 0.006
R21594 vp_p.n11428 vp_p.n11422 0.006
R21595 vp_p.n11432 vp_p.n11431 0.006
R21596 vp_p.n11442 vp_p.n11436 0.006
R21597 vp_p.n11446 vp_p.n11445 0.006
R21598 vp_p.n11456 vp_p.n11450 0.006
R21599 vp_p.n11460 vp_p.n11459 0.006
R21600 vp_p.n11470 vp_p.n11464 0.006
R21601 vp_p.n11474 vp_p.n11473 0.006
R21602 vp_p.n11484 vp_p.n11478 0.006
R21603 vp_p.n11488 vp_p.n11487 0.006
R21604 vp_p.n11498 vp_p.n11492 0.006
R21605 vp_p.n11502 vp_p.n11501 0.006
R21606 vp_p.n11512 vp_p.n11506 0.006
R21607 vp_p.n11516 vp_p.n11515 0.006
R21608 vp_p.n11526 vp_p.n11520 0.006
R21609 vp_p.n11530 vp_p.n11529 0.006
R21610 vp_p.n11540 vp_p.n11534 0.006
R21611 vp_p.n11544 vp_p.n11543 0.006
R21612 vp_p.n11554 vp_p.n11548 0.006
R21613 vp_p.n11558 vp_p.n11557 0.006
R21614 vp_p.n11568 vp_p.n11562 0.006
R21615 vp_p.n11572 vp_p.n11571 0.006
R21616 vp_p.n11582 vp_p.n11576 0.006
R21617 vp_p.n11586 vp_p.n11585 0.006
R21618 vp_p.n11596 vp_p.n11590 0.006
R21619 vp_p.n11600 vp_p.n11599 0.006
R21620 vp_p.n11605 vp_p.n11604 0.006
R21621 vp_p.n11610 vp_p.n11609 0.006
R21622 vp_p.n11615 vp_p.n11614 0.006
R21623 vp_p.n11620 vp_p.n11619 0.006
R21624 vp_p.n11625 vp_p.n11624 0.006
R21625 vp_p.n11630 vp_p.n11629 0.006
R21626 vp_p.n11635 vp_p.n11634 0.006
R21627 vp_p.n11640 vp_p.n11639 0.006
R21628 vp_p.n11645 vp_p.n11644 0.006
R21629 vp_p.n11650 vp_p.n11649 0.006
R21630 vp_p.n11655 vp_p.n11654 0.006
R21631 vp_p.n11660 vp_p.n11659 0.006
R21632 vp_p.n11587 vp_p.n11586 0.006
R21633 vp_p.n11576 vp_p.n11575 0.006
R21634 vp_p.n11573 vp_p.n11572 0.006
R21635 vp_p.n11562 vp_p.n11561 0.006
R21636 vp_p.n11559 vp_p.n11558 0.006
R21637 vp_p.n11548 vp_p.n11547 0.006
R21638 vp_p.n11545 vp_p.n11544 0.006
R21639 vp_p.n11534 vp_p.n11533 0.006
R21640 vp_p.n11531 vp_p.n11530 0.006
R21641 vp_p.n11520 vp_p.n11519 0.006
R21642 vp_p.n11517 vp_p.n11516 0.006
R21643 vp_p.n11506 vp_p.n11505 0.006
R21644 vp_p.n11503 vp_p.n11502 0.006
R21645 vp_p.n11492 vp_p.n11491 0.006
R21646 vp_p.n11489 vp_p.n11488 0.006
R21647 vp_p.n11478 vp_p.n11477 0.006
R21648 vp_p.n11475 vp_p.n11474 0.006
R21649 vp_p.n11464 vp_p.n11463 0.006
R21650 vp_p.n11461 vp_p.n11460 0.006
R21651 vp_p.n11450 vp_p.n11449 0.006
R21652 vp_p.n11447 vp_p.n11446 0.006
R21653 vp_p.n11436 vp_p.n11435 0.006
R21654 vp_p.n11433 vp_p.n11432 0.006
R21655 vp_p.n11422 vp_p.n11421 0.006
R21656 vp_p.n11419 vp_p.n11418 0.006
R21657 vp_p.n11408 vp_p.n11407 0.006
R21658 vp_p.n11405 vp_p.n11404 0.006
R21659 vp_p.n11394 vp_p.n11393 0.006
R21660 vp_p.n11391 vp_p.n11390 0.006
R21661 vp_p.n11380 vp_p.n11379 0.006
R21662 vp_p.n11377 vp_p.n11376 0.006
R21663 vp_p.n11366 vp_p.n11365 0.006
R21664 vp_p.n11363 vp_p.n11362 0.006
R21665 vp_p.n11352 vp_p.n11351 0.006
R21666 vp_p.n11349 vp_p.n11348 0.006
R21667 vp_p.n11338 vp_p.n11337 0.006
R21668 vp_p.n11335 vp_p.n11334 0.006
R21669 vp_p.n11324 vp_p.n11323 0.006
R21670 vp_p.n11321 vp_p.n11320 0.006
R21671 vp_p.n11310 vp_p.n11309 0.006
R21672 vp_p.n11307 vp_p.n11306 0.006
R21673 vp_p.n11296 vp_p.n11295 0.006
R21674 vp_p.n11293 vp_p.n11292 0.006
R21675 vp_p.n11282 vp_p.n11281 0.006
R21676 vp_p.n11279 vp_p.n11278 0.006
R21677 vp_p.n11268 vp_p.n11267 0.006
R21678 vp_p.n11265 vp_p.n11264 0.006
R21679 vp_p.n11254 vp_p.n11253 0.006
R21680 vp_p.n11251 vp_p.n11250 0.006
R21681 vp_p.n11240 vp_p.n11239 0.006
R21682 vp_p.n11237 vp_p.n11236 0.006
R21683 vp_p.n11226 vp_p.n11225 0.006
R21684 vp_p.n11223 vp_p.n11222 0.006
R21685 vp_p.n11212 vp_p.n11211 0.006
R21686 vp_p.n11209 vp_p.n11208 0.006
R21687 vp_p.n11198 vp_p.n11197 0.006
R21688 vp_p.n11195 vp_p.n11194 0.006
R21689 vp_p.n11184 vp_p.n11183 0.006
R21690 vp_p.n11181 vp_p.n11180 0.006
R21691 vp_p.n11170 vp_p.n11169 0.006
R21692 vp_p.n11167 vp_p.n11166 0.006
R21693 vp_p.n11156 vp_p.n11155 0.006
R21694 vp_p.n11153 vp_p.n11152 0.006
R21695 vp_p.n11142 vp_p.n11141 0.006
R21696 vp_p.n11139 vp_p.n11138 0.006
R21697 vp_p.n11128 vp_p.n11127 0.006
R21698 vp_p.n11125 vp_p.n11124 0.006
R21699 vp_p.n11114 vp_p.n11113 0.006
R21700 vp_p.n11111 vp_p.n11110 0.006
R21701 vp_p.n11100 vp_p.n11099 0.006
R21702 vp_p.n11097 vp_p.n11096 0.006
R21703 vp_p.n11086 vp_p.n11085 0.006
R21704 vp_p.n11083 vp_p.n11082 0.006
R21705 vp_p.n11072 vp_p.n11071 0.006
R21706 vp_p.n11069 vp_p.n11068 0.006
R21707 vp_p.n11058 vp_p.n11057 0.006
R21708 vp_p.n11055 vp_p.n11054 0.006
R21709 vp_p.n11044 vp_p.n11043 0.006
R21710 vp_p.n11041 vp_p.n11040 0.006
R21711 vp_p.n11030 vp_p.n11029 0.006
R21712 vp_p.n11027 vp_p.n11026 0.006
R21713 vp_p.n11016 vp_p.n11015 0.006
R21714 vp_p.n11013 vp_p.n11012 0.006
R21715 vp_p.n11002 vp_p.n11001 0.006
R21716 vp_p.n10999 vp_p.n10998 0.006
R21717 vp_p.n10988 vp_p.n10987 0.006
R21718 vp_p.n10985 vp_p.n10984 0.006
R21719 vp_p.n10974 vp_p.n10973 0.006
R21720 vp_p.n10971 vp_p.n10970 0.006
R21721 vp_p.n10960 vp_p.n10959 0.006
R21722 vp_p.n10957 vp_p.n10956 0.006
R21723 vp_p.n10946 vp_p.n10945 0.006
R21724 vp_p.n10943 vp_p.n10942 0.006
R21725 vp_p.n10932 vp_p.n10931 0.006
R21726 vp_p.n10929 vp_p.n10928 0.006
R21727 vp_p.n10918 vp_p.n10917 0.006
R21728 vp_p.n10915 vp_p.n10914 0.006
R21729 vp_p.n10904 vp_p.n10903 0.006
R21730 vp_p.n10901 vp_p.n10900 0.006
R21731 vp_p.n10890 vp_p.n10889 0.006
R21732 vp_p.n10887 vp_p.n10886 0.006
R21733 vp_p.n10876 vp_p.n10875 0.006
R21734 vp_p.n10873 vp_p.n10872 0.006
R21735 vp_p.n10862 vp_p.n10861 0.006
R21736 vp_p.n10859 vp_p.n10858 0.006
R21737 vp_p.n10848 vp_p.n10847 0.006
R21738 vp_p.n10845 vp_p.n10844 0.006
R21739 vp_p.n10834 vp_p.n10833 0.006
R21740 vp_p.n10831 vp_p.n10830 0.006
R21741 vp_p.n10820 vp_p.n10819 0.006
R21742 vp_p.n10817 vp_p.n10816 0.006
R21743 vp_p.n10806 vp_p.n10805 0.006
R21744 vp_p.n10803 vp_p.n10802 0.006
R21745 vp_p.n10792 vp_p.n10791 0.006
R21746 vp_p.n10789 vp_p.n10788 0.006
R21747 vp_p.n10778 vp_p.n10777 0.006
R21748 vp_p.n10775 vp_p.n10774 0.006
R21749 vp_p.n10764 vp_p.n10763 0.006
R21750 vp_p.n10761 vp_p.n10760 0.006
R21751 vp_p.n10750 vp_p.n10749 0.006
R21752 vp_p.n10747 vp_p.n10746 0.006
R21753 vp_p.n10736 vp_p.n10735 0.006
R21754 vp_p.n10733 vp_p.n10732 0.006
R21755 vp_p.n10722 vp_p.n10721 0.006
R21756 vp_p.n10719 vp_p.n10718 0.006
R21757 vp_p.n10708 vp_p.n10707 0.006
R21758 vp_p.n10705 vp_p.n10704 0.006
R21759 vp_p.n10694 vp_p.n10693 0.006
R21760 vp_p.n10691 vp_p.n10690 0.006
R21761 vp_p.n10680 vp_p.n10679 0.006
R21762 vp_p.n10677 vp_p.n10676 0.006
R21763 vp_p.n10666 vp_p.n10665 0.006
R21764 vp_p.n10663 vp_p.n10662 0.006
R21765 vp_p.n10652 vp_p.n10651 0.006
R21766 vp_p.n11590 vp_p.n11589 0.006
R21767 vp_p.n13030 vp_p.n13029 0.006
R21768 vp_p.n14399 vp_p.n14398 0.006
R21769 vp_p.n15832 vp_p.n15831 0.006
R21770 vp_p.n16311 vp_p.n16310 0.006
R21771 vp_p.n16316 vp_p.n16315 0.006
R21772 vp_p.n16327 vp_p.n16321 0.006
R21773 vp_p.n16331 vp_p.n16330 0.006
R21774 vp_p.n16341 vp_p.n16335 0.006
R21775 vp_p.n16345 vp_p.n16344 0.006
R21776 vp_p.n16355 vp_p.n16349 0.006
R21777 vp_p.n16359 vp_p.n16358 0.006
R21778 vp_p.n16369 vp_p.n16363 0.006
R21779 vp_p.n16373 vp_p.n16372 0.006
R21780 vp_p.n16383 vp_p.n16377 0.006
R21781 vp_p.n16387 vp_p.n16386 0.006
R21782 vp_p.n16397 vp_p.n16391 0.006
R21783 vp_p.n16401 vp_p.n16400 0.006
R21784 vp_p.n16411 vp_p.n16405 0.006
R21785 vp_p.n16415 vp_p.n16414 0.006
R21786 vp_p.n16425 vp_p.n16419 0.006
R21787 vp_p.n16429 vp_p.n16428 0.006
R21788 vp_p.n16439 vp_p.n16433 0.006
R21789 vp_p.n16443 vp_p.n16442 0.006
R21790 vp_p.n16453 vp_p.n16447 0.006
R21791 vp_p.n16457 vp_p.n16456 0.006
R21792 vp_p.n16467 vp_p.n16461 0.006
R21793 vp_p.n16471 vp_p.n16470 0.006
R21794 vp_p.n16481 vp_p.n16475 0.006
R21795 vp_p.n16485 vp_p.n16484 0.006
R21796 vp_p.n16495 vp_p.n16489 0.006
R21797 vp_p.n16499 vp_p.n16498 0.006
R21798 vp_p.n16509 vp_p.n16503 0.006
R21799 vp_p.n16513 vp_p.n16512 0.006
R21800 vp_p.n16523 vp_p.n16517 0.006
R21801 vp_p.n16527 vp_p.n16526 0.006
R21802 vp_p.n16537 vp_p.n16531 0.006
R21803 vp_p.n16541 vp_p.n16540 0.006
R21804 vp_p.n16551 vp_p.n16545 0.006
R21805 vp_p.n16555 vp_p.n16554 0.006
R21806 vp_p.n16565 vp_p.n16559 0.006
R21807 vp_p.n16569 vp_p.n16568 0.006
R21808 vp_p.n16579 vp_p.n16573 0.006
R21809 vp_p.n16583 vp_p.n16582 0.006
R21810 vp_p.n16593 vp_p.n16587 0.006
R21811 vp_p.n16597 vp_p.n16596 0.006
R21812 vp_p.n16607 vp_p.n16601 0.006
R21813 vp_p.n16611 vp_p.n16610 0.006
R21814 vp_p.n16621 vp_p.n16615 0.006
R21815 vp_p.n16625 vp_p.n16624 0.006
R21816 vp_p.n16635 vp_p.n16629 0.006
R21817 vp_p.n16639 vp_p.n16638 0.006
R21818 vp_p.n16649 vp_p.n16643 0.006
R21819 vp_p.n16653 vp_p.n16652 0.006
R21820 vp_p.n16663 vp_p.n16657 0.006
R21821 vp_p.n16667 vp_p.n16666 0.006
R21822 vp_p.n16677 vp_p.n16671 0.006
R21823 vp_p.n16681 vp_p.n16680 0.006
R21824 vp_p.n16691 vp_p.n16685 0.006
R21825 vp_p.n16695 vp_p.n16694 0.006
R21826 vp_p.n16705 vp_p.n16699 0.006
R21827 vp_p.n16709 vp_p.n16708 0.006
R21828 vp_p.n16719 vp_p.n16713 0.006
R21829 vp_p.n16723 vp_p.n16722 0.006
R21830 vp_p.n16733 vp_p.n16727 0.006
R21831 vp_p.n16737 vp_p.n16736 0.006
R21832 vp_p.n16747 vp_p.n16741 0.006
R21833 vp_p.n16751 vp_p.n16750 0.006
R21834 vp_p.n16761 vp_p.n16755 0.006
R21835 vp_p.n16765 vp_p.n16764 0.006
R21836 vp_p.n16775 vp_p.n16769 0.006
R21837 vp_p.n16779 vp_p.n16778 0.006
R21838 vp_p.n16789 vp_p.n16783 0.006
R21839 vp_p.n16793 vp_p.n16792 0.006
R21840 vp_p.n16803 vp_p.n16797 0.006
R21841 vp_p.n16807 vp_p.n16806 0.006
R21842 vp_p.n16817 vp_p.n16811 0.006
R21843 vp_p.n16821 vp_p.n16820 0.006
R21844 vp_p.n16831 vp_p.n16825 0.006
R21845 vp_p.n16835 vp_p.n16834 0.006
R21846 vp_p.n16845 vp_p.n16839 0.006
R21847 vp_p.n16849 vp_p.n16848 0.006
R21848 vp_p.n16859 vp_p.n16853 0.006
R21849 vp_p.n16863 vp_p.n16862 0.006
R21850 vp_p.n16873 vp_p.n16867 0.006
R21851 vp_p.n16877 vp_p.n16876 0.006
R21852 vp_p.n16887 vp_p.n16881 0.006
R21853 vp_p.n16891 vp_p.n16890 0.006
R21854 vp_p.n16901 vp_p.n16895 0.006
R21855 vp_p.n16905 vp_p.n16904 0.006
R21856 vp_p.n16915 vp_p.n16909 0.006
R21857 vp_p.n16919 vp_p.n16918 0.006
R21858 vp_p.n16929 vp_p.n16923 0.006
R21859 vp_p.n16933 vp_p.n16932 0.006
R21860 vp_p.n16943 vp_p.n16937 0.006
R21861 vp_p.n16947 vp_p.n16946 0.006
R21862 vp_p.n16957 vp_p.n16951 0.006
R21863 vp_p.n16961 vp_p.n16960 0.006
R21864 vp_p.n16971 vp_p.n16965 0.006
R21865 vp_p.n16975 vp_p.n16974 0.006
R21866 vp_p.n16985 vp_p.n16979 0.006
R21867 vp_p.n16989 vp_p.n16988 0.006
R21868 vp_p.n16999 vp_p.n16993 0.006
R21869 vp_p.n17003 vp_p.n17002 0.006
R21870 vp_p.n17013 vp_p.n17007 0.006
R21871 vp_p.n17017 vp_p.n17016 0.006
R21872 vp_p.n17027 vp_p.n17021 0.006
R21873 vp_p.n17031 vp_p.n17030 0.006
R21874 vp_p.n17041 vp_p.n17035 0.006
R21875 vp_p.n17045 vp_p.n17044 0.006
R21876 vp_p.n17055 vp_p.n17049 0.006
R21877 vp_p.n17059 vp_p.n17058 0.006
R21878 vp_p.n17069 vp_p.n17063 0.006
R21879 vp_p.n17073 vp_p.n17072 0.006
R21880 vp_p.n17083 vp_p.n17077 0.006
R21881 vp_p.n17087 vp_p.n17086 0.006
R21882 vp_p.n17097 vp_p.n17091 0.006
R21883 vp_p.n17101 vp_p.n17100 0.006
R21884 vp_p.n17111 vp_p.n17105 0.006
R21885 vp_p.n17115 vp_p.n17114 0.006
R21886 vp_p.n17125 vp_p.n17119 0.006
R21887 vp_p.n17129 vp_p.n17128 0.006
R21888 vp_p.n17139 vp_p.n17133 0.006
R21889 vp_p.n17143 vp_p.n17142 0.006
R21890 vp_p.n17153 vp_p.n17147 0.006
R21891 vp_p.n17157 vp_p.n17156 0.006
R21892 vp_p.n17167 vp_p.n17161 0.006
R21893 vp_p.n17171 vp_p.n17170 0.006
R21894 vp_p.n17181 vp_p.n17175 0.006
R21895 vp_p.n17185 vp_p.n17184 0.006
R21896 vp_p.n17195 vp_p.n17189 0.006
R21897 vp_p.n17199 vp_p.n17198 0.006
R21898 vp_p.n17209 vp_p.n17203 0.006
R21899 vp_p.n17213 vp_p.n17212 0.006
R21900 vp_p.n17223 vp_p.n17217 0.006
R21901 vp_p.n17227 vp_p.n17226 0.006
R21902 vp_p.n17237 vp_p.n17231 0.006
R21903 vp_p.n17241 vp_p.n17240 0.006
R21904 vp_p.n17251 vp_p.n17245 0.006
R21905 vp_p.n17255 vp_p.n17254 0.006
R21906 vp_p.n17259 vp_p.n17258 0.006
R21907 vp_p.n17269 vp_p.n17263 0.006
R21908 vp_p.n17273 vp_p.n17272 0.006
R21909 vp_p.n17278 vp_p.n17277 0.006
R21910 vp_p.n17283 vp_p.n17282 0.006
R21911 vp_p.n17288 vp_p.n17287 0.006
R21912 vp_p.n17293 vp_p.n17292 0.006
R21913 vp_p.n17298 vp_p.n17297 0.006
R21914 vp_p.n17303 vp_p.n17302 0.006
R21915 vp_p.n17308 vp_p.n17307 0.006
R21916 vp_p.n17313 vp_p.n17312 0.006
R21917 vp_p.n17318 vp_p.n17317 0.006
R21918 vp_p.n17323 vp_p.n17322 0.006
R21919 vp_p.n17328 vp_p.n17327 0.006
R21920 vp_p.n17260 vp_p.n17259 0.006
R21921 vp_p.n17256 vp_p.n17255 0.006
R21922 vp_p.n17245 vp_p.n17244 0.006
R21923 vp_p.n17242 vp_p.n17241 0.006
R21924 vp_p.n17231 vp_p.n17230 0.006
R21925 vp_p.n17228 vp_p.n17227 0.006
R21926 vp_p.n17217 vp_p.n17216 0.006
R21927 vp_p.n17214 vp_p.n17213 0.006
R21928 vp_p.n17203 vp_p.n17202 0.006
R21929 vp_p.n17200 vp_p.n17199 0.006
R21930 vp_p.n17189 vp_p.n17188 0.006
R21931 vp_p.n17186 vp_p.n17185 0.006
R21932 vp_p.n17175 vp_p.n17174 0.006
R21933 vp_p.n17172 vp_p.n17171 0.006
R21934 vp_p.n17161 vp_p.n17160 0.006
R21935 vp_p.n17158 vp_p.n17157 0.006
R21936 vp_p.n17147 vp_p.n17146 0.006
R21937 vp_p.n17144 vp_p.n17143 0.006
R21938 vp_p.n17133 vp_p.n17132 0.006
R21939 vp_p.n17130 vp_p.n17129 0.006
R21940 vp_p.n17119 vp_p.n17118 0.006
R21941 vp_p.n17116 vp_p.n17115 0.006
R21942 vp_p.n17105 vp_p.n17104 0.006
R21943 vp_p.n17102 vp_p.n17101 0.006
R21944 vp_p.n17091 vp_p.n17090 0.006
R21945 vp_p.n17088 vp_p.n17087 0.006
R21946 vp_p.n17077 vp_p.n17076 0.006
R21947 vp_p.n17074 vp_p.n17073 0.006
R21948 vp_p.n17063 vp_p.n17062 0.006
R21949 vp_p.n17060 vp_p.n17059 0.006
R21950 vp_p.n17049 vp_p.n17048 0.006
R21951 vp_p.n17046 vp_p.n17045 0.006
R21952 vp_p.n17035 vp_p.n17034 0.006
R21953 vp_p.n17032 vp_p.n17031 0.006
R21954 vp_p.n17021 vp_p.n17020 0.006
R21955 vp_p.n17018 vp_p.n17017 0.006
R21956 vp_p.n17007 vp_p.n17006 0.006
R21957 vp_p.n17004 vp_p.n17003 0.006
R21958 vp_p.n16993 vp_p.n16992 0.006
R21959 vp_p.n16990 vp_p.n16989 0.006
R21960 vp_p.n16979 vp_p.n16978 0.006
R21961 vp_p.n16976 vp_p.n16975 0.006
R21962 vp_p.n16965 vp_p.n16964 0.006
R21963 vp_p.n16962 vp_p.n16961 0.006
R21964 vp_p.n16951 vp_p.n16950 0.006
R21965 vp_p.n16948 vp_p.n16947 0.006
R21966 vp_p.n16937 vp_p.n16936 0.006
R21967 vp_p.n16934 vp_p.n16933 0.006
R21968 vp_p.n16923 vp_p.n16922 0.006
R21969 vp_p.n16920 vp_p.n16919 0.006
R21970 vp_p.n16909 vp_p.n16908 0.006
R21971 vp_p.n16906 vp_p.n16905 0.006
R21972 vp_p.n16895 vp_p.n16894 0.006
R21973 vp_p.n16892 vp_p.n16891 0.006
R21974 vp_p.n16881 vp_p.n16880 0.006
R21975 vp_p.n16878 vp_p.n16877 0.006
R21976 vp_p.n16867 vp_p.n16866 0.006
R21977 vp_p.n16864 vp_p.n16863 0.006
R21978 vp_p.n16853 vp_p.n16852 0.006
R21979 vp_p.n16850 vp_p.n16849 0.006
R21980 vp_p.n16839 vp_p.n16838 0.006
R21981 vp_p.n16836 vp_p.n16835 0.006
R21982 vp_p.n16825 vp_p.n16824 0.006
R21983 vp_p.n16822 vp_p.n16821 0.006
R21984 vp_p.n16811 vp_p.n16810 0.006
R21985 vp_p.n16808 vp_p.n16807 0.006
R21986 vp_p.n16797 vp_p.n16796 0.006
R21987 vp_p.n16794 vp_p.n16793 0.006
R21988 vp_p.n16783 vp_p.n16782 0.006
R21989 vp_p.n16780 vp_p.n16779 0.006
R21990 vp_p.n16769 vp_p.n16768 0.006
R21991 vp_p.n16766 vp_p.n16765 0.006
R21992 vp_p.n16755 vp_p.n16754 0.006
R21993 vp_p.n16752 vp_p.n16751 0.006
R21994 vp_p.n16741 vp_p.n16740 0.006
R21995 vp_p.n16738 vp_p.n16737 0.006
R21996 vp_p.n16727 vp_p.n16726 0.006
R21997 vp_p.n16724 vp_p.n16723 0.006
R21998 vp_p.n16713 vp_p.n16712 0.006
R21999 vp_p.n16710 vp_p.n16709 0.006
R22000 vp_p.n16699 vp_p.n16698 0.006
R22001 vp_p.n16696 vp_p.n16695 0.006
R22002 vp_p.n16685 vp_p.n16684 0.006
R22003 vp_p.n16682 vp_p.n16681 0.006
R22004 vp_p.n16671 vp_p.n16670 0.006
R22005 vp_p.n16668 vp_p.n16667 0.006
R22006 vp_p.n16657 vp_p.n16656 0.006
R22007 vp_p.n16654 vp_p.n16653 0.006
R22008 vp_p.n16643 vp_p.n16642 0.006
R22009 vp_p.n16640 vp_p.n16639 0.006
R22010 vp_p.n16629 vp_p.n16628 0.006
R22011 vp_p.n16626 vp_p.n16625 0.006
R22012 vp_p.n16615 vp_p.n16614 0.006
R22013 vp_p.n16612 vp_p.n16611 0.006
R22014 vp_p.n16601 vp_p.n16600 0.006
R22015 vp_p.n16598 vp_p.n16597 0.006
R22016 vp_p.n16587 vp_p.n16586 0.006
R22017 vp_p.n16584 vp_p.n16583 0.006
R22018 vp_p.n16573 vp_p.n16572 0.006
R22019 vp_p.n16570 vp_p.n16569 0.006
R22020 vp_p.n16559 vp_p.n16558 0.006
R22021 vp_p.n16556 vp_p.n16555 0.006
R22022 vp_p.n16545 vp_p.n16544 0.006
R22023 vp_p.n16542 vp_p.n16541 0.006
R22024 vp_p.n16531 vp_p.n16530 0.006
R22025 vp_p.n16528 vp_p.n16527 0.006
R22026 vp_p.n16517 vp_p.n16516 0.006
R22027 vp_p.n16514 vp_p.n16513 0.006
R22028 vp_p.n16503 vp_p.n16502 0.006
R22029 vp_p.n16500 vp_p.n16499 0.006
R22030 vp_p.n16489 vp_p.n16488 0.006
R22031 vp_p.n16486 vp_p.n16485 0.006
R22032 vp_p.n16475 vp_p.n16474 0.006
R22033 vp_p.n16472 vp_p.n16471 0.006
R22034 vp_p.n16461 vp_p.n16460 0.006
R22035 vp_p.n16458 vp_p.n16457 0.006
R22036 vp_p.n16447 vp_p.n16446 0.006
R22037 vp_p.n16444 vp_p.n16443 0.006
R22038 vp_p.n16433 vp_p.n16432 0.006
R22039 vp_p.n16430 vp_p.n16429 0.006
R22040 vp_p.n16419 vp_p.n16418 0.006
R22041 vp_p.n16416 vp_p.n16415 0.006
R22042 vp_p.n16405 vp_p.n16404 0.006
R22043 vp_p.n16402 vp_p.n16401 0.006
R22044 vp_p.n16391 vp_p.n16390 0.006
R22045 vp_p.n16388 vp_p.n16387 0.006
R22046 vp_p.n16377 vp_p.n16376 0.006
R22047 vp_p.n16374 vp_p.n16373 0.006
R22048 vp_p.n16363 vp_p.n16362 0.006
R22049 vp_p.n16360 vp_p.n16359 0.006
R22050 vp_p.n16349 vp_p.n16348 0.006
R22051 vp_p.n16346 vp_p.n16345 0.006
R22052 vp_p.n16335 vp_p.n16334 0.006
R22053 vp_p.n16332 vp_p.n16331 0.006
R22054 vp_p.n16321 vp_p.n16320 0.006
R22055 vp_p.n17263 vp_p.n17262 0.006
R22056 vp_p.n15837 vp_p.n15836 0.006
R22057 vp_p.n14404 vp_p.n14403 0.006
R22058 vp_p.n13035 vp_p.n13034 0.006
R22059 vp_p.n11601 vp_p.n11600 0.006
R22060 vp_p.n9205 vp_p.n9204 0.006
R22061 vp_p.n9210 vp_p.n9209 0.006
R22062 vp_p.n9221 vp_p.n9215 0.006
R22063 vp_p.n9225 vp_p.n9224 0.006
R22064 vp_p.n9235 vp_p.n9229 0.006
R22065 vp_p.n9239 vp_p.n9238 0.006
R22066 vp_p.n9249 vp_p.n9243 0.006
R22067 vp_p.n9253 vp_p.n9252 0.006
R22068 vp_p.n9263 vp_p.n9257 0.006
R22069 vp_p.n9267 vp_p.n9266 0.006
R22070 vp_p.n9277 vp_p.n9271 0.006
R22071 vp_p.n9281 vp_p.n9280 0.006
R22072 vp_p.n9291 vp_p.n9285 0.006
R22073 vp_p.n9295 vp_p.n9294 0.006
R22074 vp_p.n9305 vp_p.n9299 0.006
R22075 vp_p.n9309 vp_p.n9308 0.006
R22076 vp_p.n9319 vp_p.n9313 0.006
R22077 vp_p.n9323 vp_p.n9322 0.006
R22078 vp_p.n9333 vp_p.n9327 0.006
R22079 vp_p.n9337 vp_p.n9336 0.006
R22080 vp_p.n9347 vp_p.n9341 0.006
R22081 vp_p.n9351 vp_p.n9350 0.006
R22082 vp_p.n9361 vp_p.n9355 0.006
R22083 vp_p.n9365 vp_p.n9364 0.006
R22084 vp_p.n9375 vp_p.n9369 0.006
R22085 vp_p.n9379 vp_p.n9378 0.006
R22086 vp_p.n9389 vp_p.n9383 0.006
R22087 vp_p.n9393 vp_p.n9392 0.006
R22088 vp_p.n9403 vp_p.n9397 0.006
R22089 vp_p.n9407 vp_p.n9406 0.006
R22090 vp_p.n9417 vp_p.n9411 0.006
R22091 vp_p.n9421 vp_p.n9420 0.006
R22092 vp_p.n9431 vp_p.n9425 0.006
R22093 vp_p.n9435 vp_p.n9434 0.006
R22094 vp_p.n9445 vp_p.n9439 0.006
R22095 vp_p.n9449 vp_p.n9448 0.006
R22096 vp_p.n9459 vp_p.n9453 0.006
R22097 vp_p.n9463 vp_p.n9462 0.006
R22098 vp_p.n9473 vp_p.n9467 0.006
R22099 vp_p.n9477 vp_p.n9476 0.006
R22100 vp_p.n9487 vp_p.n9481 0.006
R22101 vp_p.n9491 vp_p.n9490 0.006
R22102 vp_p.n9501 vp_p.n9495 0.006
R22103 vp_p.n9505 vp_p.n9504 0.006
R22104 vp_p.n9515 vp_p.n9509 0.006
R22105 vp_p.n9519 vp_p.n9518 0.006
R22106 vp_p.n9529 vp_p.n9523 0.006
R22107 vp_p.n9533 vp_p.n9532 0.006
R22108 vp_p.n9543 vp_p.n9537 0.006
R22109 vp_p.n9547 vp_p.n9546 0.006
R22110 vp_p.n9557 vp_p.n9551 0.006
R22111 vp_p.n9561 vp_p.n9560 0.006
R22112 vp_p.n9571 vp_p.n9565 0.006
R22113 vp_p.n9575 vp_p.n9574 0.006
R22114 vp_p.n9585 vp_p.n9579 0.006
R22115 vp_p.n9589 vp_p.n9588 0.006
R22116 vp_p.n9599 vp_p.n9593 0.006
R22117 vp_p.n9603 vp_p.n9602 0.006
R22118 vp_p.n9613 vp_p.n9607 0.006
R22119 vp_p.n9617 vp_p.n9616 0.006
R22120 vp_p.n9627 vp_p.n9621 0.006
R22121 vp_p.n9631 vp_p.n9630 0.006
R22122 vp_p.n9641 vp_p.n9635 0.006
R22123 vp_p.n9645 vp_p.n9644 0.006
R22124 vp_p.n9655 vp_p.n9649 0.006
R22125 vp_p.n9659 vp_p.n9658 0.006
R22126 vp_p.n9669 vp_p.n9663 0.006
R22127 vp_p.n9673 vp_p.n9672 0.006
R22128 vp_p.n9683 vp_p.n9677 0.006
R22129 vp_p.n9687 vp_p.n9686 0.006
R22130 vp_p.n9697 vp_p.n9691 0.006
R22131 vp_p.n9701 vp_p.n9700 0.006
R22132 vp_p.n9711 vp_p.n9705 0.006
R22133 vp_p.n9715 vp_p.n9714 0.006
R22134 vp_p.n9725 vp_p.n9719 0.006
R22135 vp_p.n9729 vp_p.n9728 0.006
R22136 vp_p.n9739 vp_p.n9733 0.006
R22137 vp_p.n9743 vp_p.n9742 0.006
R22138 vp_p.n9753 vp_p.n9747 0.006
R22139 vp_p.n9757 vp_p.n9756 0.006
R22140 vp_p.n9767 vp_p.n9761 0.006
R22141 vp_p.n9771 vp_p.n9770 0.006
R22142 vp_p.n9781 vp_p.n9775 0.006
R22143 vp_p.n9785 vp_p.n9784 0.006
R22144 vp_p.n9795 vp_p.n9789 0.006
R22145 vp_p.n9799 vp_p.n9798 0.006
R22146 vp_p.n9809 vp_p.n9803 0.006
R22147 vp_p.n9813 vp_p.n9812 0.006
R22148 vp_p.n9823 vp_p.n9817 0.006
R22149 vp_p.n9827 vp_p.n9826 0.006
R22150 vp_p.n9837 vp_p.n9831 0.006
R22151 vp_p.n9841 vp_p.n9840 0.006
R22152 vp_p.n9851 vp_p.n9845 0.006
R22153 vp_p.n9855 vp_p.n9854 0.006
R22154 vp_p.n9865 vp_p.n9859 0.006
R22155 vp_p.n9869 vp_p.n9868 0.006
R22156 vp_p.n9879 vp_p.n9873 0.006
R22157 vp_p.n9883 vp_p.n9882 0.006
R22158 vp_p.n9893 vp_p.n9887 0.006
R22159 vp_p.n9897 vp_p.n9896 0.006
R22160 vp_p.n9907 vp_p.n9901 0.006
R22161 vp_p.n9911 vp_p.n9910 0.006
R22162 vp_p.n9921 vp_p.n9915 0.006
R22163 vp_p.n9925 vp_p.n9924 0.006
R22164 vp_p.n9935 vp_p.n9929 0.006
R22165 vp_p.n9939 vp_p.n9938 0.006
R22166 vp_p.n9949 vp_p.n9943 0.006
R22167 vp_p.n9953 vp_p.n9952 0.006
R22168 vp_p.n9963 vp_p.n9957 0.006
R22169 vp_p.n9967 vp_p.n9966 0.006
R22170 vp_p.n9977 vp_p.n9971 0.006
R22171 vp_p.n9981 vp_p.n9980 0.006
R22172 vp_p.n9991 vp_p.n9985 0.006
R22173 vp_p.n9995 vp_p.n9994 0.006
R22174 vp_p.n10005 vp_p.n9999 0.006
R22175 vp_p.n10009 vp_p.n10008 0.006
R22176 vp_p.n10019 vp_p.n10013 0.006
R22177 vp_p.n10023 vp_p.n10022 0.006
R22178 vp_p.n10033 vp_p.n10027 0.006
R22179 vp_p.n10037 vp_p.n10036 0.006
R22180 vp_p.n10047 vp_p.n10041 0.006
R22181 vp_p.n10051 vp_p.n10050 0.006
R22182 vp_p.n10061 vp_p.n10055 0.006
R22183 vp_p.n10065 vp_p.n10064 0.006
R22184 vp_p.n10075 vp_p.n10069 0.006
R22185 vp_p.n10079 vp_p.n10078 0.006
R22186 vp_p.n10089 vp_p.n10083 0.006
R22187 vp_p.n10093 vp_p.n10092 0.006
R22188 vp_p.n10103 vp_p.n10097 0.006
R22189 vp_p.n10107 vp_p.n10106 0.006
R22190 vp_p.n10117 vp_p.n10111 0.006
R22191 vp_p.n10121 vp_p.n10120 0.006
R22192 vp_p.n10131 vp_p.n10125 0.006
R22193 vp_p.n10135 vp_p.n10134 0.006
R22194 vp_p.n10145 vp_p.n10139 0.006
R22195 vp_p.n10149 vp_p.n10148 0.006
R22196 vp_p.n10159 vp_p.n10153 0.006
R22197 vp_p.n10163 vp_p.n10162 0.006
R22198 vp_p.n10173 vp_p.n10167 0.006
R22199 vp_p.n10177 vp_p.n10176 0.006
R22200 vp_p.n10182 vp_p.n10181 0.006
R22201 vp_p.n10187 vp_p.n10186 0.006
R22202 vp_p.n10192 vp_p.n10191 0.006
R22203 vp_p.n10197 vp_p.n10196 0.006
R22204 vp_p.n10202 vp_p.n10201 0.006
R22205 vp_p.n10207 vp_p.n10206 0.006
R22206 vp_p.n10212 vp_p.n10211 0.006
R22207 vp_p.n10217 vp_p.n10216 0.006
R22208 vp_p.n10222 vp_p.n10221 0.006
R22209 vp_p.n10227 vp_p.n10226 0.006
R22210 vp_p.n10164 vp_p.n10163 0.006
R22211 vp_p.n10153 vp_p.n10152 0.006
R22212 vp_p.n10150 vp_p.n10149 0.006
R22213 vp_p.n10139 vp_p.n10138 0.006
R22214 vp_p.n10136 vp_p.n10135 0.006
R22215 vp_p.n10125 vp_p.n10124 0.006
R22216 vp_p.n10122 vp_p.n10121 0.006
R22217 vp_p.n10111 vp_p.n10110 0.006
R22218 vp_p.n10108 vp_p.n10107 0.006
R22219 vp_p.n10097 vp_p.n10096 0.006
R22220 vp_p.n10094 vp_p.n10093 0.006
R22221 vp_p.n10083 vp_p.n10082 0.006
R22222 vp_p.n10080 vp_p.n10079 0.006
R22223 vp_p.n10069 vp_p.n10068 0.006
R22224 vp_p.n10066 vp_p.n10065 0.006
R22225 vp_p.n10055 vp_p.n10054 0.006
R22226 vp_p.n10052 vp_p.n10051 0.006
R22227 vp_p.n10041 vp_p.n10040 0.006
R22228 vp_p.n10038 vp_p.n10037 0.006
R22229 vp_p.n10027 vp_p.n10026 0.006
R22230 vp_p.n10024 vp_p.n10023 0.006
R22231 vp_p.n10013 vp_p.n10012 0.006
R22232 vp_p.n10010 vp_p.n10009 0.006
R22233 vp_p.n9999 vp_p.n9998 0.006
R22234 vp_p.n9996 vp_p.n9995 0.006
R22235 vp_p.n9985 vp_p.n9984 0.006
R22236 vp_p.n9982 vp_p.n9981 0.006
R22237 vp_p.n9971 vp_p.n9970 0.006
R22238 vp_p.n9968 vp_p.n9967 0.006
R22239 vp_p.n9957 vp_p.n9956 0.006
R22240 vp_p.n9954 vp_p.n9953 0.006
R22241 vp_p.n9943 vp_p.n9942 0.006
R22242 vp_p.n9940 vp_p.n9939 0.006
R22243 vp_p.n9929 vp_p.n9928 0.006
R22244 vp_p.n9926 vp_p.n9925 0.006
R22245 vp_p.n9915 vp_p.n9914 0.006
R22246 vp_p.n9912 vp_p.n9911 0.006
R22247 vp_p.n9901 vp_p.n9900 0.006
R22248 vp_p.n9898 vp_p.n9897 0.006
R22249 vp_p.n9887 vp_p.n9886 0.006
R22250 vp_p.n9884 vp_p.n9883 0.006
R22251 vp_p.n9873 vp_p.n9872 0.006
R22252 vp_p.n9870 vp_p.n9869 0.006
R22253 vp_p.n9859 vp_p.n9858 0.006
R22254 vp_p.n9856 vp_p.n9855 0.006
R22255 vp_p.n9845 vp_p.n9844 0.006
R22256 vp_p.n9842 vp_p.n9841 0.006
R22257 vp_p.n9831 vp_p.n9830 0.006
R22258 vp_p.n9828 vp_p.n9827 0.006
R22259 vp_p.n9817 vp_p.n9816 0.006
R22260 vp_p.n9814 vp_p.n9813 0.006
R22261 vp_p.n9803 vp_p.n9802 0.006
R22262 vp_p.n9800 vp_p.n9799 0.006
R22263 vp_p.n9789 vp_p.n9788 0.006
R22264 vp_p.n9786 vp_p.n9785 0.006
R22265 vp_p.n9775 vp_p.n9774 0.006
R22266 vp_p.n9772 vp_p.n9771 0.006
R22267 vp_p.n9761 vp_p.n9760 0.006
R22268 vp_p.n9758 vp_p.n9757 0.006
R22269 vp_p.n9747 vp_p.n9746 0.006
R22270 vp_p.n9744 vp_p.n9743 0.006
R22271 vp_p.n9733 vp_p.n9732 0.006
R22272 vp_p.n9730 vp_p.n9729 0.006
R22273 vp_p.n9719 vp_p.n9718 0.006
R22274 vp_p.n9716 vp_p.n9715 0.006
R22275 vp_p.n9705 vp_p.n9704 0.006
R22276 vp_p.n9702 vp_p.n9701 0.006
R22277 vp_p.n9691 vp_p.n9690 0.006
R22278 vp_p.n9688 vp_p.n9687 0.006
R22279 vp_p.n9677 vp_p.n9676 0.006
R22280 vp_p.n9674 vp_p.n9673 0.006
R22281 vp_p.n9663 vp_p.n9662 0.006
R22282 vp_p.n9660 vp_p.n9659 0.006
R22283 vp_p.n9649 vp_p.n9648 0.006
R22284 vp_p.n9646 vp_p.n9645 0.006
R22285 vp_p.n9635 vp_p.n9634 0.006
R22286 vp_p.n9632 vp_p.n9631 0.006
R22287 vp_p.n9621 vp_p.n9620 0.006
R22288 vp_p.n9618 vp_p.n9617 0.006
R22289 vp_p.n9607 vp_p.n9606 0.006
R22290 vp_p.n9604 vp_p.n9603 0.006
R22291 vp_p.n9593 vp_p.n9592 0.006
R22292 vp_p.n9590 vp_p.n9589 0.006
R22293 vp_p.n9579 vp_p.n9578 0.006
R22294 vp_p.n9576 vp_p.n9575 0.006
R22295 vp_p.n9565 vp_p.n9564 0.006
R22296 vp_p.n9562 vp_p.n9561 0.006
R22297 vp_p.n9551 vp_p.n9550 0.006
R22298 vp_p.n9548 vp_p.n9547 0.006
R22299 vp_p.n9537 vp_p.n9536 0.006
R22300 vp_p.n9534 vp_p.n9533 0.006
R22301 vp_p.n9523 vp_p.n9522 0.006
R22302 vp_p.n9520 vp_p.n9519 0.006
R22303 vp_p.n9509 vp_p.n9508 0.006
R22304 vp_p.n9506 vp_p.n9505 0.006
R22305 vp_p.n9495 vp_p.n9494 0.006
R22306 vp_p.n9492 vp_p.n9491 0.006
R22307 vp_p.n9481 vp_p.n9480 0.006
R22308 vp_p.n9478 vp_p.n9477 0.006
R22309 vp_p.n9467 vp_p.n9466 0.006
R22310 vp_p.n9464 vp_p.n9463 0.006
R22311 vp_p.n9453 vp_p.n9452 0.006
R22312 vp_p.n9450 vp_p.n9449 0.006
R22313 vp_p.n9439 vp_p.n9438 0.006
R22314 vp_p.n9436 vp_p.n9435 0.006
R22315 vp_p.n9425 vp_p.n9424 0.006
R22316 vp_p.n9422 vp_p.n9421 0.006
R22317 vp_p.n9411 vp_p.n9410 0.006
R22318 vp_p.n9408 vp_p.n9407 0.006
R22319 vp_p.n9397 vp_p.n9396 0.006
R22320 vp_p.n9394 vp_p.n9393 0.006
R22321 vp_p.n9383 vp_p.n9382 0.006
R22322 vp_p.n9380 vp_p.n9379 0.006
R22323 vp_p.n9369 vp_p.n9368 0.006
R22324 vp_p.n9366 vp_p.n9365 0.006
R22325 vp_p.n9355 vp_p.n9354 0.006
R22326 vp_p.n9352 vp_p.n9351 0.006
R22327 vp_p.n9341 vp_p.n9340 0.006
R22328 vp_p.n9338 vp_p.n9337 0.006
R22329 vp_p.n9327 vp_p.n9326 0.006
R22330 vp_p.n9324 vp_p.n9323 0.006
R22331 vp_p.n9313 vp_p.n9312 0.006
R22332 vp_p.n9310 vp_p.n9309 0.006
R22333 vp_p.n9299 vp_p.n9298 0.006
R22334 vp_p.n9296 vp_p.n9295 0.006
R22335 vp_p.n9285 vp_p.n9284 0.006
R22336 vp_p.n9282 vp_p.n9281 0.006
R22337 vp_p.n9271 vp_p.n9270 0.006
R22338 vp_p.n9268 vp_p.n9267 0.006
R22339 vp_p.n9257 vp_p.n9256 0.006
R22340 vp_p.n9254 vp_p.n9253 0.006
R22341 vp_p.n9243 vp_p.n9242 0.006
R22342 vp_p.n9240 vp_p.n9239 0.006
R22343 vp_p.n9229 vp_p.n9228 0.006
R22344 vp_p.n9226 vp_p.n9225 0.006
R22345 vp_p.n9215 vp_p.n9214 0.006
R22346 vp_p.n10167 vp_p.n10166 0.006
R22347 vp_p.n11606 vp_p.n11605 0.006
R22348 vp_p.n13040 vp_p.n13039 0.006
R22349 vp_p.n14409 vp_p.n14408 0.006
R22350 vp_p.n15842 vp_p.n15841 0.006
R22351 vp_p.n17274 vp_p.n17273 0.006
R22352 vp_p.n17738 vp_p.n17737 0.006
R22353 vp_p.n17743 vp_p.n17742 0.006
R22354 vp_p.n17754 vp_p.n17748 0.006
R22355 vp_p.n17758 vp_p.n17757 0.006
R22356 vp_p.n17768 vp_p.n17762 0.006
R22357 vp_p.n17772 vp_p.n17771 0.006
R22358 vp_p.n17782 vp_p.n17776 0.006
R22359 vp_p.n17786 vp_p.n17785 0.006
R22360 vp_p.n17796 vp_p.n17790 0.006
R22361 vp_p.n17800 vp_p.n17799 0.006
R22362 vp_p.n17810 vp_p.n17804 0.006
R22363 vp_p.n17814 vp_p.n17813 0.006
R22364 vp_p.n17824 vp_p.n17818 0.006
R22365 vp_p.n17828 vp_p.n17827 0.006
R22366 vp_p.n17838 vp_p.n17832 0.006
R22367 vp_p.n17842 vp_p.n17841 0.006
R22368 vp_p.n17852 vp_p.n17846 0.006
R22369 vp_p.n17856 vp_p.n17855 0.006
R22370 vp_p.n17866 vp_p.n17860 0.006
R22371 vp_p.n17870 vp_p.n17869 0.006
R22372 vp_p.n17880 vp_p.n17874 0.006
R22373 vp_p.n17884 vp_p.n17883 0.006
R22374 vp_p.n17894 vp_p.n17888 0.006
R22375 vp_p.n17898 vp_p.n17897 0.006
R22376 vp_p.n17908 vp_p.n17902 0.006
R22377 vp_p.n17912 vp_p.n17911 0.006
R22378 vp_p.n17922 vp_p.n17916 0.006
R22379 vp_p.n17926 vp_p.n17925 0.006
R22380 vp_p.n17936 vp_p.n17930 0.006
R22381 vp_p.n17940 vp_p.n17939 0.006
R22382 vp_p.n17950 vp_p.n17944 0.006
R22383 vp_p.n17954 vp_p.n17953 0.006
R22384 vp_p.n17964 vp_p.n17958 0.006
R22385 vp_p.n17968 vp_p.n17967 0.006
R22386 vp_p.n17978 vp_p.n17972 0.006
R22387 vp_p.n17982 vp_p.n17981 0.006
R22388 vp_p.n17992 vp_p.n17986 0.006
R22389 vp_p.n17996 vp_p.n17995 0.006
R22390 vp_p.n18006 vp_p.n18000 0.006
R22391 vp_p.n18010 vp_p.n18009 0.006
R22392 vp_p.n18020 vp_p.n18014 0.006
R22393 vp_p.n18024 vp_p.n18023 0.006
R22394 vp_p.n18034 vp_p.n18028 0.006
R22395 vp_p.n18038 vp_p.n18037 0.006
R22396 vp_p.n18048 vp_p.n18042 0.006
R22397 vp_p.n18052 vp_p.n18051 0.006
R22398 vp_p.n18062 vp_p.n18056 0.006
R22399 vp_p.n18066 vp_p.n18065 0.006
R22400 vp_p.n18076 vp_p.n18070 0.006
R22401 vp_p.n18080 vp_p.n18079 0.006
R22402 vp_p.n18090 vp_p.n18084 0.006
R22403 vp_p.n18094 vp_p.n18093 0.006
R22404 vp_p.n18104 vp_p.n18098 0.006
R22405 vp_p.n18108 vp_p.n18107 0.006
R22406 vp_p.n18118 vp_p.n18112 0.006
R22407 vp_p.n18122 vp_p.n18121 0.006
R22408 vp_p.n18132 vp_p.n18126 0.006
R22409 vp_p.n18136 vp_p.n18135 0.006
R22410 vp_p.n18146 vp_p.n18140 0.006
R22411 vp_p.n18150 vp_p.n18149 0.006
R22412 vp_p.n18160 vp_p.n18154 0.006
R22413 vp_p.n18164 vp_p.n18163 0.006
R22414 vp_p.n18174 vp_p.n18168 0.006
R22415 vp_p.n18178 vp_p.n18177 0.006
R22416 vp_p.n18188 vp_p.n18182 0.006
R22417 vp_p.n18192 vp_p.n18191 0.006
R22418 vp_p.n18202 vp_p.n18196 0.006
R22419 vp_p.n18206 vp_p.n18205 0.006
R22420 vp_p.n18216 vp_p.n18210 0.006
R22421 vp_p.n18220 vp_p.n18219 0.006
R22422 vp_p.n18230 vp_p.n18224 0.006
R22423 vp_p.n18234 vp_p.n18233 0.006
R22424 vp_p.n18244 vp_p.n18238 0.006
R22425 vp_p.n18248 vp_p.n18247 0.006
R22426 vp_p.n18258 vp_p.n18252 0.006
R22427 vp_p.n18262 vp_p.n18261 0.006
R22428 vp_p.n18272 vp_p.n18266 0.006
R22429 vp_p.n18276 vp_p.n18275 0.006
R22430 vp_p.n18286 vp_p.n18280 0.006
R22431 vp_p.n18290 vp_p.n18289 0.006
R22432 vp_p.n18300 vp_p.n18294 0.006
R22433 vp_p.n18304 vp_p.n18303 0.006
R22434 vp_p.n18314 vp_p.n18308 0.006
R22435 vp_p.n18318 vp_p.n18317 0.006
R22436 vp_p.n18328 vp_p.n18322 0.006
R22437 vp_p.n18332 vp_p.n18331 0.006
R22438 vp_p.n18342 vp_p.n18336 0.006
R22439 vp_p.n18346 vp_p.n18345 0.006
R22440 vp_p.n18356 vp_p.n18350 0.006
R22441 vp_p.n18360 vp_p.n18359 0.006
R22442 vp_p.n18370 vp_p.n18364 0.006
R22443 vp_p.n18374 vp_p.n18373 0.006
R22444 vp_p.n18384 vp_p.n18378 0.006
R22445 vp_p.n18388 vp_p.n18387 0.006
R22446 vp_p.n18398 vp_p.n18392 0.006
R22447 vp_p.n18402 vp_p.n18401 0.006
R22448 vp_p.n18412 vp_p.n18406 0.006
R22449 vp_p.n18416 vp_p.n18415 0.006
R22450 vp_p.n18426 vp_p.n18420 0.006
R22451 vp_p.n18430 vp_p.n18429 0.006
R22452 vp_p.n18440 vp_p.n18434 0.006
R22453 vp_p.n18444 vp_p.n18443 0.006
R22454 vp_p.n18454 vp_p.n18448 0.006
R22455 vp_p.n18458 vp_p.n18457 0.006
R22456 vp_p.n18468 vp_p.n18462 0.006
R22457 vp_p.n18472 vp_p.n18471 0.006
R22458 vp_p.n18482 vp_p.n18476 0.006
R22459 vp_p.n18486 vp_p.n18485 0.006
R22460 vp_p.n18496 vp_p.n18490 0.006
R22461 vp_p.n18500 vp_p.n18499 0.006
R22462 vp_p.n18510 vp_p.n18504 0.006
R22463 vp_p.n18514 vp_p.n18513 0.006
R22464 vp_p.n18524 vp_p.n18518 0.006
R22465 vp_p.n18528 vp_p.n18527 0.006
R22466 vp_p.n18538 vp_p.n18532 0.006
R22467 vp_p.n18542 vp_p.n18541 0.006
R22468 vp_p.n18552 vp_p.n18546 0.006
R22469 vp_p.n18556 vp_p.n18555 0.006
R22470 vp_p.n18566 vp_p.n18560 0.006
R22471 vp_p.n18570 vp_p.n18569 0.006
R22472 vp_p.n18580 vp_p.n18574 0.006
R22473 vp_p.n18584 vp_p.n18583 0.006
R22474 vp_p.n18594 vp_p.n18588 0.006
R22475 vp_p.n18598 vp_p.n18597 0.006
R22476 vp_p.n18608 vp_p.n18602 0.006
R22477 vp_p.n18612 vp_p.n18611 0.006
R22478 vp_p.n18622 vp_p.n18616 0.006
R22479 vp_p.n18626 vp_p.n18625 0.006
R22480 vp_p.n18636 vp_p.n18630 0.006
R22481 vp_p.n18640 vp_p.n18639 0.006
R22482 vp_p.n18650 vp_p.n18644 0.006
R22483 vp_p.n18654 vp_p.n18653 0.006
R22484 vp_p.n18664 vp_p.n18658 0.006
R22485 vp_p.n18668 vp_p.n18667 0.006
R22486 vp_p.n18678 vp_p.n18672 0.006
R22487 vp_p.n18682 vp_p.n18681 0.006
R22488 vp_p.n18692 vp_p.n18686 0.006
R22489 vp_p.n18696 vp_p.n18695 0.006
R22490 vp_p.n18700 vp_p.n18699 0.006
R22491 vp_p.n18710 vp_p.n18704 0.006
R22492 vp_p.n18714 vp_p.n18713 0.006
R22493 vp_p.n18719 vp_p.n18718 0.006
R22494 vp_p.n18724 vp_p.n18723 0.006
R22495 vp_p.n18729 vp_p.n18728 0.006
R22496 vp_p.n18734 vp_p.n18733 0.006
R22497 vp_p.n18739 vp_p.n18738 0.006
R22498 vp_p.n18744 vp_p.n18743 0.006
R22499 vp_p.n18749 vp_p.n18748 0.006
R22500 vp_p.n18754 vp_p.n18753 0.006
R22501 vp_p.n18759 vp_p.n18758 0.006
R22502 vp_p.n18701 vp_p.n18700 0.006
R22503 vp_p.n18697 vp_p.n18696 0.006
R22504 vp_p.n18686 vp_p.n18685 0.006
R22505 vp_p.n18683 vp_p.n18682 0.006
R22506 vp_p.n18672 vp_p.n18671 0.006
R22507 vp_p.n18669 vp_p.n18668 0.006
R22508 vp_p.n18658 vp_p.n18657 0.006
R22509 vp_p.n18655 vp_p.n18654 0.006
R22510 vp_p.n18644 vp_p.n18643 0.006
R22511 vp_p.n18641 vp_p.n18640 0.006
R22512 vp_p.n18630 vp_p.n18629 0.006
R22513 vp_p.n18627 vp_p.n18626 0.006
R22514 vp_p.n18616 vp_p.n18615 0.006
R22515 vp_p.n18613 vp_p.n18612 0.006
R22516 vp_p.n18602 vp_p.n18601 0.006
R22517 vp_p.n18599 vp_p.n18598 0.006
R22518 vp_p.n18588 vp_p.n18587 0.006
R22519 vp_p.n18585 vp_p.n18584 0.006
R22520 vp_p.n18574 vp_p.n18573 0.006
R22521 vp_p.n18571 vp_p.n18570 0.006
R22522 vp_p.n18560 vp_p.n18559 0.006
R22523 vp_p.n18557 vp_p.n18556 0.006
R22524 vp_p.n18546 vp_p.n18545 0.006
R22525 vp_p.n18543 vp_p.n18542 0.006
R22526 vp_p.n18532 vp_p.n18531 0.006
R22527 vp_p.n18529 vp_p.n18528 0.006
R22528 vp_p.n18518 vp_p.n18517 0.006
R22529 vp_p.n18515 vp_p.n18514 0.006
R22530 vp_p.n18504 vp_p.n18503 0.006
R22531 vp_p.n18501 vp_p.n18500 0.006
R22532 vp_p.n18490 vp_p.n18489 0.006
R22533 vp_p.n18487 vp_p.n18486 0.006
R22534 vp_p.n18476 vp_p.n18475 0.006
R22535 vp_p.n18473 vp_p.n18472 0.006
R22536 vp_p.n18462 vp_p.n18461 0.006
R22537 vp_p.n18459 vp_p.n18458 0.006
R22538 vp_p.n18448 vp_p.n18447 0.006
R22539 vp_p.n18445 vp_p.n18444 0.006
R22540 vp_p.n18434 vp_p.n18433 0.006
R22541 vp_p.n18431 vp_p.n18430 0.006
R22542 vp_p.n18420 vp_p.n18419 0.006
R22543 vp_p.n18417 vp_p.n18416 0.006
R22544 vp_p.n18406 vp_p.n18405 0.006
R22545 vp_p.n18403 vp_p.n18402 0.006
R22546 vp_p.n18392 vp_p.n18391 0.006
R22547 vp_p.n18389 vp_p.n18388 0.006
R22548 vp_p.n18378 vp_p.n18377 0.006
R22549 vp_p.n18375 vp_p.n18374 0.006
R22550 vp_p.n18364 vp_p.n18363 0.006
R22551 vp_p.n18361 vp_p.n18360 0.006
R22552 vp_p.n18350 vp_p.n18349 0.006
R22553 vp_p.n18347 vp_p.n18346 0.006
R22554 vp_p.n18336 vp_p.n18335 0.006
R22555 vp_p.n18333 vp_p.n18332 0.006
R22556 vp_p.n18322 vp_p.n18321 0.006
R22557 vp_p.n18319 vp_p.n18318 0.006
R22558 vp_p.n18308 vp_p.n18307 0.006
R22559 vp_p.n18305 vp_p.n18304 0.006
R22560 vp_p.n18294 vp_p.n18293 0.006
R22561 vp_p.n18291 vp_p.n18290 0.006
R22562 vp_p.n18280 vp_p.n18279 0.006
R22563 vp_p.n18277 vp_p.n18276 0.006
R22564 vp_p.n18266 vp_p.n18265 0.006
R22565 vp_p.n18263 vp_p.n18262 0.006
R22566 vp_p.n18252 vp_p.n18251 0.006
R22567 vp_p.n18249 vp_p.n18248 0.006
R22568 vp_p.n18238 vp_p.n18237 0.006
R22569 vp_p.n18235 vp_p.n18234 0.006
R22570 vp_p.n18224 vp_p.n18223 0.006
R22571 vp_p.n18221 vp_p.n18220 0.006
R22572 vp_p.n18210 vp_p.n18209 0.006
R22573 vp_p.n18207 vp_p.n18206 0.006
R22574 vp_p.n18196 vp_p.n18195 0.006
R22575 vp_p.n18193 vp_p.n18192 0.006
R22576 vp_p.n18182 vp_p.n18181 0.006
R22577 vp_p.n18179 vp_p.n18178 0.006
R22578 vp_p.n18168 vp_p.n18167 0.006
R22579 vp_p.n18165 vp_p.n18164 0.006
R22580 vp_p.n18154 vp_p.n18153 0.006
R22581 vp_p.n18151 vp_p.n18150 0.006
R22582 vp_p.n18140 vp_p.n18139 0.006
R22583 vp_p.n18137 vp_p.n18136 0.006
R22584 vp_p.n18126 vp_p.n18125 0.006
R22585 vp_p.n18123 vp_p.n18122 0.006
R22586 vp_p.n18112 vp_p.n18111 0.006
R22587 vp_p.n18109 vp_p.n18108 0.006
R22588 vp_p.n18098 vp_p.n18097 0.006
R22589 vp_p.n18095 vp_p.n18094 0.006
R22590 vp_p.n18084 vp_p.n18083 0.006
R22591 vp_p.n18081 vp_p.n18080 0.006
R22592 vp_p.n18070 vp_p.n18069 0.006
R22593 vp_p.n18067 vp_p.n18066 0.006
R22594 vp_p.n18056 vp_p.n18055 0.006
R22595 vp_p.n18053 vp_p.n18052 0.006
R22596 vp_p.n18042 vp_p.n18041 0.006
R22597 vp_p.n18039 vp_p.n18038 0.006
R22598 vp_p.n18028 vp_p.n18027 0.006
R22599 vp_p.n18025 vp_p.n18024 0.006
R22600 vp_p.n18014 vp_p.n18013 0.006
R22601 vp_p.n18011 vp_p.n18010 0.006
R22602 vp_p.n18000 vp_p.n17999 0.006
R22603 vp_p.n17997 vp_p.n17996 0.006
R22604 vp_p.n17986 vp_p.n17985 0.006
R22605 vp_p.n17983 vp_p.n17982 0.006
R22606 vp_p.n17972 vp_p.n17971 0.006
R22607 vp_p.n17969 vp_p.n17968 0.006
R22608 vp_p.n17958 vp_p.n17957 0.006
R22609 vp_p.n17955 vp_p.n17954 0.006
R22610 vp_p.n17944 vp_p.n17943 0.006
R22611 vp_p.n17941 vp_p.n17940 0.006
R22612 vp_p.n17930 vp_p.n17929 0.006
R22613 vp_p.n17927 vp_p.n17926 0.006
R22614 vp_p.n17916 vp_p.n17915 0.006
R22615 vp_p.n17913 vp_p.n17912 0.006
R22616 vp_p.n17902 vp_p.n17901 0.006
R22617 vp_p.n17899 vp_p.n17898 0.006
R22618 vp_p.n17888 vp_p.n17887 0.006
R22619 vp_p.n17885 vp_p.n17884 0.006
R22620 vp_p.n17874 vp_p.n17873 0.006
R22621 vp_p.n17871 vp_p.n17870 0.006
R22622 vp_p.n17860 vp_p.n17859 0.006
R22623 vp_p.n17857 vp_p.n17856 0.006
R22624 vp_p.n17846 vp_p.n17845 0.006
R22625 vp_p.n17843 vp_p.n17842 0.006
R22626 vp_p.n17832 vp_p.n17831 0.006
R22627 vp_p.n17829 vp_p.n17828 0.006
R22628 vp_p.n17818 vp_p.n17817 0.006
R22629 vp_p.n17815 vp_p.n17814 0.006
R22630 vp_p.n17804 vp_p.n17803 0.006
R22631 vp_p.n17801 vp_p.n17800 0.006
R22632 vp_p.n17790 vp_p.n17789 0.006
R22633 vp_p.n17787 vp_p.n17786 0.006
R22634 vp_p.n17776 vp_p.n17775 0.006
R22635 vp_p.n17773 vp_p.n17772 0.006
R22636 vp_p.n17762 vp_p.n17761 0.006
R22637 vp_p.n17759 vp_p.n17758 0.006
R22638 vp_p.n17748 vp_p.n17747 0.006
R22639 vp_p.n18704 vp_p.n18703 0.006
R22640 vp_p.n17279 vp_p.n17278 0.006
R22641 vp_p.n15847 vp_p.n15846 0.006
R22642 vp_p.n14414 vp_p.n14413 0.006
R22643 vp_p.n13045 vp_p.n13044 0.006
R22644 vp_p.n11611 vp_p.n11610 0.006
R22645 vp_p.n10178 vp_p.n10177 0.006
R22646 vp_p.n459 vp_p.n458 0.006
R22647 vp_p.n464 vp_p.n463 0.006
R22648 vp_p.n475 vp_p.n469 0.006
R22649 vp_p.n479 vp_p.n478 0.006
R22650 vp_p.n489 vp_p.n483 0.006
R22651 vp_p.n493 vp_p.n492 0.006
R22652 vp_p.n503 vp_p.n497 0.006
R22653 vp_p.n507 vp_p.n506 0.006
R22654 vp_p.n517 vp_p.n511 0.006
R22655 vp_p.n521 vp_p.n520 0.006
R22656 vp_p.n531 vp_p.n525 0.006
R22657 vp_p.n535 vp_p.n534 0.006
R22658 vp_p.n545 vp_p.n539 0.006
R22659 vp_p.n549 vp_p.n548 0.006
R22660 vp_p.n559 vp_p.n553 0.006
R22661 vp_p.n563 vp_p.n562 0.006
R22662 vp_p.n573 vp_p.n567 0.006
R22663 vp_p.n577 vp_p.n576 0.006
R22664 vp_p.n587 vp_p.n581 0.006
R22665 vp_p.n591 vp_p.n590 0.006
R22666 vp_p.n601 vp_p.n595 0.006
R22667 vp_p.n605 vp_p.n604 0.006
R22668 vp_p.n615 vp_p.n609 0.006
R22669 vp_p.n619 vp_p.n618 0.006
R22670 vp_p.n629 vp_p.n623 0.006
R22671 vp_p.n633 vp_p.n632 0.006
R22672 vp_p.n643 vp_p.n637 0.006
R22673 vp_p.n647 vp_p.n646 0.006
R22674 vp_p.n657 vp_p.n651 0.006
R22675 vp_p.n661 vp_p.n660 0.006
R22676 vp_p.n671 vp_p.n665 0.006
R22677 vp_p.n675 vp_p.n674 0.006
R22678 vp_p.n685 vp_p.n679 0.006
R22679 vp_p.n689 vp_p.n688 0.006
R22680 vp_p.n699 vp_p.n693 0.006
R22681 vp_p.n703 vp_p.n702 0.006
R22682 vp_p.n713 vp_p.n707 0.006
R22683 vp_p.n717 vp_p.n716 0.006
R22684 vp_p.n727 vp_p.n721 0.006
R22685 vp_p.n731 vp_p.n730 0.006
R22686 vp_p.n741 vp_p.n735 0.006
R22687 vp_p.n745 vp_p.n744 0.006
R22688 vp_p.n755 vp_p.n749 0.006
R22689 vp_p.n759 vp_p.n758 0.006
R22690 vp_p.n769 vp_p.n763 0.006
R22691 vp_p.n773 vp_p.n772 0.006
R22692 vp_p.n783 vp_p.n777 0.006
R22693 vp_p.n787 vp_p.n786 0.006
R22694 vp_p.n797 vp_p.n791 0.006
R22695 vp_p.n801 vp_p.n800 0.006
R22696 vp_p.n811 vp_p.n805 0.006
R22697 vp_p.n815 vp_p.n814 0.006
R22698 vp_p.n825 vp_p.n819 0.006
R22699 vp_p.n829 vp_p.n828 0.006
R22700 vp_p.n839 vp_p.n833 0.006
R22701 vp_p.n843 vp_p.n842 0.006
R22702 vp_p.n853 vp_p.n847 0.006
R22703 vp_p.n857 vp_p.n856 0.006
R22704 vp_p.n867 vp_p.n861 0.006
R22705 vp_p.n871 vp_p.n870 0.006
R22706 vp_p.n881 vp_p.n875 0.006
R22707 vp_p.n885 vp_p.n884 0.006
R22708 vp_p.n895 vp_p.n889 0.006
R22709 vp_p.n899 vp_p.n898 0.006
R22710 vp_p.n909 vp_p.n903 0.006
R22711 vp_p.n913 vp_p.n912 0.006
R22712 vp_p.n923 vp_p.n917 0.006
R22713 vp_p.n927 vp_p.n926 0.006
R22714 vp_p.n937 vp_p.n931 0.006
R22715 vp_p.n941 vp_p.n940 0.006
R22716 vp_p.n951 vp_p.n945 0.006
R22717 vp_p.n955 vp_p.n954 0.006
R22718 vp_p.n965 vp_p.n959 0.006
R22719 vp_p.n969 vp_p.n968 0.006
R22720 vp_p.n979 vp_p.n973 0.006
R22721 vp_p.n983 vp_p.n982 0.006
R22722 vp_p.n993 vp_p.n987 0.006
R22723 vp_p.n997 vp_p.n996 0.006
R22724 vp_p.n1007 vp_p.n1001 0.006
R22725 vp_p.n1011 vp_p.n1010 0.006
R22726 vp_p.n1021 vp_p.n1015 0.006
R22727 vp_p.n1025 vp_p.n1024 0.006
R22728 vp_p.n1035 vp_p.n1029 0.006
R22729 vp_p.n1039 vp_p.n1038 0.006
R22730 vp_p.n1049 vp_p.n1043 0.006
R22731 vp_p.n1053 vp_p.n1052 0.006
R22732 vp_p.n1063 vp_p.n1057 0.006
R22733 vp_p.n1067 vp_p.n1066 0.006
R22734 vp_p.n1077 vp_p.n1071 0.006
R22735 vp_p.n1081 vp_p.n1080 0.006
R22736 vp_p.n1091 vp_p.n1085 0.006
R22737 vp_p.n1095 vp_p.n1094 0.006
R22738 vp_p.n1105 vp_p.n1099 0.006
R22739 vp_p.n1109 vp_p.n1108 0.006
R22740 vp_p.n1119 vp_p.n1113 0.006
R22741 vp_p.n1123 vp_p.n1122 0.006
R22742 vp_p.n1133 vp_p.n1127 0.006
R22743 vp_p.n1137 vp_p.n1136 0.006
R22744 vp_p.n1147 vp_p.n1141 0.006
R22745 vp_p.n1151 vp_p.n1150 0.006
R22746 vp_p.n1161 vp_p.n1155 0.006
R22747 vp_p.n1165 vp_p.n1164 0.006
R22748 vp_p.n1175 vp_p.n1169 0.006
R22749 vp_p.n1179 vp_p.n1178 0.006
R22750 vp_p.n1189 vp_p.n1183 0.006
R22751 vp_p.n1193 vp_p.n1192 0.006
R22752 vp_p.n1203 vp_p.n1197 0.006
R22753 vp_p.n1207 vp_p.n1206 0.006
R22754 vp_p.n1217 vp_p.n1211 0.006
R22755 vp_p.n1221 vp_p.n1220 0.006
R22756 vp_p.n1231 vp_p.n1225 0.006
R22757 vp_p.n1235 vp_p.n1234 0.006
R22758 vp_p.n1245 vp_p.n1239 0.006
R22759 vp_p.n1249 vp_p.n1248 0.006
R22760 vp_p.n1259 vp_p.n1253 0.006
R22761 vp_p.n1263 vp_p.n1262 0.006
R22762 vp_p.n1273 vp_p.n1267 0.006
R22763 vp_p.n1277 vp_p.n1276 0.006
R22764 vp_p.n1287 vp_p.n1281 0.006
R22765 vp_p.n1291 vp_p.n1290 0.006
R22766 vp_p.n1301 vp_p.n1295 0.006
R22767 vp_p.n1305 vp_p.n1304 0.006
R22768 vp_p.n1315 vp_p.n1309 0.006
R22769 vp_p.n1319 vp_p.n1318 0.006
R22770 vp_p.n1329 vp_p.n1323 0.006
R22771 vp_p.n1333 vp_p.n1332 0.006
R22772 vp_p.n1343 vp_p.n1337 0.006
R22773 vp_p.n1347 vp_p.n1346 0.006
R22774 vp_p.n1357 vp_p.n1351 0.006
R22775 vp_p.n1361 vp_p.n1360 0.006
R22776 vp_p.n1371 vp_p.n1365 0.006
R22777 vp_p.n1375 vp_p.n1374 0.006
R22778 vp_p.n1385 vp_p.n1379 0.006
R22779 vp_p.n1389 vp_p.n1388 0.006
R22780 vp_p.n1399 vp_p.n1393 0.006
R22781 vp_p.n1403 vp_p.n1402 0.006
R22782 vp_p.n1413 vp_p.n1407 0.006
R22783 vp_p.n1417 vp_p.n1416 0.006
R22784 vp_p.n1427 vp_p.n1421 0.006
R22785 vp_p.n1431 vp_p.n1430 0.006
R22786 vp_p.n1441 vp_p.n1435 0.006
R22787 vp_p.n1445 vp_p.n1444 0.006
R22788 vp_p.n1450 vp_p.n1449 0.006
R22789 vp_p.n1455 vp_p.n1454 0.006
R22790 vp_p.n1460 vp_p.n1459 0.006
R22791 vp_p.n1465 vp_p.n1464 0.006
R22792 vp_p.n1470 vp_p.n1469 0.006
R22793 vp_p.n1475 vp_p.n1474 0.006
R22794 vp_p.n1480 vp_p.n1479 0.006
R22795 vp_p.n1485 vp_p.n1484 0.006
R22796 vp_p.n1432 vp_p.n1431 0.006
R22797 vp_p.n1421 vp_p.n1420 0.006
R22798 vp_p.n1418 vp_p.n1417 0.006
R22799 vp_p.n1407 vp_p.n1406 0.006
R22800 vp_p.n1404 vp_p.n1403 0.006
R22801 vp_p.n1393 vp_p.n1392 0.006
R22802 vp_p.n1390 vp_p.n1389 0.006
R22803 vp_p.n1379 vp_p.n1378 0.006
R22804 vp_p.n1376 vp_p.n1375 0.006
R22805 vp_p.n1365 vp_p.n1364 0.006
R22806 vp_p.n1362 vp_p.n1361 0.006
R22807 vp_p.n1351 vp_p.n1350 0.006
R22808 vp_p.n1348 vp_p.n1347 0.006
R22809 vp_p.n1337 vp_p.n1336 0.006
R22810 vp_p.n1334 vp_p.n1333 0.006
R22811 vp_p.n1323 vp_p.n1322 0.006
R22812 vp_p.n1320 vp_p.n1319 0.006
R22813 vp_p.n1309 vp_p.n1308 0.006
R22814 vp_p.n1306 vp_p.n1305 0.006
R22815 vp_p.n1295 vp_p.n1294 0.006
R22816 vp_p.n1292 vp_p.n1291 0.006
R22817 vp_p.n1281 vp_p.n1280 0.006
R22818 vp_p.n1278 vp_p.n1277 0.006
R22819 vp_p.n1267 vp_p.n1266 0.006
R22820 vp_p.n1264 vp_p.n1263 0.006
R22821 vp_p.n1253 vp_p.n1252 0.006
R22822 vp_p.n1250 vp_p.n1249 0.006
R22823 vp_p.n1239 vp_p.n1238 0.006
R22824 vp_p.n1236 vp_p.n1235 0.006
R22825 vp_p.n1225 vp_p.n1224 0.006
R22826 vp_p.n1222 vp_p.n1221 0.006
R22827 vp_p.n1211 vp_p.n1210 0.006
R22828 vp_p.n1208 vp_p.n1207 0.006
R22829 vp_p.n1197 vp_p.n1196 0.006
R22830 vp_p.n1194 vp_p.n1193 0.006
R22831 vp_p.n1183 vp_p.n1182 0.006
R22832 vp_p.n1180 vp_p.n1179 0.006
R22833 vp_p.n1169 vp_p.n1168 0.006
R22834 vp_p.n1166 vp_p.n1165 0.006
R22835 vp_p.n1155 vp_p.n1154 0.006
R22836 vp_p.n1152 vp_p.n1151 0.006
R22837 vp_p.n1141 vp_p.n1140 0.006
R22838 vp_p.n1138 vp_p.n1137 0.006
R22839 vp_p.n1127 vp_p.n1126 0.006
R22840 vp_p.n1124 vp_p.n1123 0.006
R22841 vp_p.n1113 vp_p.n1112 0.006
R22842 vp_p.n1110 vp_p.n1109 0.006
R22843 vp_p.n1099 vp_p.n1098 0.006
R22844 vp_p.n1096 vp_p.n1095 0.006
R22845 vp_p.n1085 vp_p.n1084 0.006
R22846 vp_p.n1082 vp_p.n1081 0.006
R22847 vp_p.n1071 vp_p.n1070 0.006
R22848 vp_p.n1068 vp_p.n1067 0.006
R22849 vp_p.n1057 vp_p.n1056 0.006
R22850 vp_p.n1054 vp_p.n1053 0.006
R22851 vp_p.n1043 vp_p.n1042 0.006
R22852 vp_p.n1040 vp_p.n1039 0.006
R22853 vp_p.n1029 vp_p.n1028 0.006
R22854 vp_p.n1026 vp_p.n1025 0.006
R22855 vp_p.n1015 vp_p.n1014 0.006
R22856 vp_p.n1012 vp_p.n1011 0.006
R22857 vp_p.n1001 vp_p.n1000 0.006
R22858 vp_p.n998 vp_p.n997 0.006
R22859 vp_p.n987 vp_p.n986 0.006
R22860 vp_p.n984 vp_p.n983 0.006
R22861 vp_p.n973 vp_p.n972 0.006
R22862 vp_p.n970 vp_p.n969 0.006
R22863 vp_p.n959 vp_p.n958 0.006
R22864 vp_p.n956 vp_p.n955 0.006
R22865 vp_p.n945 vp_p.n944 0.006
R22866 vp_p.n942 vp_p.n941 0.006
R22867 vp_p.n931 vp_p.n930 0.006
R22868 vp_p.n928 vp_p.n927 0.006
R22869 vp_p.n917 vp_p.n916 0.006
R22870 vp_p.n914 vp_p.n913 0.006
R22871 vp_p.n903 vp_p.n902 0.006
R22872 vp_p.n900 vp_p.n899 0.006
R22873 vp_p.n889 vp_p.n888 0.006
R22874 vp_p.n886 vp_p.n885 0.006
R22875 vp_p.n875 vp_p.n874 0.006
R22876 vp_p.n872 vp_p.n871 0.006
R22877 vp_p.n861 vp_p.n860 0.006
R22878 vp_p.n858 vp_p.n857 0.006
R22879 vp_p.n847 vp_p.n846 0.006
R22880 vp_p.n844 vp_p.n843 0.006
R22881 vp_p.n833 vp_p.n832 0.006
R22882 vp_p.n830 vp_p.n829 0.006
R22883 vp_p.n819 vp_p.n818 0.006
R22884 vp_p.n816 vp_p.n815 0.006
R22885 vp_p.n805 vp_p.n804 0.006
R22886 vp_p.n802 vp_p.n801 0.006
R22887 vp_p.n791 vp_p.n790 0.006
R22888 vp_p.n788 vp_p.n787 0.006
R22889 vp_p.n777 vp_p.n776 0.006
R22890 vp_p.n774 vp_p.n773 0.006
R22891 vp_p.n763 vp_p.n762 0.006
R22892 vp_p.n760 vp_p.n759 0.006
R22893 vp_p.n749 vp_p.n748 0.006
R22894 vp_p.n746 vp_p.n745 0.006
R22895 vp_p.n735 vp_p.n734 0.006
R22896 vp_p.n732 vp_p.n731 0.006
R22897 vp_p.n721 vp_p.n720 0.006
R22898 vp_p.n718 vp_p.n717 0.006
R22899 vp_p.n707 vp_p.n706 0.006
R22900 vp_p.n704 vp_p.n703 0.006
R22901 vp_p.n693 vp_p.n692 0.006
R22902 vp_p.n690 vp_p.n689 0.006
R22903 vp_p.n679 vp_p.n678 0.006
R22904 vp_p.n676 vp_p.n675 0.006
R22905 vp_p.n665 vp_p.n664 0.006
R22906 vp_p.n662 vp_p.n661 0.006
R22907 vp_p.n651 vp_p.n650 0.006
R22908 vp_p.n648 vp_p.n647 0.006
R22909 vp_p.n637 vp_p.n636 0.006
R22910 vp_p.n634 vp_p.n633 0.006
R22911 vp_p.n623 vp_p.n622 0.006
R22912 vp_p.n620 vp_p.n619 0.006
R22913 vp_p.n609 vp_p.n608 0.006
R22914 vp_p.n606 vp_p.n605 0.006
R22915 vp_p.n595 vp_p.n594 0.006
R22916 vp_p.n592 vp_p.n591 0.006
R22917 vp_p.n581 vp_p.n580 0.006
R22918 vp_p.n578 vp_p.n577 0.006
R22919 vp_p.n567 vp_p.n566 0.006
R22920 vp_p.n564 vp_p.n563 0.006
R22921 vp_p.n553 vp_p.n552 0.006
R22922 vp_p.n550 vp_p.n549 0.006
R22923 vp_p.n539 vp_p.n538 0.006
R22924 vp_p.n536 vp_p.n535 0.006
R22925 vp_p.n525 vp_p.n524 0.006
R22926 vp_p.n522 vp_p.n521 0.006
R22927 vp_p.n511 vp_p.n510 0.006
R22928 vp_p.n508 vp_p.n507 0.006
R22929 vp_p.n497 vp_p.n496 0.006
R22930 vp_p.n494 vp_p.n493 0.006
R22931 vp_p.n483 vp_p.n482 0.006
R22932 vp_p.n480 vp_p.n479 0.006
R22933 vp_p.n469 vp_p.n468 0.006
R22934 vp_p.n1435 vp_p.n1434 0.006
R22935 vp_p.n10183 vp_p.n10182 0.006
R22936 vp_p.n11616 vp_p.n11615 0.006
R22937 vp_p.n13050 vp_p.n13049 0.006
R22938 vp_p.n14419 vp_p.n14418 0.006
R22939 vp_p.n15852 vp_p.n15851 0.006
R22940 vp_p.n17284 vp_p.n17283 0.006
R22941 vp_p.n18715 vp_p.n18714 0.006
R22942 vp_p.n19164 vp_p.n19163 0.006
R22943 vp_p.n19169 vp_p.n19168 0.006
R22944 vp_p.n19180 vp_p.n19174 0.006
R22945 vp_p.n19184 vp_p.n19183 0.006
R22946 vp_p.n19194 vp_p.n19188 0.006
R22947 vp_p.n19198 vp_p.n19197 0.006
R22948 vp_p.n19208 vp_p.n19202 0.006
R22949 vp_p.n19212 vp_p.n19211 0.006
R22950 vp_p.n19222 vp_p.n19216 0.006
R22951 vp_p.n19226 vp_p.n19225 0.006
R22952 vp_p.n19236 vp_p.n19230 0.006
R22953 vp_p.n19240 vp_p.n19239 0.006
R22954 vp_p.n19250 vp_p.n19244 0.006
R22955 vp_p.n19254 vp_p.n19253 0.006
R22956 vp_p.n19264 vp_p.n19258 0.006
R22957 vp_p.n19268 vp_p.n19267 0.006
R22958 vp_p.n19278 vp_p.n19272 0.006
R22959 vp_p.n19282 vp_p.n19281 0.006
R22960 vp_p.n19292 vp_p.n19286 0.006
R22961 vp_p.n19296 vp_p.n19295 0.006
R22962 vp_p.n19306 vp_p.n19300 0.006
R22963 vp_p.n19310 vp_p.n19309 0.006
R22964 vp_p.n19320 vp_p.n19314 0.006
R22965 vp_p.n19324 vp_p.n19323 0.006
R22966 vp_p.n19334 vp_p.n19328 0.006
R22967 vp_p.n19338 vp_p.n19337 0.006
R22968 vp_p.n19348 vp_p.n19342 0.006
R22969 vp_p.n19352 vp_p.n19351 0.006
R22970 vp_p.n19362 vp_p.n19356 0.006
R22971 vp_p.n19366 vp_p.n19365 0.006
R22972 vp_p.n19376 vp_p.n19370 0.006
R22973 vp_p.n19380 vp_p.n19379 0.006
R22974 vp_p.n19390 vp_p.n19384 0.006
R22975 vp_p.n19394 vp_p.n19393 0.006
R22976 vp_p.n19404 vp_p.n19398 0.006
R22977 vp_p.n19408 vp_p.n19407 0.006
R22978 vp_p.n19418 vp_p.n19412 0.006
R22979 vp_p.n19422 vp_p.n19421 0.006
R22980 vp_p.n19432 vp_p.n19426 0.006
R22981 vp_p.n19436 vp_p.n19435 0.006
R22982 vp_p.n19446 vp_p.n19440 0.006
R22983 vp_p.n19450 vp_p.n19449 0.006
R22984 vp_p.n19460 vp_p.n19454 0.006
R22985 vp_p.n19464 vp_p.n19463 0.006
R22986 vp_p.n19474 vp_p.n19468 0.006
R22987 vp_p.n19478 vp_p.n19477 0.006
R22988 vp_p.n19488 vp_p.n19482 0.006
R22989 vp_p.n19492 vp_p.n19491 0.006
R22990 vp_p.n19502 vp_p.n19496 0.006
R22991 vp_p.n19506 vp_p.n19505 0.006
R22992 vp_p.n19516 vp_p.n19510 0.006
R22993 vp_p.n19520 vp_p.n19519 0.006
R22994 vp_p.n19530 vp_p.n19524 0.006
R22995 vp_p.n19534 vp_p.n19533 0.006
R22996 vp_p.n19544 vp_p.n19538 0.006
R22997 vp_p.n19548 vp_p.n19547 0.006
R22998 vp_p.n19558 vp_p.n19552 0.006
R22999 vp_p.n19562 vp_p.n19561 0.006
R23000 vp_p.n19572 vp_p.n19566 0.006
R23001 vp_p.n19576 vp_p.n19575 0.006
R23002 vp_p.n19586 vp_p.n19580 0.006
R23003 vp_p.n19590 vp_p.n19589 0.006
R23004 vp_p.n19600 vp_p.n19594 0.006
R23005 vp_p.n19604 vp_p.n19603 0.006
R23006 vp_p.n19614 vp_p.n19608 0.006
R23007 vp_p.n19618 vp_p.n19617 0.006
R23008 vp_p.n19628 vp_p.n19622 0.006
R23009 vp_p.n19632 vp_p.n19631 0.006
R23010 vp_p.n19642 vp_p.n19636 0.006
R23011 vp_p.n19646 vp_p.n19645 0.006
R23012 vp_p.n19656 vp_p.n19650 0.006
R23013 vp_p.n19660 vp_p.n19659 0.006
R23014 vp_p.n19670 vp_p.n19664 0.006
R23015 vp_p.n19674 vp_p.n19673 0.006
R23016 vp_p.n19684 vp_p.n19678 0.006
R23017 vp_p.n19688 vp_p.n19687 0.006
R23018 vp_p.n19698 vp_p.n19692 0.006
R23019 vp_p.n19702 vp_p.n19701 0.006
R23020 vp_p.n19712 vp_p.n19706 0.006
R23021 vp_p.n19716 vp_p.n19715 0.006
R23022 vp_p.n19726 vp_p.n19720 0.006
R23023 vp_p.n19730 vp_p.n19729 0.006
R23024 vp_p.n19740 vp_p.n19734 0.006
R23025 vp_p.n19744 vp_p.n19743 0.006
R23026 vp_p.n19754 vp_p.n19748 0.006
R23027 vp_p.n19758 vp_p.n19757 0.006
R23028 vp_p.n19768 vp_p.n19762 0.006
R23029 vp_p.n19772 vp_p.n19771 0.006
R23030 vp_p.n19782 vp_p.n19776 0.006
R23031 vp_p.n19786 vp_p.n19785 0.006
R23032 vp_p.n19796 vp_p.n19790 0.006
R23033 vp_p.n19800 vp_p.n19799 0.006
R23034 vp_p.n19810 vp_p.n19804 0.006
R23035 vp_p.n19814 vp_p.n19813 0.006
R23036 vp_p.n19824 vp_p.n19818 0.006
R23037 vp_p.n19828 vp_p.n19827 0.006
R23038 vp_p.n19838 vp_p.n19832 0.006
R23039 vp_p.n19842 vp_p.n19841 0.006
R23040 vp_p.n19852 vp_p.n19846 0.006
R23041 vp_p.n19856 vp_p.n19855 0.006
R23042 vp_p.n19866 vp_p.n19860 0.006
R23043 vp_p.n19870 vp_p.n19869 0.006
R23044 vp_p.n19880 vp_p.n19874 0.006
R23045 vp_p.n19884 vp_p.n19883 0.006
R23046 vp_p.n19894 vp_p.n19888 0.006
R23047 vp_p.n19898 vp_p.n19897 0.006
R23048 vp_p.n19908 vp_p.n19902 0.006
R23049 vp_p.n19912 vp_p.n19911 0.006
R23050 vp_p.n19922 vp_p.n19916 0.006
R23051 vp_p.n19926 vp_p.n19925 0.006
R23052 vp_p.n19936 vp_p.n19930 0.006
R23053 vp_p.n19940 vp_p.n19939 0.006
R23054 vp_p.n19950 vp_p.n19944 0.006
R23055 vp_p.n19954 vp_p.n19953 0.006
R23056 vp_p.n19964 vp_p.n19958 0.006
R23057 vp_p.n19968 vp_p.n19967 0.006
R23058 vp_p.n19978 vp_p.n19972 0.006
R23059 vp_p.n19982 vp_p.n19981 0.006
R23060 vp_p.n19992 vp_p.n19986 0.006
R23061 vp_p.n19996 vp_p.n19995 0.006
R23062 vp_p.n20006 vp_p.n20000 0.006
R23063 vp_p.n20010 vp_p.n20009 0.006
R23064 vp_p.n20020 vp_p.n20014 0.006
R23065 vp_p.n20024 vp_p.n20023 0.006
R23066 vp_p.n20034 vp_p.n20028 0.006
R23067 vp_p.n20038 vp_p.n20037 0.006
R23068 vp_p.n20048 vp_p.n20042 0.006
R23069 vp_p.n20052 vp_p.n20051 0.006
R23070 vp_p.n20062 vp_p.n20056 0.006
R23071 vp_p.n20066 vp_p.n20065 0.006
R23072 vp_p.n20076 vp_p.n20070 0.006
R23073 vp_p.n20080 vp_p.n20079 0.006
R23074 vp_p.n20090 vp_p.n20084 0.006
R23075 vp_p.n20094 vp_p.n20093 0.006
R23076 vp_p.n20104 vp_p.n20098 0.006
R23077 vp_p.n20108 vp_p.n20107 0.006
R23078 vp_p.n20118 vp_p.n20112 0.006
R23079 vp_p.n20122 vp_p.n20121 0.006
R23080 vp_p.n20132 vp_p.n20126 0.006
R23081 vp_p.n20136 vp_p.n20135 0.006
R23082 vp_p.n20140 vp_p.n20139 0.006
R23083 vp_p.n20150 vp_p.n20144 0.006
R23084 vp_p.n20154 vp_p.n20153 0.006
R23085 vp_p.n20159 vp_p.n20158 0.006
R23086 vp_p.n20164 vp_p.n20163 0.006
R23087 vp_p.n20169 vp_p.n20168 0.006
R23088 vp_p.n20174 vp_p.n20173 0.006
R23089 vp_p.n20179 vp_p.n20178 0.006
R23090 vp_p.n20184 vp_p.n20183 0.006
R23091 vp_p.n20189 vp_p.n20188 0.006
R23092 vp_p.n20141 vp_p.n20140 0.006
R23093 vp_p.n20137 vp_p.n20136 0.006
R23094 vp_p.n20126 vp_p.n20125 0.006
R23095 vp_p.n20123 vp_p.n20122 0.006
R23096 vp_p.n20112 vp_p.n20111 0.006
R23097 vp_p.n20109 vp_p.n20108 0.006
R23098 vp_p.n20098 vp_p.n20097 0.006
R23099 vp_p.n20095 vp_p.n20094 0.006
R23100 vp_p.n20084 vp_p.n20083 0.006
R23101 vp_p.n20081 vp_p.n20080 0.006
R23102 vp_p.n20070 vp_p.n20069 0.006
R23103 vp_p.n20067 vp_p.n20066 0.006
R23104 vp_p.n20056 vp_p.n20055 0.006
R23105 vp_p.n20053 vp_p.n20052 0.006
R23106 vp_p.n20042 vp_p.n20041 0.006
R23107 vp_p.n20039 vp_p.n20038 0.006
R23108 vp_p.n20028 vp_p.n20027 0.006
R23109 vp_p.n20025 vp_p.n20024 0.006
R23110 vp_p.n20014 vp_p.n20013 0.006
R23111 vp_p.n20011 vp_p.n20010 0.006
R23112 vp_p.n20000 vp_p.n19999 0.006
R23113 vp_p.n19997 vp_p.n19996 0.006
R23114 vp_p.n19986 vp_p.n19985 0.006
R23115 vp_p.n19983 vp_p.n19982 0.006
R23116 vp_p.n19972 vp_p.n19971 0.006
R23117 vp_p.n19969 vp_p.n19968 0.006
R23118 vp_p.n19958 vp_p.n19957 0.006
R23119 vp_p.n19955 vp_p.n19954 0.006
R23120 vp_p.n19944 vp_p.n19943 0.006
R23121 vp_p.n19941 vp_p.n19940 0.006
R23122 vp_p.n19930 vp_p.n19929 0.006
R23123 vp_p.n19927 vp_p.n19926 0.006
R23124 vp_p.n19916 vp_p.n19915 0.006
R23125 vp_p.n19913 vp_p.n19912 0.006
R23126 vp_p.n19902 vp_p.n19901 0.006
R23127 vp_p.n19899 vp_p.n19898 0.006
R23128 vp_p.n19888 vp_p.n19887 0.006
R23129 vp_p.n19885 vp_p.n19884 0.006
R23130 vp_p.n19874 vp_p.n19873 0.006
R23131 vp_p.n19871 vp_p.n19870 0.006
R23132 vp_p.n19860 vp_p.n19859 0.006
R23133 vp_p.n19857 vp_p.n19856 0.006
R23134 vp_p.n19846 vp_p.n19845 0.006
R23135 vp_p.n19843 vp_p.n19842 0.006
R23136 vp_p.n19832 vp_p.n19831 0.006
R23137 vp_p.n19829 vp_p.n19828 0.006
R23138 vp_p.n19818 vp_p.n19817 0.006
R23139 vp_p.n19815 vp_p.n19814 0.006
R23140 vp_p.n19804 vp_p.n19803 0.006
R23141 vp_p.n19801 vp_p.n19800 0.006
R23142 vp_p.n19790 vp_p.n19789 0.006
R23143 vp_p.n19787 vp_p.n19786 0.006
R23144 vp_p.n19776 vp_p.n19775 0.006
R23145 vp_p.n19773 vp_p.n19772 0.006
R23146 vp_p.n19762 vp_p.n19761 0.006
R23147 vp_p.n19759 vp_p.n19758 0.006
R23148 vp_p.n19748 vp_p.n19747 0.006
R23149 vp_p.n19745 vp_p.n19744 0.006
R23150 vp_p.n19734 vp_p.n19733 0.006
R23151 vp_p.n19731 vp_p.n19730 0.006
R23152 vp_p.n19720 vp_p.n19719 0.006
R23153 vp_p.n19717 vp_p.n19716 0.006
R23154 vp_p.n19706 vp_p.n19705 0.006
R23155 vp_p.n19703 vp_p.n19702 0.006
R23156 vp_p.n19692 vp_p.n19691 0.006
R23157 vp_p.n19689 vp_p.n19688 0.006
R23158 vp_p.n19678 vp_p.n19677 0.006
R23159 vp_p.n19675 vp_p.n19674 0.006
R23160 vp_p.n19664 vp_p.n19663 0.006
R23161 vp_p.n19661 vp_p.n19660 0.006
R23162 vp_p.n19650 vp_p.n19649 0.006
R23163 vp_p.n19647 vp_p.n19646 0.006
R23164 vp_p.n19636 vp_p.n19635 0.006
R23165 vp_p.n19633 vp_p.n19632 0.006
R23166 vp_p.n19622 vp_p.n19621 0.006
R23167 vp_p.n19619 vp_p.n19618 0.006
R23168 vp_p.n19608 vp_p.n19607 0.006
R23169 vp_p.n19605 vp_p.n19604 0.006
R23170 vp_p.n19594 vp_p.n19593 0.006
R23171 vp_p.n19591 vp_p.n19590 0.006
R23172 vp_p.n19580 vp_p.n19579 0.006
R23173 vp_p.n19577 vp_p.n19576 0.006
R23174 vp_p.n19566 vp_p.n19565 0.006
R23175 vp_p.n19563 vp_p.n19562 0.006
R23176 vp_p.n19552 vp_p.n19551 0.006
R23177 vp_p.n19549 vp_p.n19548 0.006
R23178 vp_p.n19538 vp_p.n19537 0.006
R23179 vp_p.n19535 vp_p.n19534 0.006
R23180 vp_p.n19524 vp_p.n19523 0.006
R23181 vp_p.n19521 vp_p.n19520 0.006
R23182 vp_p.n19510 vp_p.n19509 0.006
R23183 vp_p.n19507 vp_p.n19506 0.006
R23184 vp_p.n19496 vp_p.n19495 0.006
R23185 vp_p.n19493 vp_p.n19492 0.006
R23186 vp_p.n19482 vp_p.n19481 0.006
R23187 vp_p.n19479 vp_p.n19478 0.006
R23188 vp_p.n19468 vp_p.n19467 0.006
R23189 vp_p.n19465 vp_p.n19464 0.006
R23190 vp_p.n19454 vp_p.n19453 0.006
R23191 vp_p.n19451 vp_p.n19450 0.006
R23192 vp_p.n19440 vp_p.n19439 0.006
R23193 vp_p.n19437 vp_p.n19436 0.006
R23194 vp_p.n19426 vp_p.n19425 0.006
R23195 vp_p.n19423 vp_p.n19422 0.006
R23196 vp_p.n19412 vp_p.n19411 0.006
R23197 vp_p.n19409 vp_p.n19408 0.006
R23198 vp_p.n19398 vp_p.n19397 0.006
R23199 vp_p.n19395 vp_p.n19394 0.006
R23200 vp_p.n19384 vp_p.n19383 0.006
R23201 vp_p.n19381 vp_p.n19380 0.006
R23202 vp_p.n19370 vp_p.n19369 0.006
R23203 vp_p.n19367 vp_p.n19366 0.006
R23204 vp_p.n19356 vp_p.n19355 0.006
R23205 vp_p.n19353 vp_p.n19352 0.006
R23206 vp_p.n19342 vp_p.n19341 0.006
R23207 vp_p.n19339 vp_p.n19338 0.006
R23208 vp_p.n19328 vp_p.n19327 0.006
R23209 vp_p.n19325 vp_p.n19324 0.006
R23210 vp_p.n19314 vp_p.n19313 0.006
R23211 vp_p.n19311 vp_p.n19310 0.006
R23212 vp_p.n19300 vp_p.n19299 0.006
R23213 vp_p.n19297 vp_p.n19296 0.006
R23214 vp_p.n19286 vp_p.n19285 0.006
R23215 vp_p.n19283 vp_p.n19282 0.006
R23216 vp_p.n19272 vp_p.n19271 0.006
R23217 vp_p.n19269 vp_p.n19268 0.006
R23218 vp_p.n19258 vp_p.n19257 0.006
R23219 vp_p.n19255 vp_p.n19254 0.006
R23220 vp_p.n19244 vp_p.n19243 0.006
R23221 vp_p.n19241 vp_p.n19240 0.006
R23222 vp_p.n19230 vp_p.n19229 0.006
R23223 vp_p.n19227 vp_p.n19226 0.006
R23224 vp_p.n19216 vp_p.n19215 0.006
R23225 vp_p.n19213 vp_p.n19212 0.006
R23226 vp_p.n19202 vp_p.n19201 0.006
R23227 vp_p.n19199 vp_p.n19198 0.006
R23228 vp_p.n19188 vp_p.n19187 0.006
R23229 vp_p.n19185 vp_p.n19184 0.006
R23230 vp_p.n19174 vp_p.n19173 0.006
R23231 vp_p.n20144 vp_p.n20143 0.006
R23232 vp_p.n18720 vp_p.n18719 0.006
R23233 vp_p.n17289 vp_p.n17288 0.006
R23234 vp_p.n15857 vp_p.n15856 0.006
R23235 vp_p.n14424 vp_p.n14423 0.006
R23236 vp_p.n13055 vp_p.n13054 0.006
R23237 vp_p.n11621 vp_p.n11620 0.006
R23238 vp_p.n10188 vp_p.n10187 0.006
R23239 vp_p.n1446 vp_p.n1445 0.006
R23240 vp_p.n1885 vp_p.n1884 0.006
R23241 vp_p.n1890 vp_p.n1889 0.006
R23242 vp_p.n1901 vp_p.n1895 0.006
R23243 vp_p.n1905 vp_p.n1904 0.006
R23244 vp_p.n1915 vp_p.n1909 0.006
R23245 vp_p.n1919 vp_p.n1918 0.006
R23246 vp_p.n1929 vp_p.n1923 0.006
R23247 vp_p.n1933 vp_p.n1932 0.006
R23248 vp_p.n1943 vp_p.n1937 0.006
R23249 vp_p.n1947 vp_p.n1946 0.006
R23250 vp_p.n1957 vp_p.n1951 0.006
R23251 vp_p.n1961 vp_p.n1960 0.006
R23252 vp_p.n1971 vp_p.n1965 0.006
R23253 vp_p.n1975 vp_p.n1974 0.006
R23254 vp_p.n1985 vp_p.n1979 0.006
R23255 vp_p.n1989 vp_p.n1988 0.006
R23256 vp_p.n1999 vp_p.n1993 0.006
R23257 vp_p.n2003 vp_p.n2002 0.006
R23258 vp_p.n2013 vp_p.n2007 0.006
R23259 vp_p.n2017 vp_p.n2016 0.006
R23260 vp_p.n2027 vp_p.n2021 0.006
R23261 vp_p.n2031 vp_p.n2030 0.006
R23262 vp_p.n2041 vp_p.n2035 0.006
R23263 vp_p.n2045 vp_p.n2044 0.006
R23264 vp_p.n2055 vp_p.n2049 0.006
R23265 vp_p.n2059 vp_p.n2058 0.006
R23266 vp_p.n2069 vp_p.n2063 0.006
R23267 vp_p.n2073 vp_p.n2072 0.006
R23268 vp_p.n2083 vp_p.n2077 0.006
R23269 vp_p.n2087 vp_p.n2086 0.006
R23270 vp_p.n2097 vp_p.n2091 0.006
R23271 vp_p.n2101 vp_p.n2100 0.006
R23272 vp_p.n2111 vp_p.n2105 0.006
R23273 vp_p.n2115 vp_p.n2114 0.006
R23274 vp_p.n2125 vp_p.n2119 0.006
R23275 vp_p.n2129 vp_p.n2128 0.006
R23276 vp_p.n2139 vp_p.n2133 0.006
R23277 vp_p.n2143 vp_p.n2142 0.006
R23278 vp_p.n2153 vp_p.n2147 0.006
R23279 vp_p.n2157 vp_p.n2156 0.006
R23280 vp_p.n2167 vp_p.n2161 0.006
R23281 vp_p.n2171 vp_p.n2170 0.006
R23282 vp_p.n2181 vp_p.n2175 0.006
R23283 vp_p.n2185 vp_p.n2184 0.006
R23284 vp_p.n2195 vp_p.n2189 0.006
R23285 vp_p.n2199 vp_p.n2198 0.006
R23286 vp_p.n2209 vp_p.n2203 0.006
R23287 vp_p.n2213 vp_p.n2212 0.006
R23288 vp_p.n2223 vp_p.n2217 0.006
R23289 vp_p.n2227 vp_p.n2226 0.006
R23290 vp_p.n2237 vp_p.n2231 0.006
R23291 vp_p.n2241 vp_p.n2240 0.006
R23292 vp_p.n2251 vp_p.n2245 0.006
R23293 vp_p.n2255 vp_p.n2254 0.006
R23294 vp_p.n2265 vp_p.n2259 0.006
R23295 vp_p.n2269 vp_p.n2268 0.006
R23296 vp_p.n2279 vp_p.n2273 0.006
R23297 vp_p.n2283 vp_p.n2282 0.006
R23298 vp_p.n2293 vp_p.n2287 0.006
R23299 vp_p.n2297 vp_p.n2296 0.006
R23300 vp_p.n2307 vp_p.n2301 0.006
R23301 vp_p.n2311 vp_p.n2310 0.006
R23302 vp_p.n2321 vp_p.n2315 0.006
R23303 vp_p.n2325 vp_p.n2324 0.006
R23304 vp_p.n2335 vp_p.n2329 0.006
R23305 vp_p.n2339 vp_p.n2338 0.006
R23306 vp_p.n2349 vp_p.n2343 0.006
R23307 vp_p.n2353 vp_p.n2352 0.006
R23308 vp_p.n2363 vp_p.n2357 0.006
R23309 vp_p.n2367 vp_p.n2366 0.006
R23310 vp_p.n2377 vp_p.n2371 0.006
R23311 vp_p.n2381 vp_p.n2380 0.006
R23312 vp_p.n2391 vp_p.n2385 0.006
R23313 vp_p.n2395 vp_p.n2394 0.006
R23314 vp_p.n2405 vp_p.n2399 0.006
R23315 vp_p.n2409 vp_p.n2408 0.006
R23316 vp_p.n2419 vp_p.n2413 0.006
R23317 vp_p.n2423 vp_p.n2422 0.006
R23318 vp_p.n2433 vp_p.n2427 0.006
R23319 vp_p.n2437 vp_p.n2436 0.006
R23320 vp_p.n2447 vp_p.n2441 0.006
R23321 vp_p.n2451 vp_p.n2450 0.006
R23322 vp_p.n2461 vp_p.n2455 0.006
R23323 vp_p.n2465 vp_p.n2464 0.006
R23324 vp_p.n2475 vp_p.n2469 0.006
R23325 vp_p.n2479 vp_p.n2478 0.006
R23326 vp_p.n2489 vp_p.n2483 0.006
R23327 vp_p.n2493 vp_p.n2492 0.006
R23328 vp_p.n2503 vp_p.n2497 0.006
R23329 vp_p.n2507 vp_p.n2506 0.006
R23330 vp_p.n2517 vp_p.n2511 0.006
R23331 vp_p.n2521 vp_p.n2520 0.006
R23332 vp_p.n2531 vp_p.n2525 0.006
R23333 vp_p.n2535 vp_p.n2534 0.006
R23334 vp_p.n2545 vp_p.n2539 0.006
R23335 vp_p.n2549 vp_p.n2548 0.006
R23336 vp_p.n2559 vp_p.n2553 0.006
R23337 vp_p.n2563 vp_p.n2562 0.006
R23338 vp_p.n2573 vp_p.n2567 0.006
R23339 vp_p.n2577 vp_p.n2576 0.006
R23340 vp_p.n2587 vp_p.n2581 0.006
R23341 vp_p.n2591 vp_p.n2590 0.006
R23342 vp_p.n2601 vp_p.n2595 0.006
R23343 vp_p.n2605 vp_p.n2604 0.006
R23344 vp_p.n2615 vp_p.n2609 0.006
R23345 vp_p.n2619 vp_p.n2618 0.006
R23346 vp_p.n2629 vp_p.n2623 0.006
R23347 vp_p.n2633 vp_p.n2632 0.006
R23348 vp_p.n2643 vp_p.n2637 0.006
R23349 vp_p.n2647 vp_p.n2646 0.006
R23350 vp_p.n2657 vp_p.n2651 0.006
R23351 vp_p.n2661 vp_p.n2660 0.006
R23352 vp_p.n2671 vp_p.n2665 0.006
R23353 vp_p.n2675 vp_p.n2674 0.006
R23354 vp_p.n2685 vp_p.n2679 0.006
R23355 vp_p.n2689 vp_p.n2688 0.006
R23356 vp_p.n2699 vp_p.n2693 0.006
R23357 vp_p.n2703 vp_p.n2702 0.006
R23358 vp_p.n2713 vp_p.n2707 0.006
R23359 vp_p.n2717 vp_p.n2716 0.006
R23360 vp_p.n2727 vp_p.n2721 0.006
R23361 vp_p.n2731 vp_p.n2730 0.006
R23362 vp_p.n2741 vp_p.n2735 0.006
R23363 vp_p.n2745 vp_p.n2744 0.006
R23364 vp_p.n2755 vp_p.n2749 0.006
R23365 vp_p.n2759 vp_p.n2758 0.006
R23366 vp_p.n2769 vp_p.n2763 0.006
R23367 vp_p.n2773 vp_p.n2772 0.006
R23368 vp_p.n2783 vp_p.n2777 0.006
R23369 vp_p.n2787 vp_p.n2786 0.006
R23370 vp_p.n2797 vp_p.n2791 0.006
R23371 vp_p.n2801 vp_p.n2800 0.006
R23372 vp_p.n2811 vp_p.n2805 0.006
R23373 vp_p.n2815 vp_p.n2814 0.006
R23374 vp_p.n2825 vp_p.n2819 0.006
R23375 vp_p.n2829 vp_p.n2828 0.006
R23376 vp_p.n2839 vp_p.n2833 0.006
R23377 vp_p.n2843 vp_p.n2842 0.006
R23378 vp_p.n2853 vp_p.n2847 0.006
R23379 vp_p.n2857 vp_p.n2856 0.006
R23380 vp_p.n2867 vp_p.n2861 0.006
R23381 vp_p.n2871 vp_p.n2870 0.006
R23382 vp_p.n2881 vp_p.n2875 0.006
R23383 vp_p.n2885 vp_p.n2884 0.006
R23384 vp_p.n2890 vp_p.n2889 0.006
R23385 vp_p.n2895 vp_p.n2894 0.006
R23386 vp_p.n2900 vp_p.n2899 0.006
R23387 vp_p.n2905 vp_p.n2904 0.006
R23388 vp_p.n2910 vp_p.n2909 0.006
R23389 vp_p.n2915 vp_p.n2914 0.006
R23390 vp_p.n2872 vp_p.n2871 0.006
R23391 vp_p.n2861 vp_p.n2860 0.006
R23392 vp_p.n2858 vp_p.n2857 0.006
R23393 vp_p.n2847 vp_p.n2846 0.006
R23394 vp_p.n2844 vp_p.n2843 0.006
R23395 vp_p.n2833 vp_p.n2832 0.006
R23396 vp_p.n2830 vp_p.n2829 0.006
R23397 vp_p.n2819 vp_p.n2818 0.006
R23398 vp_p.n2816 vp_p.n2815 0.006
R23399 vp_p.n2805 vp_p.n2804 0.006
R23400 vp_p.n2802 vp_p.n2801 0.006
R23401 vp_p.n2791 vp_p.n2790 0.006
R23402 vp_p.n2788 vp_p.n2787 0.006
R23403 vp_p.n2777 vp_p.n2776 0.006
R23404 vp_p.n2774 vp_p.n2773 0.006
R23405 vp_p.n2763 vp_p.n2762 0.006
R23406 vp_p.n2760 vp_p.n2759 0.006
R23407 vp_p.n2749 vp_p.n2748 0.006
R23408 vp_p.n2746 vp_p.n2745 0.006
R23409 vp_p.n2735 vp_p.n2734 0.006
R23410 vp_p.n2732 vp_p.n2731 0.006
R23411 vp_p.n2721 vp_p.n2720 0.006
R23412 vp_p.n2718 vp_p.n2717 0.006
R23413 vp_p.n2707 vp_p.n2706 0.006
R23414 vp_p.n2704 vp_p.n2703 0.006
R23415 vp_p.n2693 vp_p.n2692 0.006
R23416 vp_p.n2690 vp_p.n2689 0.006
R23417 vp_p.n2679 vp_p.n2678 0.006
R23418 vp_p.n2676 vp_p.n2675 0.006
R23419 vp_p.n2665 vp_p.n2664 0.006
R23420 vp_p.n2662 vp_p.n2661 0.006
R23421 vp_p.n2651 vp_p.n2650 0.006
R23422 vp_p.n2648 vp_p.n2647 0.006
R23423 vp_p.n2637 vp_p.n2636 0.006
R23424 vp_p.n2634 vp_p.n2633 0.006
R23425 vp_p.n2623 vp_p.n2622 0.006
R23426 vp_p.n2620 vp_p.n2619 0.006
R23427 vp_p.n2609 vp_p.n2608 0.006
R23428 vp_p.n2606 vp_p.n2605 0.006
R23429 vp_p.n2595 vp_p.n2594 0.006
R23430 vp_p.n2592 vp_p.n2591 0.006
R23431 vp_p.n2581 vp_p.n2580 0.006
R23432 vp_p.n2578 vp_p.n2577 0.006
R23433 vp_p.n2567 vp_p.n2566 0.006
R23434 vp_p.n2564 vp_p.n2563 0.006
R23435 vp_p.n2553 vp_p.n2552 0.006
R23436 vp_p.n2550 vp_p.n2549 0.006
R23437 vp_p.n2539 vp_p.n2538 0.006
R23438 vp_p.n2536 vp_p.n2535 0.006
R23439 vp_p.n2525 vp_p.n2524 0.006
R23440 vp_p.n2522 vp_p.n2521 0.006
R23441 vp_p.n2511 vp_p.n2510 0.006
R23442 vp_p.n2508 vp_p.n2507 0.006
R23443 vp_p.n2497 vp_p.n2496 0.006
R23444 vp_p.n2494 vp_p.n2493 0.006
R23445 vp_p.n2483 vp_p.n2482 0.006
R23446 vp_p.n2480 vp_p.n2479 0.006
R23447 vp_p.n2469 vp_p.n2468 0.006
R23448 vp_p.n2466 vp_p.n2465 0.006
R23449 vp_p.n2455 vp_p.n2454 0.006
R23450 vp_p.n2452 vp_p.n2451 0.006
R23451 vp_p.n2441 vp_p.n2440 0.006
R23452 vp_p.n2438 vp_p.n2437 0.006
R23453 vp_p.n2427 vp_p.n2426 0.006
R23454 vp_p.n2424 vp_p.n2423 0.006
R23455 vp_p.n2413 vp_p.n2412 0.006
R23456 vp_p.n2410 vp_p.n2409 0.006
R23457 vp_p.n2399 vp_p.n2398 0.006
R23458 vp_p.n2396 vp_p.n2395 0.006
R23459 vp_p.n2385 vp_p.n2384 0.006
R23460 vp_p.n2382 vp_p.n2381 0.006
R23461 vp_p.n2371 vp_p.n2370 0.006
R23462 vp_p.n2368 vp_p.n2367 0.006
R23463 vp_p.n2357 vp_p.n2356 0.006
R23464 vp_p.n2354 vp_p.n2353 0.006
R23465 vp_p.n2343 vp_p.n2342 0.006
R23466 vp_p.n2340 vp_p.n2339 0.006
R23467 vp_p.n2329 vp_p.n2328 0.006
R23468 vp_p.n2326 vp_p.n2325 0.006
R23469 vp_p.n2315 vp_p.n2314 0.006
R23470 vp_p.n2312 vp_p.n2311 0.006
R23471 vp_p.n2301 vp_p.n2300 0.006
R23472 vp_p.n2298 vp_p.n2297 0.006
R23473 vp_p.n2287 vp_p.n2286 0.006
R23474 vp_p.n2284 vp_p.n2283 0.006
R23475 vp_p.n2273 vp_p.n2272 0.006
R23476 vp_p.n2270 vp_p.n2269 0.006
R23477 vp_p.n2259 vp_p.n2258 0.006
R23478 vp_p.n2256 vp_p.n2255 0.006
R23479 vp_p.n2245 vp_p.n2244 0.006
R23480 vp_p.n2242 vp_p.n2241 0.006
R23481 vp_p.n2231 vp_p.n2230 0.006
R23482 vp_p.n2228 vp_p.n2227 0.006
R23483 vp_p.n2217 vp_p.n2216 0.006
R23484 vp_p.n2214 vp_p.n2213 0.006
R23485 vp_p.n2203 vp_p.n2202 0.006
R23486 vp_p.n2200 vp_p.n2199 0.006
R23487 vp_p.n2189 vp_p.n2188 0.006
R23488 vp_p.n2186 vp_p.n2185 0.006
R23489 vp_p.n2175 vp_p.n2174 0.006
R23490 vp_p.n2172 vp_p.n2171 0.006
R23491 vp_p.n2161 vp_p.n2160 0.006
R23492 vp_p.n2158 vp_p.n2157 0.006
R23493 vp_p.n2147 vp_p.n2146 0.006
R23494 vp_p.n2144 vp_p.n2143 0.006
R23495 vp_p.n2133 vp_p.n2132 0.006
R23496 vp_p.n2130 vp_p.n2129 0.006
R23497 vp_p.n2119 vp_p.n2118 0.006
R23498 vp_p.n2116 vp_p.n2115 0.006
R23499 vp_p.n2105 vp_p.n2104 0.006
R23500 vp_p.n2102 vp_p.n2101 0.006
R23501 vp_p.n2091 vp_p.n2090 0.006
R23502 vp_p.n2088 vp_p.n2087 0.006
R23503 vp_p.n2077 vp_p.n2076 0.006
R23504 vp_p.n2074 vp_p.n2073 0.006
R23505 vp_p.n2063 vp_p.n2062 0.006
R23506 vp_p.n2060 vp_p.n2059 0.006
R23507 vp_p.n2049 vp_p.n2048 0.006
R23508 vp_p.n2046 vp_p.n2045 0.006
R23509 vp_p.n2035 vp_p.n2034 0.006
R23510 vp_p.n2032 vp_p.n2031 0.006
R23511 vp_p.n2021 vp_p.n2020 0.006
R23512 vp_p.n2018 vp_p.n2017 0.006
R23513 vp_p.n2007 vp_p.n2006 0.006
R23514 vp_p.n2004 vp_p.n2003 0.006
R23515 vp_p.n1993 vp_p.n1992 0.006
R23516 vp_p.n1990 vp_p.n1989 0.006
R23517 vp_p.n1979 vp_p.n1978 0.006
R23518 vp_p.n1976 vp_p.n1975 0.006
R23519 vp_p.n1965 vp_p.n1964 0.006
R23520 vp_p.n1962 vp_p.n1961 0.006
R23521 vp_p.n1951 vp_p.n1950 0.006
R23522 vp_p.n1948 vp_p.n1947 0.006
R23523 vp_p.n1937 vp_p.n1936 0.006
R23524 vp_p.n1934 vp_p.n1933 0.006
R23525 vp_p.n1923 vp_p.n1922 0.006
R23526 vp_p.n1920 vp_p.n1919 0.006
R23527 vp_p.n1909 vp_p.n1908 0.006
R23528 vp_p.n1906 vp_p.n1905 0.006
R23529 vp_p.n1895 vp_p.n1894 0.006
R23530 vp_p.n2875 vp_p.n2874 0.006
R23531 vp_p.n1451 vp_p.n1450 0.006
R23532 vp_p.n10193 vp_p.n10192 0.006
R23533 vp_p.n11626 vp_p.n11625 0.006
R23534 vp_p.n13060 vp_p.n13059 0.006
R23535 vp_p.n14429 vp_p.n14428 0.006
R23536 vp_p.n15862 vp_p.n15861 0.006
R23537 vp_p.n17294 vp_p.n17293 0.006
R23538 vp_p.n18725 vp_p.n18724 0.006
R23539 vp_p.n20155 vp_p.n20154 0.006
R23540 vp_p.n20589 vp_p.n20588 0.006
R23541 vp_p.n20594 vp_p.n20593 0.006
R23542 vp_p.n20605 vp_p.n20599 0.006
R23543 vp_p.n20609 vp_p.n20608 0.006
R23544 vp_p.n20619 vp_p.n20613 0.006
R23545 vp_p.n20623 vp_p.n20622 0.006
R23546 vp_p.n20633 vp_p.n20627 0.006
R23547 vp_p.n20637 vp_p.n20636 0.006
R23548 vp_p.n20647 vp_p.n20641 0.006
R23549 vp_p.n20651 vp_p.n20650 0.006
R23550 vp_p.n20661 vp_p.n20655 0.006
R23551 vp_p.n20665 vp_p.n20664 0.006
R23552 vp_p.n20675 vp_p.n20669 0.006
R23553 vp_p.n20679 vp_p.n20678 0.006
R23554 vp_p.n20689 vp_p.n20683 0.006
R23555 vp_p.n20693 vp_p.n20692 0.006
R23556 vp_p.n20703 vp_p.n20697 0.006
R23557 vp_p.n20707 vp_p.n20706 0.006
R23558 vp_p.n20717 vp_p.n20711 0.006
R23559 vp_p.n20721 vp_p.n20720 0.006
R23560 vp_p.n20731 vp_p.n20725 0.006
R23561 vp_p.n20735 vp_p.n20734 0.006
R23562 vp_p.n20745 vp_p.n20739 0.006
R23563 vp_p.n20749 vp_p.n20748 0.006
R23564 vp_p.n20759 vp_p.n20753 0.006
R23565 vp_p.n20763 vp_p.n20762 0.006
R23566 vp_p.n20773 vp_p.n20767 0.006
R23567 vp_p.n20777 vp_p.n20776 0.006
R23568 vp_p.n20787 vp_p.n20781 0.006
R23569 vp_p.n20791 vp_p.n20790 0.006
R23570 vp_p.n20801 vp_p.n20795 0.006
R23571 vp_p.n20805 vp_p.n20804 0.006
R23572 vp_p.n20815 vp_p.n20809 0.006
R23573 vp_p.n20819 vp_p.n20818 0.006
R23574 vp_p.n20829 vp_p.n20823 0.006
R23575 vp_p.n20833 vp_p.n20832 0.006
R23576 vp_p.n20843 vp_p.n20837 0.006
R23577 vp_p.n20847 vp_p.n20846 0.006
R23578 vp_p.n20857 vp_p.n20851 0.006
R23579 vp_p.n20861 vp_p.n20860 0.006
R23580 vp_p.n20871 vp_p.n20865 0.006
R23581 vp_p.n20875 vp_p.n20874 0.006
R23582 vp_p.n20885 vp_p.n20879 0.006
R23583 vp_p.n20889 vp_p.n20888 0.006
R23584 vp_p.n20899 vp_p.n20893 0.006
R23585 vp_p.n20903 vp_p.n20902 0.006
R23586 vp_p.n20913 vp_p.n20907 0.006
R23587 vp_p.n20917 vp_p.n20916 0.006
R23588 vp_p.n20927 vp_p.n20921 0.006
R23589 vp_p.n20931 vp_p.n20930 0.006
R23590 vp_p.n20941 vp_p.n20935 0.006
R23591 vp_p.n20945 vp_p.n20944 0.006
R23592 vp_p.n20955 vp_p.n20949 0.006
R23593 vp_p.n20959 vp_p.n20958 0.006
R23594 vp_p.n20969 vp_p.n20963 0.006
R23595 vp_p.n20973 vp_p.n20972 0.006
R23596 vp_p.n20983 vp_p.n20977 0.006
R23597 vp_p.n20987 vp_p.n20986 0.006
R23598 vp_p.n20997 vp_p.n20991 0.006
R23599 vp_p.n21001 vp_p.n21000 0.006
R23600 vp_p.n21011 vp_p.n21005 0.006
R23601 vp_p.n21015 vp_p.n21014 0.006
R23602 vp_p.n21025 vp_p.n21019 0.006
R23603 vp_p.n21029 vp_p.n21028 0.006
R23604 vp_p.n21039 vp_p.n21033 0.006
R23605 vp_p.n21043 vp_p.n21042 0.006
R23606 vp_p.n21053 vp_p.n21047 0.006
R23607 vp_p.n21057 vp_p.n21056 0.006
R23608 vp_p.n21067 vp_p.n21061 0.006
R23609 vp_p.n21071 vp_p.n21070 0.006
R23610 vp_p.n21081 vp_p.n21075 0.006
R23611 vp_p.n21085 vp_p.n21084 0.006
R23612 vp_p.n21095 vp_p.n21089 0.006
R23613 vp_p.n21099 vp_p.n21098 0.006
R23614 vp_p.n21109 vp_p.n21103 0.006
R23615 vp_p.n21113 vp_p.n21112 0.006
R23616 vp_p.n21123 vp_p.n21117 0.006
R23617 vp_p.n21127 vp_p.n21126 0.006
R23618 vp_p.n21137 vp_p.n21131 0.006
R23619 vp_p.n21141 vp_p.n21140 0.006
R23620 vp_p.n21151 vp_p.n21145 0.006
R23621 vp_p.n21155 vp_p.n21154 0.006
R23622 vp_p.n21165 vp_p.n21159 0.006
R23623 vp_p.n21169 vp_p.n21168 0.006
R23624 vp_p.n21179 vp_p.n21173 0.006
R23625 vp_p.n21183 vp_p.n21182 0.006
R23626 vp_p.n21193 vp_p.n21187 0.006
R23627 vp_p.n21197 vp_p.n21196 0.006
R23628 vp_p.n21207 vp_p.n21201 0.006
R23629 vp_p.n21211 vp_p.n21210 0.006
R23630 vp_p.n21221 vp_p.n21215 0.006
R23631 vp_p.n21225 vp_p.n21224 0.006
R23632 vp_p.n21235 vp_p.n21229 0.006
R23633 vp_p.n21239 vp_p.n21238 0.006
R23634 vp_p.n21249 vp_p.n21243 0.006
R23635 vp_p.n21253 vp_p.n21252 0.006
R23636 vp_p.n21263 vp_p.n21257 0.006
R23637 vp_p.n21267 vp_p.n21266 0.006
R23638 vp_p.n21277 vp_p.n21271 0.006
R23639 vp_p.n21281 vp_p.n21280 0.006
R23640 vp_p.n21291 vp_p.n21285 0.006
R23641 vp_p.n21295 vp_p.n21294 0.006
R23642 vp_p.n21305 vp_p.n21299 0.006
R23643 vp_p.n21309 vp_p.n21308 0.006
R23644 vp_p.n21319 vp_p.n21313 0.006
R23645 vp_p.n21323 vp_p.n21322 0.006
R23646 vp_p.n21333 vp_p.n21327 0.006
R23647 vp_p.n21337 vp_p.n21336 0.006
R23648 vp_p.n21347 vp_p.n21341 0.006
R23649 vp_p.n21351 vp_p.n21350 0.006
R23650 vp_p.n21361 vp_p.n21355 0.006
R23651 vp_p.n21365 vp_p.n21364 0.006
R23652 vp_p.n21375 vp_p.n21369 0.006
R23653 vp_p.n21379 vp_p.n21378 0.006
R23654 vp_p.n21389 vp_p.n21383 0.006
R23655 vp_p.n21393 vp_p.n21392 0.006
R23656 vp_p.n21403 vp_p.n21397 0.006
R23657 vp_p.n21407 vp_p.n21406 0.006
R23658 vp_p.n21417 vp_p.n21411 0.006
R23659 vp_p.n21421 vp_p.n21420 0.006
R23660 vp_p.n21431 vp_p.n21425 0.006
R23661 vp_p.n21435 vp_p.n21434 0.006
R23662 vp_p.n21445 vp_p.n21439 0.006
R23663 vp_p.n21449 vp_p.n21448 0.006
R23664 vp_p.n21459 vp_p.n21453 0.006
R23665 vp_p.n21463 vp_p.n21462 0.006
R23666 vp_p.n21473 vp_p.n21467 0.006
R23667 vp_p.n21477 vp_p.n21476 0.006
R23668 vp_p.n21487 vp_p.n21481 0.006
R23669 vp_p.n21491 vp_p.n21490 0.006
R23670 vp_p.n21501 vp_p.n21495 0.006
R23671 vp_p.n21505 vp_p.n21504 0.006
R23672 vp_p.n21515 vp_p.n21509 0.006
R23673 vp_p.n21519 vp_p.n21518 0.006
R23674 vp_p.n21529 vp_p.n21523 0.006
R23675 vp_p.n21533 vp_p.n21532 0.006
R23676 vp_p.n21543 vp_p.n21537 0.006
R23677 vp_p.n21547 vp_p.n21546 0.006
R23678 vp_p.n21557 vp_p.n21551 0.006
R23679 vp_p.n21561 vp_p.n21560 0.006
R23680 vp_p.n21571 vp_p.n21565 0.006
R23681 vp_p.n21575 vp_p.n21574 0.006
R23682 vp_p.n21579 vp_p.n21578 0.006
R23683 vp_p.n21589 vp_p.n21583 0.006
R23684 vp_p.n21593 vp_p.n21592 0.006
R23685 vp_p.n21598 vp_p.n21597 0.006
R23686 vp_p.n21603 vp_p.n21602 0.006
R23687 vp_p.n21608 vp_p.n21607 0.006
R23688 vp_p.n21613 vp_p.n21612 0.006
R23689 vp_p.n21618 vp_p.n21617 0.006
R23690 vp_p.n21580 vp_p.n21579 0.006
R23691 vp_p.n21576 vp_p.n21575 0.006
R23692 vp_p.n21565 vp_p.n21564 0.006
R23693 vp_p.n21562 vp_p.n21561 0.006
R23694 vp_p.n21551 vp_p.n21550 0.006
R23695 vp_p.n21548 vp_p.n21547 0.006
R23696 vp_p.n21537 vp_p.n21536 0.006
R23697 vp_p.n21534 vp_p.n21533 0.006
R23698 vp_p.n21523 vp_p.n21522 0.006
R23699 vp_p.n21520 vp_p.n21519 0.006
R23700 vp_p.n21509 vp_p.n21508 0.006
R23701 vp_p.n21506 vp_p.n21505 0.006
R23702 vp_p.n21495 vp_p.n21494 0.006
R23703 vp_p.n21492 vp_p.n21491 0.006
R23704 vp_p.n21481 vp_p.n21480 0.006
R23705 vp_p.n21478 vp_p.n21477 0.006
R23706 vp_p.n21467 vp_p.n21466 0.006
R23707 vp_p.n21464 vp_p.n21463 0.006
R23708 vp_p.n21453 vp_p.n21452 0.006
R23709 vp_p.n21450 vp_p.n21449 0.006
R23710 vp_p.n21439 vp_p.n21438 0.006
R23711 vp_p.n21436 vp_p.n21435 0.006
R23712 vp_p.n21425 vp_p.n21424 0.006
R23713 vp_p.n21422 vp_p.n21421 0.006
R23714 vp_p.n21411 vp_p.n21410 0.006
R23715 vp_p.n21408 vp_p.n21407 0.006
R23716 vp_p.n21397 vp_p.n21396 0.006
R23717 vp_p.n21394 vp_p.n21393 0.006
R23718 vp_p.n21383 vp_p.n21382 0.006
R23719 vp_p.n21380 vp_p.n21379 0.006
R23720 vp_p.n21369 vp_p.n21368 0.006
R23721 vp_p.n21366 vp_p.n21365 0.006
R23722 vp_p.n21355 vp_p.n21354 0.006
R23723 vp_p.n21352 vp_p.n21351 0.006
R23724 vp_p.n21341 vp_p.n21340 0.006
R23725 vp_p.n21338 vp_p.n21337 0.006
R23726 vp_p.n21327 vp_p.n21326 0.006
R23727 vp_p.n21324 vp_p.n21323 0.006
R23728 vp_p.n21313 vp_p.n21312 0.006
R23729 vp_p.n21310 vp_p.n21309 0.006
R23730 vp_p.n21299 vp_p.n21298 0.006
R23731 vp_p.n21296 vp_p.n21295 0.006
R23732 vp_p.n21285 vp_p.n21284 0.006
R23733 vp_p.n21282 vp_p.n21281 0.006
R23734 vp_p.n21271 vp_p.n21270 0.006
R23735 vp_p.n21268 vp_p.n21267 0.006
R23736 vp_p.n21257 vp_p.n21256 0.006
R23737 vp_p.n21254 vp_p.n21253 0.006
R23738 vp_p.n21243 vp_p.n21242 0.006
R23739 vp_p.n21240 vp_p.n21239 0.006
R23740 vp_p.n21229 vp_p.n21228 0.006
R23741 vp_p.n21226 vp_p.n21225 0.006
R23742 vp_p.n21215 vp_p.n21214 0.006
R23743 vp_p.n21212 vp_p.n21211 0.006
R23744 vp_p.n21201 vp_p.n21200 0.006
R23745 vp_p.n21198 vp_p.n21197 0.006
R23746 vp_p.n21187 vp_p.n21186 0.006
R23747 vp_p.n21184 vp_p.n21183 0.006
R23748 vp_p.n21173 vp_p.n21172 0.006
R23749 vp_p.n21170 vp_p.n21169 0.006
R23750 vp_p.n21159 vp_p.n21158 0.006
R23751 vp_p.n21156 vp_p.n21155 0.006
R23752 vp_p.n21145 vp_p.n21144 0.006
R23753 vp_p.n21142 vp_p.n21141 0.006
R23754 vp_p.n21131 vp_p.n21130 0.006
R23755 vp_p.n21128 vp_p.n21127 0.006
R23756 vp_p.n21117 vp_p.n21116 0.006
R23757 vp_p.n21114 vp_p.n21113 0.006
R23758 vp_p.n21103 vp_p.n21102 0.006
R23759 vp_p.n21100 vp_p.n21099 0.006
R23760 vp_p.n21089 vp_p.n21088 0.006
R23761 vp_p.n21086 vp_p.n21085 0.006
R23762 vp_p.n21075 vp_p.n21074 0.006
R23763 vp_p.n21072 vp_p.n21071 0.006
R23764 vp_p.n21061 vp_p.n21060 0.006
R23765 vp_p.n21058 vp_p.n21057 0.006
R23766 vp_p.n21047 vp_p.n21046 0.006
R23767 vp_p.n21044 vp_p.n21043 0.006
R23768 vp_p.n21033 vp_p.n21032 0.006
R23769 vp_p.n21030 vp_p.n21029 0.006
R23770 vp_p.n21019 vp_p.n21018 0.006
R23771 vp_p.n21016 vp_p.n21015 0.006
R23772 vp_p.n21005 vp_p.n21004 0.006
R23773 vp_p.n21002 vp_p.n21001 0.006
R23774 vp_p.n20991 vp_p.n20990 0.006
R23775 vp_p.n20988 vp_p.n20987 0.006
R23776 vp_p.n20977 vp_p.n20976 0.006
R23777 vp_p.n20974 vp_p.n20973 0.006
R23778 vp_p.n20963 vp_p.n20962 0.006
R23779 vp_p.n20960 vp_p.n20959 0.006
R23780 vp_p.n20949 vp_p.n20948 0.006
R23781 vp_p.n20946 vp_p.n20945 0.006
R23782 vp_p.n20935 vp_p.n20934 0.006
R23783 vp_p.n20932 vp_p.n20931 0.006
R23784 vp_p.n20921 vp_p.n20920 0.006
R23785 vp_p.n20918 vp_p.n20917 0.006
R23786 vp_p.n20907 vp_p.n20906 0.006
R23787 vp_p.n20904 vp_p.n20903 0.006
R23788 vp_p.n20893 vp_p.n20892 0.006
R23789 vp_p.n20890 vp_p.n20889 0.006
R23790 vp_p.n20879 vp_p.n20878 0.006
R23791 vp_p.n20876 vp_p.n20875 0.006
R23792 vp_p.n20865 vp_p.n20864 0.006
R23793 vp_p.n20862 vp_p.n20861 0.006
R23794 vp_p.n20851 vp_p.n20850 0.006
R23795 vp_p.n20848 vp_p.n20847 0.006
R23796 vp_p.n20837 vp_p.n20836 0.006
R23797 vp_p.n20834 vp_p.n20833 0.006
R23798 vp_p.n20823 vp_p.n20822 0.006
R23799 vp_p.n20820 vp_p.n20819 0.006
R23800 vp_p.n20809 vp_p.n20808 0.006
R23801 vp_p.n20806 vp_p.n20805 0.006
R23802 vp_p.n20795 vp_p.n20794 0.006
R23803 vp_p.n20792 vp_p.n20791 0.006
R23804 vp_p.n20781 vp_p.n20780 0.006
R23805 vp_p.n20778 vp_p.n20777 0.006
R23806 vp_p.n20767 vp_p.n20766 0.006
R23807 vp_p.n20764 vp_p.n20763 0.006
R23808 vp_p.n20753 vp_p.n20752 0.006
R23809 vp_p.n20750 vp_p.n20749 0.006
R23810 vp_p.n20739 vp_p.n20738 0.006
R23811 vp_p.n20736 vp_p.n20735 0.006
R23812 vp_p.n20725 vp_p.n20724 0.006
R23813 vp_p.n20722 vp_p.n20721 0.006
R23814 vp_p.n20711 vp_p.n20710 0.006
R23815 vp_p.n20708 vp_p.n20707 0.006
R23816 vp_p.n20697 vp_p.n20696 0.006
R23817 vp_p.n20694 vp_p.n20693 0.006
R23818 vp_p.n20683 vp_p.n20682 0.006
R23819 vp_p.n20680 vp_p.n20679 0.006
R23820 vp_p.n20669 vp_p.n20668 0.006
R23821 vp_p.n20666 vp_p.n20665 0.006
R23822 vp_p.n20655 vp_p.n20654 0.006
R23823 vp_p.n20652 vp_p.n20651 0.006
R23824 vp_p.n20641 vp_p.n20640 0.006
R23825 vp_p.n20638 vp_p.n20637 0.006
R23826 vp_p.n20627 vp_p.n20626 0.006
R23827 vp_p.n20624 vp_p.n20623 0.006
R23828 vp_p.n20613 vp_p.n20612 0.006
R23829 vp_p.n20610 vp_p.n20609 0.006
R23830 vp_p.n20599 vp_p.n20598 0.006
R23831 vp_p.n21583 vp_p.n21582 0.006
R23832 vp_p.n20160 vp_p.n20159 0.006
R23833 vp_p.n18730 vp_p.n18729 0.006
R23834 vp_p.n17299 vp_p.n17298 0.006
R23835 vp_p.n15867 vp_p.n15866 0.006
R23836 vp_p.n14434 vp_p.n14433 0.006
R23837 vp_p.n13065 vp_p.n13064 0.006
R23838 vp_p.n11631 vp_p.n11630 0.006
R23839 vp_p.n10198 vp_p.n10197 0.006
R23840 vp_p.n1456 vp_p.n1455 0.006
R23841 vp_p.n2886 vp_p.n2885 0.006
R23842 vp_p.n3310 vp_p.n3309 0.006
R23843 vp_p.n3315 vp_p.n3314 0.006
R23844 vp_p.n3326 vp_p.n3320 0.006
R23845 vp_p.n3330 vp_p.n3329 0.006
R23846 vp_p.n3340 vp_p.n3334 0.006
R23847 vp_p.n3344 vp_p.n3343 0.006
R23848 vp_p.n3354 vp_p.n3348 0.006
R23849 vp_p.n3358 vp_p.n3357 0.006
R23850 vp_p.n3368 vp_p.n3362 0.006
R23851 vp_p.n3372 vp_p.n3371 0.006
R23852 vp_p.n3382 vp_p.n3376 0.006
R23853 vp_p.n3386 vp_p.n3385 0.006
R23854 vp_p.n3396 vp_p.n3390 0.006
R23855 vp_p.n3400 vp_p.n3399 0.006
R23856 vp_p.n3410 vp_p.n3404 0.006
R23857 vp_p.n3414 vp_p.n3413 0.006
R23858 vp_p.n3424 vp_p.n3418 0.006
R23859 vp_p.n3428 vp_p.n3427 0.006
R23860 vp_p.n3438 vp_p.n3432 0.006
R23861 vp_p.n3442 vp_p.n3441 0.006
R23862 vp_p.n3452 vp_p.n3446 0.006
R23863 vp_p.n3456 vp_p.n3455 0.006
R23864 vp_p.n3466 vp_p.n3460 0.006
R23865 vp_p.n3470 vp_p.n3469 0.006
R23866 vp_p.n3480 vp_p.n3474 0.006
R23867 vp_p.n3484 vp_p.n3483 0.006
R23868 vp_p.n3494 vp_p.n3488 0.006
R23869 vp_p.n3498 vp_p.n3497 0.006
R23870 vp_p.n3508 vp_p.n3502 0.006
R23871 vp_p.n3512 vp_p.n3511 0.006
R23872 vp_p.n3522 vp_p.n3516 0.006
R23873 vp_p.n3526 vp_p.n3525 0.006
R23874 vp_p.n3536 vp_p.n3530 0.006
R23875 vp_p.n3540 vp_p.n3539 0.006
R23876 vp_p.n3550 vp_p.n3544 0.006
R23877 vp_p.n3554 vp_p.n3553 0.006
R23878 vp_p.n3564 vp_p.n3558 0.006
R23879 vp_p.n3568 vp_p.n3567 0.006
R23880 vp_p.n3578 vp_p.n3572 0.006
R23881 vp_p.n3582 vp_p.n3581 0.006
R23882 vp_p.n3592 vp_p.n3586 0.006
R23883 vp_p.n3596 vp_p.n3595 0.006
R23884 vp_p.n3606 vp_p.n3600 0.006
R23885 vp_p.n3610 vp_p.n3609 0.006
R23886 vp_p.n3620 vp_p.n3614 0.006
R23887 vp_p.n3624 vp_p.n3623 0.006
R23888 vp_p.n3634 vp_p.n3628 0.006
R23889 vp_p.n3638 vp_p.n3637 0.006
R23890 vp_p.n3648 vp_p.n3642 0.006
R23891 vp_p.n3652 vp_p.n3651 0.006
R23892 vp_p.n3662 vp_p.n3656 0.006
R23893 vp_p.n3666 vp_p.n3665 0.006
R23894 vp_p.n3676 vp_p.n3670 0.006
R23895 vp_p.n3680 vp_p.n3679 0.006
R23896 vp_p.n3690 vp_p.n3684 0.006
R23897 vp_p.n3694 vp_p.n3693 0.006
R23898 vp_p.n3704 vp_p.n3698 0.006
R23899 vp_p.n3708 vp_p.n3707 0.006
R23900 vp_p.n3718 vp_p.n3712 0.006
R23901 vp_p.n3722 vp_p.n3721 0.006
R23902 vp_p.n3732 vp_p.n3726 0.006
R23903 vp_p.n3736 vp_p.n3735 0.006
R23904 vp_p.n3746 vp_p.n3740 0.006
R23905 vp_p.n3750 vp_p.n3749 0.006
R23906 vp_p.n3760 vp_p.n3754 0.006
R23907 vp_p.n3764 vp_p.n3763 0.006
R23908 vp_p.n3774 vp_p.n3768 0.006
R23909 vp_p.n3778 vp_p.n3777 0.006
R23910 vp_p.n3788 vp_p.n3782 0.006
R23911 vp_p.n3792 vp_p.n3791 0.006
R23912 vp_p.n3802 vp_p.n3796 0.006
R23913 vp_p.n3806 vp_p.n3805 0.006
R23914 vp_p.n3816 vp_p.n3810 0.006
R23915 vp_p.n3820 vp_p.n3819 0.006
R23916 vp_p.n3830 vp_p.n3824 0.006
R23917 vp_p.n3834 vp_p.n3833 0.006
R23918 vp_p.n3844 vp_p.n3838 0.006
R23919 vp_p.n3848 vp_p.n3847 0.006
R23920 vp_p.n3858 vp_p.n3852 0.006
R23921 vp_p.n3862 vp_p.n3861 0.006
R23922 vp_p.n3872 vp_p.n3866 0.006
R23923 vp_p.n3876 vp_p.n3875 0.006
R23924 vp_p.n3886 vp_p.n3880 0.006
R23925 vp_p.n3890 vp_p.n3889 0.006
R23926 vp_p.n3900 vp_p.n3894 0.006
R23927 vp_p.n3904 vp_p.n3903 0.006
R23928 vp_p.n3914 vp_p.n3908 0.006
R23929 vp_p.n3918 vp_p.n3917 0.006
R23930 vp_p.n3928 vp_p.n3922 0.006
R23931 vp_p.n3932 vp_p.n3931 0.006
R23932 vp_p.n3942 vp_p.n3936 0.006
R23933 vp_p.n3946 vp_p.n3945 0.006
R23934 vp_p.n3956 vp_p.n3950 0.006
R23935 vp_p.n3960 vp_p.n3959 0.006
R23936 vp_p.n3970 vp_p.n3964 0.006
R23937 vp_p.n3974 vp_p.n3973 0.006
R23938 vp_p.n3984 vp_p.n3978 0.006
R23939 vp_p.n3988 vp_p.n3987 0.006
R23940 vp_p.n3998 vp_p.n3992 0.006
R23941 vp_p.n4002 vp_p.n4001 0.006
R23942 vp_p.n4012 vp_p.n4006 0.006
R23943 vp_p.n4016 vp_p.n4015 0.006
R23944 vp_p.n4026 vp_p.n4020 0.006
R23945 vp_p.n4030 vp_p.n4029 0.006
R23946 vp_p.n4040 vp_p.n4034 0.006
R23947 vp_p.n4044 vp_p.n4043 0.006
R23948 vp_p.n4054 vp_p.n4048 0.006
R23949 vp_p.n4058 vp_p.n4057 0.006
R23950 vp_p.n4068 vp_p.n4062 0.006
R23951 vp_p.n4072 vp_p.n4071 0.006
R23952 vp_p.n4082 vp_p.n4076 0.006
R23953 vp_p.n4086 vp_p.n4085 0.006
R23954 vp_p.n4096 vp_p.n4090 0.006
R23955 vp_p.n4100 vp_p.n4099 0.006
R23956 vp_p.n4110 vp_p.n4104 0.006
R23957 vp_p.n4114 vp_p.n4113 0.006
R23958 vp_p.n4124 vp_p.n4118 0.006
R23959 vp_p.n4128 vp_p.n4127 0.006
R23960 vp_p.n4138 vp_p.n4132 0.006
R23961 vp_p.n4142 vp_p.n4141 0.006
R23962 vp_p.n4152 vp_p.n4146 0.006
R23963 vp_p.n4156 vp_p.n4155 0.006
R23964 vp_p.n4166 vp_p.n4160 0.006
R23965 vp_p.n4170 vp_p.n4169 0.006
R23966 vp_p.n4180 vp_p.n4174 0.006
R23967 vp_p.n4184 vp_p.n4183 0.006
R23968 vp_p.n4194 vp_p.n4188 0.006
R23969 vp_p.n4198 vp_p.n4197 0.006
R23970 vp_p.n4208 vp_p.n4202 0.006
R23971 vp_p.n4212 vp_p.n4211 0.006
R23972 vp_p.n4222 vp_p.n4216 0.006
R23973 vp_p.n4226 vp_p.n4225 0.006
R23974 vp_p.n4236 vp_p.n4230 0.006
R23975 vp_p.n4240 vp_p.n4239 0.006
R23976 vp_p.n4250 vp_p.n4244 0.006
R23977 vp_p.n4254 vp_p.n4253 0.006
R23978 vp_p.n4264 vp_p.n4258 0.006
R23979 vp_p.n4268 vp_p.n4267 0.006
R23980 vp_p.n4278 vp_p.n4272 0.006
R23981 vp_p.n4282 vp_p.n4281 0.006
R23982 vp_p.n4292 vp_p.n4286 0.006
R23983 vp_p.n4296 vp_p.n4295 0.006
R23984 vp_p.n4306 vp_p.n4300 0.006
R23985 vp_p.n4310 vp_p.n4309 0.006
R23986 vp_p.n4320 vp_p.n4314 0.006
R23987 vp_p.n4324 vp_p.n4323 0.006
R23988 vp_p.n4329 vp_p.n4328 0.006
R23989 vp_p.n4334 vp_p.n4333 0.006
R23990 vp_p.n4339 vp_p.n4338 0.006
R23991 vp_p.n4344 vp_p.n4343 0.006
R23992 vp_p.n4311 vp_p.n4310 0.006
R23993 vp_p.n4300 vp_p.n4299 0.006
R23994 vp_p.n4297 vp_p.n4296 0.006
R23995 vp_p.n4286 vp_p.n4285 0.006
R23996 vp_p.n4283 vp_p.n4282 0.006
R23997 vp_p.n4272 vp_p.n4271 0.006
R23998 vp_p.n4269 vp_p.n4268 0.006
R23999 vp_p.n4258 vp_p.n4257 0.006
R24000 vp_p.n4255 vp_p.n4254 0.006
R24001 vp_p.n4244 vp_p.n4243 0.006
R24002 vp_p.n4241 vp_p.n4240 0.006
R24003 vp_p.n4230 vp_p.n4229 0.006
R24004 vp_p.n4227 vp_p.n4226 0.006
R24005 vp_p.n4216 vp_p.n4215 0.006
R24006 vp_p.n4213 vp_p.n4212 0.006
R24007 vp_p.n4202 vp_p.n4201 0.006
R24008 vp_p.n4199 vp_p.n4198 0.006
R24009 vp_p.n4188 vp_p.n4187 0.006
R24010 vp_p.n4185 vp_p.n4184 0.006
R24011 vp_p.n4174 vp_p.n4173 0.006
R24012 vp_p.n4171 vp_p.n4170 0.006
R24013 vp_p.n4160 vp_p.n4159 0.006
R24014 vp_p.n4157 vp_p.n4156 0.006
R24015 vp_p.n4146 vp_p.n4145 0.006
R24016 vp_p.n4143 vp_p.n4142 0.006
R24017 vp_p.n4132 vp_p.n4131 0.006
R24018 vp_p.n4129 vp_p.n4128 0.006
R24019 vp_p.n4118 vp_p.n4117 0.006
R24020 vp_p.n4115 vp_p.n4114 0.006
R24021 vp_p.n4104 vp_p.n4103 0.006
R24022 vp_p.n4101 vp_p.n4100 0.006
R24023 vp_p.n4090 vp_p.n4089 0.006
R24024 vp_p.n4087 vp_p.n4086 0.006
R24025 vp_p.n4076 vp_p.n4075 0.006
R24026 vp_p.n4073 vp_p.n4072 0.006
R24027 vp_p.n4062 vp_p.n4061 0.006
R24028 vp_p.n4059 vp_p.n4058 0.006
R24029 vp_p.n4048 vp_p.n4047 0.006
R24030 vp_p.n4045 vp_p.n4044 0.006
R24031 vp_p.n4034 vp_p.n4033 0.006
R24032 vp_p.n4031 vp_p.n4030 0.006
R24033 vp_p.n4020 vp_p.n4019 0.006
R24034 vp_p.n4017 vp_p.n4016 0.006
R24035 vp_p.n4006 vp_p.n4005 0.006
R24036 vp_p.n4003 vp_p.n4002 0.006
R24037 vp_p.n3992 vp_p.n3991 0.006
R24038 vp_p.n3989 vp_p.n3988 0.006
R24039 vp_p.n3978 vp_p.n3977 0.006
R24040 vp_p.n3975 vp_p.n3974 0.006
R24041 vp_p.n3964 vp_p.n3963 0.006
R24042 vp_p.n3961 vp_p.n3960 0.006
R24043 vp_p.n3950 vp_p.n3949 0.006
R24044 vp_p.n3947 vp_p.n3946 0.006
R24045 vp_p.n3936 vp_p.n3935 0.006
R24046 vp_p.n3933 vp_p.n3932 0.006
R24047 vp_p.n3922 vp_p.n3921 0.006
R24048 vp_p.n3919 vp_p.n3918 0.006
R24049 vp_p.n3908 vp_p.n3907 0.006
R24050 vp_p.n3905 vp_p.n3904 0.006
R24051 vp_p.n3894 vp_p.n3893 0.006
R24052 vp_p.n3891 vp_p.n3890 0.006
R24053 vp_p.n3880 vp_p.n3879 0.006
R24054 vp_p.n3877 vp_p.n3876 0.006
R24055 vp_p.n3866 vp_p.n3865 0.006
R24056 vp_p.n3863 vp_p.n3862 0.006
R24057 vp_p.n3852 vp_p.n3851 0.006
R24058 vp_p.n3849 vp_p.n3848 0.006
R24059 vp_p.n3838 vp_p.n3837 0.006
R24060 vp_p.n3835 vp_p.n3834 0.006
R24061 vp_p.n3824 vp_p.n3823 0.006
R24062 vp_p.n3821 vp_p.n3820 0.006
R24063 vp_p.n3810 vp_p.n3809 0.006
R24064 vp_p.n3807 vp_p.n3806 0.006
R24065 vp_p.n3796 vp_p.n3795 0.006
R24066 vp_p.n3793 vp_p.n3792 0.006
R24067 vp_p.n3782 vp_p.n3781 0.006
R24068 vp_p.n3779 vp_p.n3778 0.006
R24069 vp_p.n3768 vp_p.n3767 0.006
R24070 vp_p.n3765 vp_p.n3764 0.006
R24071 vp_p.n3754 vp_p.n3753 0.006
R24072 vp_p.n3751 vp_p.n3750 0.006
R24073 vp_p.n3740 vp_p.n3739 0.006
R24074 vp_p.n3737 vp_p.n3736 0.006
R24075 vp_p.n3726 vp_p.n3725 0.006
R24076 vp_p.n3723 vp_p.n3722 0.006
R24077 vp_p.n3712 vp_p.n3711 0.006
R24078 vp_p.n3709 vp_p.n3708 0.006
R24079 vp_p.n3698 vp_p.n3697 0.006
R24080 vp_p.n3695 vp_p.n3694 0.006
R24081 vp_p.n3684 vp_p.n3683 0.006
R24082 vp_p.n3681 vp_p.n3680 0.006
R24083 vp_p.n3670 vp_p.n3669 0.006
R24084 vp_p.n3667 vp_p.n3666 0.006
R24085 vp_p.n3656 vp_p.n3655 0.006
R24086 vp_p.n3653 vp_p.n3652 0.006
R24087 vp_p.n3642 vp_p.n3641 0.006
R24088 vp_p.n3639 vp_p.n3638 0.006
R24089 vp_p.n3628 vp_p.n3627 0.006
R24090 vp_p.n3625 vp_p.n3624 0.006
R24091 vp_p.n3614 vp_p.n3613 0.006
R24092 vp_p.n3611 vp_p.n3610 0.006
R24093 vp_p.n3600 vp_p.n3599 0.006
R24094 vp_p.n3597 vp_p.n3596 0.006
R24095 vp_p.n3586 vp_p.n3585 0.006
R24096 vp_p.n3583 vp_p.n3582 0.006
R24097 vp_p.n3572 vp_p.n3571 0.006
R24098 vp_p.n3569 vp_p.n3568 0.006
R24099 vp_p.n3558 vp_p.n3557 0.006
R24100 vp_p.n3555 vp_p.n3554 0.006
R24101 vp_p.n3544 vp_p.n3543 0.006
R24102 vp_p.n3541 vp_p.n3540 0.006
R24103 vp_p.n3530 vp_p.n3529 0.006
R24104 vp_p.n3527 vp_p.n3526 0.006
R24105 vp_p.n3516 vp_p.n3515 0.006
R24106 vp_p.n3513 vp_p.n3512 0.006
R24107 vp_p.n3502 vp_p.n3501 0.006
R24108 vp_p.n3499 vp_p.n3498 0.006
R24109 vp_p.n3488 vp_p.n3487 0.006
R24110 vp_p.n3485 vp_p.n3484 0.006
R24111 vp_p.n3474 vp_p.n3473 0.006
R24112 vp_p.n3471 vp_p.n3470 0.006
R24113 vp_p.n3460 vp_p.n3459 0.006
R24114 vp_p.n3457 vp_p.n3456 0.006
R24115 vp_p.n3446 vp_p.n3445 0.006
R24116 vp_p.n3443 vp_p.n3442 0.006
R24117 vp_p.n3432 vp_p.n3431 0.006
R24118 vp_p.n3429 vp_p.n3428 0.006
R24119 vp_p.n3418 vp_p.n3417 0.006
R24120 vp_p.n3415 vp_p.n3414 0.006
R24121 vp_p.n3404 vp_p.n3403 0.006
R24122 vp_p.n3401 vp_p.n3400 0.006
R24123 vp_p.n3390 vp_p.n3389 0.006
R24124 vp_p.n3387 vp_p.n3386 0.006
R24125 vp_p.n3376 vp_p.n3375 0.006
R24126 vp_p.n3373 vp_p.n3372 0.006
R24127 vp_p.n3362 vp_p.n3361 0.006
R24128 vp_p.n3359 vp_p.n3358 0.006
R24129 vp_p.n3348 vp_p.n3347 0.006
R24130 vp_p.n3345 vp_p.n3344 0.006
R24131 vp_p.n3334 vp_p.n3333 0.006
R24132 vp_p.n3331 vp_p.n3330 0.006
R24133 vp_p.n3320 vp_p.n3319 0.006
R24134 vp_p.n4314 vp_p.n4313 0.006
R24135 vp_p.n2891 vp_p.n2890 0.006
R24136 vp_p.n1461 vp_p.n1460 0.006
R24137 vp_p.n10203 vp_p.n10202 0.006
R24138 vp_p.n11636 vp_p.n11635 0.006
R24139 vp_p.n13070 vp_p.n13069 0.006
R24140 vp_p.n14439 vp_p.n14438 0.006
R24141 vp_p.n15872 vp_p.n15871 0.006
R24142 vp_p.n17304 vp_p.n17303 0.006
R24143 vp_p.n18735 vp_p.n18734 0.006
R24144 vp_p.n20165 vp_p.n20164 0.006
R24145 vp_p.n21594 vp_p.n21593 0.006
R24146 vp_p.n22013 vp_p.n22012 0.006
R24147 vp_p.n22018 vp_p.n22017 0.006
R24148 vp_p.n22029 vp_p.n22023 0.006
R24149 vp_p.n22033 vp_p.n22032 0.006
R24150 vp_p.n22043 vp_p.n22037 0.006
R24151 vp_p.n22047 vp_p.n22046 0.006
R24152 vp_p.n22057 vp_p.n22051 0.006
R24153 vp_p.n22061 vp_p.n22060 0.006
R24154 vp_p.n22071 vp_p.n22065 0.006
R24155 vp_p.n22075 vp_p.n22074 0.006
R24156 vp_p.n22085 vp_p.n22079 0.006
R24157 vp_p.n22089 vp_p.n22088 0.006
R24158 vp_p.n22099 vp_p.n22093 0.006
R24159 vp_p.n22103 vp_p.n22102 0.006
R24160 vp_p.n22113 vp_p.n22107 0.006
R24161 vp_p.n22117 vp_p.n22116 0.006
R24162 vp_p.n22127 vp_p.n22121 0.006
R24163 vp_p.n22131 vp_p.n22130 0.006
R24164 vp_p.n22141 vp_p.n22135 0.006
R24165 vp_p.n22145 vp_p.n22144 0.006
R24166 vp_p.n22155 vp_p.n22149 0.006
R24167 vp_p.n22159 vp_p.n22158 0.006
R24168 vp_p.n22169 vp_p.n22163 0.006
R24169 vp_p.n22173 vp_p.n22172 0.006
R24170 vp_p.n22183 vp_p.n22177 0.006
R24171 vp_p.n22187 vp_p.n22186 0.006
R24172 vp_p.n22197 vp_p.n22191 0.006
R24173 vp_p.n22201 vp_p.n22200 0.006
R24174 vp_p.n22211 vp_p.n22205 0.006
R24175 vp_p.n22215 vp_p.n22214 0.006
R24176 vp_p.n22225 vp_p.n22219 0.006
R24177 vp_p.n22229 vp_p.n22228 0.006
R24178 vp_p.n22239 vp_p.n22233 0.006
R24179 vp_p.n22243 vp_p.n22242 0.006
R24180 vp_p.n22253 vp_p.n22247 0.006
R24181 vp_p.n22257 vp_p.n22256 0.006
R24182 vp_p.n22267 vp_p.n22261 0.006
R24183 vp_p.n22271 vp_p.n22270 0.006
R24184 vp_p.n22281 vp_p.n22275 0.006
R24185 vp_p.n22285 vp_p.n22284 0.006
R24186 vp_p.n22295 vp_p.n22289 0.006
R24187 vp_p.n22299 vp_p.n22298 0.006
R24188 vp_p.n22309 vp_p.n22303 0.006
R24189 vp_p.n22313 vp_p.n22312 0.006
R24190 vp_p.n22323 vp_p.n22317 0.006
R24191 vp_p.n22327 vp_p.n22326 0.006
R24192 vp_p.n22337 vp_p.n22331 0.006
R24193 vp_p.n22341 vp_p.n22340 0.006
R24194 vp_p.n22351 vp_p.n22345 0.006
R24195 vp_p.n22355 vp_p.n22354 0.006
R24196 vp_p.n22365 vp_p.n22359 0.006
R24197 vp_p.n22369 vp_p.n22368 0.006
R24198 vp_p.n22379 vp_p.n22373 0.006
R24199 vp_p.n22383 vp_p.n22382 0.006
R24200 vp_p.n22393 vp_p.n22387 0.006
R24201 vp_p.n22397 vp_p.n22396 0.006
R24202 vp_p.n22407 vp_p.n22401 0.006
R24203 vp_p.n22411 vp_p.n22410 0.006
R24204 vp_p.n22421 vp_p.n22415 0.006
R24205 vp_p.n22425 vp_p.n22424 0.006
R24206 vp_p.n22435 vp_p.n22429 0.006
R24207 vp_p.n22439 vp_p.n22438 0.006
R24208 vp_p.n22449 vp_p.n22443 0.006
R24209 vp_p.n22453 vp_p.n22452 0.006
R24210 vp_p.n22463 vp_p.n22457 0.006
R24211 vp_p.n22467 vp_p.n22466 0.006
R24212 vp_p.n22477 vp_p.n22471 0.006
R24213 vp_p.n22481 vp_p.n22480 0.006
R24214 vp_p.n22491 vp_p.n22485 0.006
R24215 vp_p.n22495 vp_p.n22494 0.006
R24216 vp_p.n22505 vp_p.n22499 0.006
R24217 vp_p.n22509 vp_p.n22508 0.006
R24218 vp_p.n22519 vp_p.n22513 0.006
R24219 vp_p.n22523 vp_p.n22522 0.006
R24220 vp_p.n22533 vp_p.n22527 0.006
R24221 vp_p.n22537 vp_p.n22536 0.006
R24222 vp_p.n22547 vp_p.n22541 0.006
R24223 vp_p.n22551 vp_p.n22550 0.006
R24224 vp_p.n22561 vp_p.n22555 0.006
R24225 vp_p.n22565 vp_p.n22564 0.006
R24226 vp_p.n22575 vp_p.n22569 0.006
R24227 vp_p.n22579 vp_p.n22578 0.006
R24228 vp_p.n22589 vp_p.n22583 0.006
R24229 vp_p.n22593 vp_p.n22592 0.006
R24230 vp_p.n22603 vp_p.n22597 0.006
R24231 vp_p.n22607 vp_p.n22606 0.006
R24232 vp_p.n22617 vp_p.n22611 0.006
R24233 vp_p.n22621 vp_p.n22620 0.006
R24234 vp_p.n22631 vp_p.n22625 0.006
R24235 vp_p.n22635 vp_p.n22634 0.006
R24236 vp_p.n22645 vp_p.n22639 0.006
R24237 vp_p.n22649 vp_p.n22648 0.006
R24238 vp_p.n22659 vp_p.n22653 0.006
R24239 vp_p.n22663 vp_p.n22662 0.006
R24240 vp_p.n22673 vp_p.n22667 0.006
R24241 vp_p.n22677 vp_p.n22676 0.006
R24242 vp_p.n22687 vp_p.n22681 0.006
R24243 vp_p.n22691 vp_p.n22690 0.006
R24244 vp_p.n22701 vp_p.n22695 0.006
R24245 vp_p.n22705 vp_p.n22704 0.006
R24246 vp_p.n22715 vp_p.n22709 0.006
R24247 vp_p.n22719 vp_p.n22718 0.006
R24248 vp_p.n22729 vp_p.n22723 0.006
R24249 vp_p.n22733 vp_p.n22732 0.006
R24250 vp_p.n22743 vp_p.n22737 0.006
R24251 vp_p.n22747 vp_p.n22746 0.006
R24252 vp_p.n22757 vp_p.n22751 0.006
R24253 vp_p.n22761 vp_p.n22760 0.006
R24254 vp_p.n22771 vp_p.n22765 0.006
R24255 vp_p.n22775 vp_p.n22774 0.006
R24256 vp_p.n22785 vp_p.n22779 0.006
R24257 vp_p.n22789 vp_p.n22788 0.006
R24258 vp_p.n22799 vp_p.n22793 0.006
R24259 vp_p.n22803 vp_p.n22802 0.006
R24260 vp_p.n22813 vp_p.n22807 0.006
R24261 vp_p.n22817 vp_p.n22816 0.006
R24262 vp_p.n22827 vp_p.n22821 0.006
R24263 vp_p.n22831 vp_p.n22830 0.006
R24264 vp_p.n22841 vp_p.n22835 0.006
R24265 vp_p.n22845 vp_p.n22844 0.006
R24266 vp_p.n22855 vp_p.n22849 0.006
R24267 vp_p.n22859 vp_p.n22858 0.006
R24268 vp_p.n22869 vp_p.n22863 0.006
R24269 vp_p.n22873 vp_p.n22872 0.006
R24270 vp_p.n22883 vp_p.n22877 0.006
R24271 vp_p.n22887 vp_p.n22886 0.006
R24272 vp_p.n22897 vp_p.n22891 0.006
R24273 vp_p.n22901 vp_p.n22900 0.006
R24274 vp_p.n22911 vp_p.n22905 0.006
R24275 vp_p.n22915 vp_p.n22914 0.006
R24276 vp_p.n22925 vp_p.n22919 0.006
R24277 vp_p.n22929 vp_p.n22928 0.006
R24278 vp_p.n22939 vp_p.n22933 0.006
R24279 vp_p.n22943 vp_p.n22942 0.006
R24280 vp_p.n22953 vp_p.n22947 0.006
R24281 vp_p.n22957 vp_p.n22956 0.006
R24282 vp_p.n22967 vp_p.n22961 0.006
R24283 vp_p.n22971 vp_p.n22970 0.006
R24284 vp_p.n22981 vp_p.n22975 0.006
R24285 vp_p.n22985 vp_p.n22984 0.006
R24286 vp_p.n22995 vp_p.n22989 0.006
R24287 vp_p.n22999 vp_p.n22998 0.006
R24288 vp_p.n23009 vp_p.n23003 0.006
R24289 vp_p.n23013 vp_p.n23012 0.006
R24290 vp_p.n23017 vp_p.n23016 0.006
R24291 vp_p.n23027 vp_p.n23021 0.006
R24292 vp_p.n23031 vp_p.n23030 0.006
R24293 vp_p.n23036 vp_p.n23035 0.006
R24294 vp_p.n23041 vp_p.n23040 0.006
R24295 vp_p.n23046 vp_p.n23045 0.006
R24296 vp_p.n23018 vp_p.n23017 0.006
R24297 vp_p.n23014 vp_p.n23013 0.006
R24298 vp_p.n23003 vp_p.n23002 0.006
R24299 vp_p.n23000 vp_p.n22999 0.006
R24300 vp_p.n22989 vp_p.n22988 0.006
R24301 vp_p.n22986 vp_p.n22985 0.006
R24302 vp_p.n22975 vp_p.n22974 0.006
R24303 vp_p.n22972 vp_p.n22971 0.006
R24304 vp_p.n22961 vp_p.n22960 0.006
R24305 vp_p.n22958 vp_p.n22957 0.006
R24306 vp_p.n22947 vp_p.n22946 0.006
R24307 vp_p.n22944 vp_p.n22943 0.006
R24308 vp_p.n22933 vp_p.n22932 0.006
R24309 vp_p.n22930 vp_p.n22929 0.006
R24310 vp_p.n22919 vp_p.n22918 0.006
R24311 vp_p.n22916 vp_p.n22915 0.006
R24312 vp_p.n22905 vp_p.n22904 0.006
R24313 vp_p.n22902 vp_p.n22901 0.006
R24314 vp_p.n22891 vp_p.n22890 0.006
R24315 vp_p.n22888 vp_p.n22887 0.006
R24316 vp_p.n22877 vp_p.n22876 0.006
R24317 vp_p.n22874 vp_p.n22873 0.006
R24318 vp_p.n22863 vp_p.n22862 0.006
R24319 vp_p.n22860 vp_p.n22859 0.006
R24320 vp_p.n22849 vp_p.n22848 0.006
R24321 vp_p.n22846 vp_p.n22845 0.006
R24322 vp_p.n22835 vp_p.n22834 0.006
R24323 vp_p.n22832 vp_p.n22831 0.006
R24324 vp_p.n22821 vp_p.n22820 0.006
R24325 vp_p.n22818 vp_p.n22817 0.006
R24326 vp_p.n22807 vp_p.n22806 0.006
R24327 vp_p.n22804 vp_p.n22803 0.006
R24328 vp_p.n22793 vp_p.n22792 0.006
R24329 vp_p.n22790 vp_p.n22789 0.006
R24330 vp_p.n22779 vp_p.n22778 0.006
R24331 vp_p.n22776 vp_p.n22775 0.006
R24332 vp_p.n22765 vp_p.n22764 0.006
R24333 vp_p.n22762 vp_p.n22761 0.006
R24334 vp_p.n22751 vp_p.n22750 0.006
R24335 vp_p.n22748 vp_p.n22747 0.006
R24336 vp_p.n22737 vp_p.n22736 0.006
R24337 vp_p.n22734 vp_p.n22733 0.006
R24338 vp_p.n22723 vp_p.n22722 0.006
R24339 vp_p.n22720 vp_p.n22719 0.006
R24340 vp_p.n22709 vp_p.n22708 0.006
R24341 vp_p.n22706 vp_p.n22705 0.006
R24342 vp_p.n22695 vp_p.n22694 0.006
R24343 vp_p.n22692 vp_p.n22691 0.006
R24344 vp_p.n22681 vp_p.n22680 0.006
R24345 vp_p.n22678 vp_p.n22677 0.006
R24346 vp_p.n22667 vp_p.n22666 0.006
R24347 vp_p.n22664 vp_p.n22663 0.006
R24348 vp_p.n22653 vp_p.n22652 0.006
R24349 vp_p.n22650 vp_p.n22649 0.006
R24350 vp_p.n22639 vp_p.n22638 0.006
R24351 vp_p.n22636 vp_p.n22635 0.006
R24352 vp_p.n22625 vp_p.n22624 0.006
R24353 vp_p.n22622 vp_p.n22621 0.006
R24354 vp_p.n22611 vp_p.n22610 0.006
R24355 vp_p.n22608 vp_p.n22607 0.006
R24356 vp_p.n22597 vp_p.n22596 0.006
R24357 vp_p.n22594 vp_p.n22593 0.006
R24358 vp_p.n22583 vp_p.n22582 0.006
R24359 vp_p.n22580 vp_p.n22579 0.006
R24360 vp_p.n22569 vp_p.n22568 0.006
R24361 vp_p.n22566 vp_p.n22565 0.006
R24362 vp_p.n22555 vp_p.n22554 0.006
R24363 vp_p.n22552 vp_p.n22551 0.006
R24364 vp_p.n22541 vp_p.n22540 0.006
R24365 vp_p.n22538 vp_p.n22537 0.006
R24366 vp_p.n22527 vp_p.n22526 0.006
R24367 vp_p.n22524 vp_p.n22523 0.006
R24368 vp_p.n22513 vp_p.n22512 0.006
R24369 vp_p.n22510 vp_p.n22509 0.006
R24370 vp_p.n22499 vp_p.n22498 0.006
R24371 vp_p.n22496 vp_p.n22495 0.006
R24372 vp_p.n22485 vp_p.n22484 0.006
R24373 vp_p.n22482 vp_p.n22481 0.006
R24374 vp_p.n22471 vp_p.n22470 0.006
R24375 vp_p.n22468 vp_p.n22467 0.006
R24376 vp_p.n22457 vp_p.n22456 0.006
R24377 vp_p.n22454 vp_p.n22453 0.006
R24378 vp_p.n22443 vp_p.n22442 0.006
R24379 vp_p.n22440 vp_p.n22439 0.006
R24380 vp_p.n22429 vp_p.n22428 0.006
R24381 vp_p.n22426 vp_p.n22425 0.006
R24382 vp_p.n22415 vp_p.n22414 0.006
R24383 vp_p.n22412 vp_p.n22411 0.006
R24384 vp_p.n22401 vp_p.n22400 0.006
R24385 vp_p.n22398 vp_p.n22397 0.006
R24386 vp_p.n22387 vp_p.n22386 0.006
R24387 vp_p.n22384 vp_p.n22383 0.006
R24388 vp_p.n22373 vp_p.n22372 0.006
R24389 vp_p.n22370 vp_p.n22369 0.006
R24390 vp_p.n22359 vp_p.n22358 0.006
R24391 vp_p.n22356 vp_p.n22355 0.006
R24392 vp_p.n22345 vp_p.n22344 0.006
R24393 vp_p.n22342 vp_p.n22341 0.006
R24394 vp_p.n22331 vp_p.n22330 0.006
R24395 vp_p.n22328 vp_p.n22327 0.006
R24396 vp_p.n22317 vp_p.n22316 0.006
R24397 vp_p.n22314 vp_p.n22313 0.006
R24398 vp_p.n22303 vp_p.n22302 0.006
R24399 vp_p.n22300 vp_p.n22299 0.006
R24400 vp_p.n22289 vp_p.n22288 0.006
R24401 vp_p.n22286 vp_p.n22285 0.006
R24402 vp_p.n22275 vp_p.n22274 0.006
R24403 vp_p.n22272 vp_p.n22271 0.006
R24404 vp_p.n22261 vp_p.n22260 0.006
R24405 vp_p.n22258 vp_p.n22257 0.006
R24406 vp_p.n22247 vp_p.n22246 0.006
R24407 vp_p.n22244 vp_p.n22243 0.006
R24408 vp_p.n22233 vp_p.n22232 0.006
R24409 vp_p.n22230 vp_p.n22229 0.006
R24410 vp_p.n22219 vp_p.n22218 0.006
R24411 vp_p.n22216 vp_p.n22215 0.006
R24412 vp_p.n22205 vp_p.n22204 0.006
R24413 vp_p.n22202 vp_p.n22201 0.006
R24414 vp_p.n22191 vp_p.n22190 0.006
R24415 vp_p.n22188 vp_p.n22187 0.006
R24416 vp_p.n22177 vp_p.n22176 0.006
R24417 vp_p.n22174 vp_p.n22173 0.006
R24418 vp_p.n22163 vp_p.n22162 0.006
R24419 vp_p.n22160 vp_p.n22159 0.006
R24420 vp_p.n22149 vp_p.n22148 0.006
R24421 vp_p.n22146 vp_p.n22145 0.006
R24422 vp_p.n22135 vp_p.n22134 0.006
R24423 vp_p.n22132 vp_p.n22131 0.006
R24424 vp_p.n22121 vp_p.n22120 0.006
R24425 vp_p.n22118 vp_p.n22117 0.006
R24426 vp_p.n22107 vp_p.n22106 0.006
R24427 vp_p.n22104 vp_p.n22103 0.006
R24428 vp_p.n22093 vp_p.n22092 0.006
R24429 vp_p.n22090 vp_p.n22089 0.006
R24430 vp_p.n22079 vp_p.n22078 0.006
R24431 vp_p.n22076 vp_p.n22075 0.006
R24432 vp_p.n22065 vp_p.n22064 0.006
R24433 vp_p.n22062 vp_p.n22061 0.006
R24434 vp_p.n22051 vp_p.n22050 0.006
R24435 vp_p.n22048 vp_p.n22047 0.006
R24436 vp_p.n22037 vp_p.n22036 0.006
R24437 vp_p.n22034 vp_p.n22033 0.006
R24438 vp_p.n22023 vp_p.n22022 0.006
R24439 vp_p.n23021 vp_p.n23020 0.006
R24440 vp_p.n21599 vp_p.n21598 0.006
R24441 vp_p.n20170 vp_p.n20169 0.006
R24442 vp_p.n18740 vp_p.n18739 0.006
R24443 vp_p.n17309 vp_p.n17308 0.006
R24444 vp_p.n15877 vp_p.n15876 0.006
R24445 vp_p.n14444 vp_p.n14443 0.006
R24446 vp_p.n13075 vp_p.n13074 0.006
R24447 vp_p.n11641 vp_p.n11640 0.006
R24448 vp_p.n10208 vp_p.n10207 0.006
R24449 vp_p.n1466 vp_p.n1465 0.006
R24450 vp_p.n2896 vp_p.n2895 0.006
R24451 vp_p.n4325 vp_p.n4324 0.006
R24452 vp_p.n4734 vp_p.n4733 0.006
R24453 vp_p.n4739 vp_p.n4738 0.006
R24454 vp_p.n4750 vp_p.n4744 0.006
R24455 vp_p.n4754 vp_p.n4753 0.006
R24456 vp_p.n4764 vp_p.n4758 0.006
R24457 vp_p.n4768 vp_p.n4767 0.006
R24458 vp_p.n4778 vp_p.n4772 0.006
R24459 vp_p.n4782 vp_p.n4781 0.006
R24460 vp_p.n4792 vp_p.n4786 0.006
R24461 vp_p.n4796 vp_p.n4795 0.006
R24462 vp_p.n4806 vp_p.n4800 0.006
R24463 vp_p.n4810 vp_p.n4809 0.006
R24464 vp_p.n4820 vp_p.n4814 0.006
R24465 vp_p.n4824 vp_p.n4823 0.006
R24466 vp_p.n4834 vp_p.n4828 0.006
R24467 vp_p.n4838 vp_p.n4837 0.006
R24468 vp_p.n4848 vp_p.n4842 0.006
R24469 vp_p.n4852 vp_p.n4851 0.006
R24470 vp_p.n4862 vp_p.n4856 0.006
R24471 vp_p.n4866 vp_p.n4865 0.006
R24472 vp_p.n4876 vp_p.n4870 0.006
R24473 vp_p.n4880 vp_p.n4879 0.006
R24474 vp_p.n4890 vp_p.n4884 0.006
R24475 vp_p.n4894 vp_p.n4893 0.006
R24476 vp_p.n4904 vp_p.n4898 0.006
R24477 vp_p.n4908 vp_p.n4907 0.006
R24478 vp_p.n4918 vp_p.n4912 0.006
R24479 vp_p.n4922 vp_p.n4921 0.006
R24480 vp_p.n4932 vp_p.n4926 0.006
R24481 vp_p.n4936 vp_p.n4935 0.006
R24482 vp_p.n4946 vp_p.n4940 0.006
R24483 vp_p.n4950 vp_p.n4949 0.006
R24484 vp_p.n4960 vp_p.n4954 0.006
R24485 vp_p.n4964 vp_p.n4963 0.006
R24486 vp_p.n4974 vp_p.n4968 0.006
R24487 vp_p.n4978 vp_p.n4977 0.006
R24488 vp_p.n4988 vp_p.n4982 0.006
R24489 vp_p.n4992 vp_p.n4991 0.006
R24490 vp_p.n5002 vp_p.n4996 0.006
R24491 vp_p.n5006 vp_p.n5005 0.006
R24492 vp_p.n5016 vp_p.n5010 0.006
R24493 vp_p.n5020 vp_p.n5019 0.006
R24494 vp_p.n5030 vp_p.n5024 0.006
R24495 vp_p.n5034 vp_p.n5033 0.006
R24496 vp_p.n5044 vp_p.n5038 0.006
R24497 vp_p.n5048 vp_p.n5047 0.006
R24498 vp_p.n5058 vp_p.n5052 0.006
R24499 vp_p.n5062 vp_p.n5061 0.006
R24500 vp_p.n5072 vp_p.n5066 0.006
R24501 vp_p.n5076 vp_p.n5075 0.006
R24502 vp_p.n5086 vp_p.n5080 0.006
R24503 vp_p.n5090 vp_p.n5089 0.006
R24504 vp_p.n5100 vp_p.n5094 0.006
R24505 vp_p.n5104 vp_p.n5103 0.006
R24506 vp_p.n5114 vp_p.n5108 0.006
R24507 vp_p.n5118 vp_p.n5117 0.006
R24508 vp_p.n5128 vp_p.n5122 0.006
R24509 vp_p.n5132 vp_p.n5131 0.006
R24510 vp_p.n5142 vp_p.n5136 0.006
R24511 vp_p.n5146 vp_p.n5145 0.006
R24512 vp_p.n5156 vp_p.n5150 0.006
R24513 vp_p.n5160 vp_p.n5159 0.006
R24514 vp_p.n5170 vp_p.n5164 0.006
R24515 vp_p.n5174 vp_p.n5173 0.006
R24516 vp_p.n5184 vp_p.n5178 0.006
R24517 vp_p.n5188 vp_p.n5187 0.006
R24518 vp_p.n5198 vp_p.n5192 0.006
R24519 vp_p.n5202 vp_p.n5201 0.006
R24520 vp_p.n5212 vp_p.n5206 0.006
R24521 vp_p.n5216 vp_p.n5215 0.006
R24522 vp_p.n5226 vp_p.n5220 0.006
R24523 vp_p.n5230 vp_p.n5229 0.006
R24524 vp_p.n5240 vp_p.n5234 0.006
R24525 vp_p.n5244 vp_p.n5243 0.006
R24526 vp_p.n5254 vp_p.n5248 0.006
R24527 vp_p.n5258 vp_p.n5257 0.006
R24528 vp_p.n5268 vp_p.n5262 0.006
R24529 vp_p.n5272 vp_p.n5271 0.006
R24530 vp_p.n5282 vp_p.n5276 0.006
R24531 vp_p.n5286 vp_p.n5285 0.006
R24532 vp_p.n5296 vp_p.n5290 0.006
R24533 vp_p.n5300 vp_p.n5299 0.006
R24534 vp_p.n5310 vp_p.n5304 0.006
R24535 vp_p.n5314 vp_p.n5313 0.006
R24536 vp_p.n5324 vp_p.n5318 0.006
R24537 vp_p.n5328 vp_p.n5327 0.006
R24538 vp_p.n5338 vp_p.n5332 0.006
R24539 vp_p.n5342 vp_p.n5341 0.006
R24540 vp_p.n5352 vp_p.n5346 0.006
R24541 vp_p.n5356 vp_p.n5355 0.006
R24542 vp_p.n5366 vp_p.n5360 0.006
R24543 vp_p.n5370 vp_p.n5369 0.006
R24544 vp_p.n5380 vp_p.n5374 0.006
R24545 vp_p.n5384 vp_p.n5383 0.006
R24546 vp_p.n5394 vp_p.n5388 0.006
R24547 vp_p.n5398 vp_p.n5397 0.006
R24548 vp_p.n5408 vp_p.n5402 0.006
R24549 vp_p.n5412 vp_p.n5411 0.006
R24550 vp_p.n5422 vp_p.n5416 0.006
R24551 vp_p.n5426 vp_p.n5425 0.006
R24552 vp_p.n5436 vp_p.n5430 0.006
R24553 vp_p.n5440 vp_p.n5439 0.006
R24554 vp_p.n5450 vp_p.n5444 0.006
R24555 vp_p.n5454 vp_p.n5453 0.006
R24556 vp_p.n5464 vp_p.n5458 0.006
R24557 vp_p.n5468 vp_p.n5467 0.006
R24558 vp_p.n5478 vp_p.n5472 0.006
R24559 vp_p.n5482 vp_p.n5481 0.006
R24560 vp_p.n5492 vp_p.n5486 0.006
R24561 vp_p.n5496 vp_p.n5495 0.006
R24562 vp_p.n5506 vp_p.n5500 0.006
R24563 vp_p.n5510 vp_p.n5509 0.006
R24564 vp_p.n5520 vp_p.n5514 0.006
R24565 vp_p.n5524 vp_p.n5523 0.006
R24566 vp_p.n5534 vp_p.n5528 0.006
R24567 vp_p.n5538 vp_p.n5537 0.006
R24568 vp_p.n5548 vp_p.n5542 0.006
R24569 vp_p.n5552 vp_p.n5551 0.006
R24570 vp_p.n5562 vp_p.n5556 0.006
R24571 vp_p.n5566 vp_p.n5565 0.006
R24572 vp_p.n5576 vp_p.n5570 0.006
R24573 vp_p.n5580 vp_p.n5579 0.006
R24574 vp_p.n5590 vp_p.n5584 0.006
R24575 vp_p.n5594 vp_p.n5593 0.006
R24576 vp_p.n5604 vp_p.n5598 0.006
R24577 vp_p.n5608 vp_p.n5607 0.006
R24578 vp_p.n5618 vp_p.n5612 0.006
R24579 vp_p.n5622 vp_p.n5621 0.006
R24580 vp_p.n5632 vp_p.n5626 0.006
R24581 vp_p.n5636 vp_p.n5635 0.006
R24582 vp_p.n5646 vp_p.n5640 0.006
R24583 vp_p.n5650 vp_p.n5649 0.006
R24584 vp_p.n5660 vp_p.n5654 0.006
R24585 vp_p.n5664 vp_p.n5663 0.006
R24586 vp_p.n5674 vp_p.n5668 0.006
R24587 vp_p.n5678 vp_p.n5677 0.006
R24588 vp_p.n5688 vp_p.n5682 0.006
R24589 vp_p.n5692 vp_p.n5691 0.006
R24590 vp_p.n5702 vp_p.n5696 0.006
R24591 vp_p.n5706 vp_p.n5705 0.006
R24592 vp_p.n5716 vp_p.n5710 0.006
R24593 vp_p.n5720 vp_p.n5719 0.006
R24594 vp_p.n5730 vp_p.n5724 0.006
R24595 vp_p.n5734 vp_p.n5733 0.006
R24596 vp_p.n5744 vp_p.n5738 0.006
R24597 vp_p.n5748 vp_p.n5747 0.006
R24598 vp_p.n5758 vp_p.n5752 0.006
R24599 vp_p.n5762 vp_p.n5761 0.006
R24600 vp_p.n5767 vp_p.n5766 0.006
R24601 vp_p.n5772 vp_p.n5771 0.006
R24602 vp_p.n5749 vp_p.n5748 0.006
R24603 vp_p.n5738 vp_p.n5737 0.006
R24604 vp_p.n5735 vp_p.n5734 0.006
R24605 vp_p.n5724 vp_p.n5723 0.006
R24606 vp_p.n5721 vp_p.n5720 0.006
R24607 vp_p.n5710 vp_p.n5709 0.006
R24608 vp_p.n5707 vp_p.n5706 0.006
R24609 vp_p.n5696 vp_p.n5695 0.006
R24610 vp_p.n5693 vp_p.n5692 0.006
R24611 vp_p.n5682 vp_p.n5681 0.006
R24612 vp_p.n5679 vp_p.n5678 0.006
R24613 vp_p.n5668 vp_p.n5667 0.006
R24614 vp_p.n5665 vp_p.n5664 0.006
R24615 vp_p.n5654 vp_p.n5653 0.006
R24616 vp_p.n5651 vp_p.n5650 0.006
R24617 vp_p.n5640 vp_p.n5639 0.006
R24618 vp_p.n5637 vp_p.n5636 0.006
R24619 vp_p.n5626 vp_p.n5625 0.006
R24620 vp_p.n5623 vp_p.n5622 0.006
R24621 vp_p.n5612 vp_p.n5611 0.006
R24622 vp_p.n5609 vp_p.n5608 0.006
R24623 vp_p.n5598 vp_p.n5597 0.006
R24624 vp_p.n5595 vp_p.n5594 0.006
R24625 vp_p.n5584 vp_p.n5583 0.006
R24626 vp_p.n5581 vp_p.n5580 0.006
R24627 vp_p.n5570 vp_p.n5569 0.006
R24628 vp_p.n5567 vp_p.n5566 0.006
R24629 vp_p.n5556 vp_p.n5555 0.006
R24630 vp_p.n5553 vp_p.n5552 0.006
R24631 vp_p.n5542 vp_p.n5541 0.006
R24632 vp_p.n5539 vp_p.n5538 0.006
R24633 vp_p.n5528 vp_p.n5527 0.006
R24634 vp_p.n5525 vp_p.n5524 0.006
R24635 vp_p.n5514 vp_p.n5513 0.006
R24636 vp_p.n5511 vp_p.n5510 0.006
R24637 vp_p.n5500 vp_p.n5499 0.006
R24638 vp_p.n5497 vp_p.n5496 0.006
R24639 vp_p.n5486 vp_p.n5485 0.006
R24640 vp_p.n5483 vp_p.n5482 0.006
R24641 vp_p.n5472 vp_p.n5471 0.006
R24642 vp_p.n5469 vp_p.n5468 0.006
R24643 vp_p.n5458 vp_p.n5457 0.006
R24644 vp_p.n5455 vp_p.n5454 0.006
R24645 vp_p.n5444 vp_p.n5443 0.006
R24646 vp_p.n5441 vp_p.n5440 0.006
R24647 vp_p.n5430 vp_p.n5429 0.006
R24648 vp_p.n5427 vp_p.n5426 0.006
R24649 vp_p.n5416 vp_p.n5415 0.006
R24650 vp_p.n5413 vp_p.n5412 0.006
R24651 vp_p.n5402 vp_p.n5401 0.006
R24652 vp_p.n5399 vp_p.n5398 0.006
R24653 vp_p.n5388 vp_p.n5387 0.006
R24654 vp_p.n5385 vp_p.n5384 0.006
R24655 vp_p.n5374 vp_p.n5373 0.006
R24656 vp_p.n5371 vp_p.n5370 0.006
R24657 vp_p.n5360 vp_p.n5359 0.006
R24658 vp_p.n5357 vp_p.n5356 0.006
R24659 vp_p.n5346 vp_p.n5345 0.006
R24660 vp_p.n5343 vp_p.n5342 0.006
R24661 vp_p.n5332 vp_p.n5331 0.006
R24662 vp_p.n5329 vp_p.n5328 0.006
R24663 vp_p.n5318 vp_p.n5317 0.006
R24664 vp_p.n5315 vp_p.n5314 0.006
R24665 vp_p.n5304 vp_p.n5303 0.006
R24666 vp_p.n5301 vp_p.n5300 0.006
R24667 vp_p.n5290 vp_p.n5289 0.006
R24668 vp_p.n5287 vp_p.n5286 0.006
R24669 vp_p.n5276 vp_p.n5275 0.006
R24670 vp_p.n5273 vp_p.n5272 0.006
R24671 vp_p.n5262 vp_p.n5261 0.006
R24672 vp_p.n5259 vp_p.n5258 0.006
R24673 vp_p.n5248 vp_p.n5247 0.006
R24674 vp_p.n5245 vp_p.n5244 0.006
R24675 vp_p.n5234 vp_p.n5233 0.006
R24676 vp_p.n5231 vp_p.n5230 0.006
R24677 vp_p.n5220 vp_p.n5219 0.006
R24678 vp_p.n5217 vp_p.n5216 0.006
R24679 vp_p.n5206 vp_p.n5205 0.006
R24680 vp_p.n5203 vp_p.n5202 0.006
R24681 vp_p.n5192 vp_p.n5191 0.006
R24682 vp_p.n5189 vp_p.n5188 0.006
R24683 vp_p.n5178 vp_p.n5177 0.006
R24684 vp_p.n5175 vp_p.n5174 0.006
R24685 vp_p.n5164 vp_p.n5163 0.006
R24686 vp_p.n5161 vp_p.n5160 0.006
R24687 vp_p.n5150 vp_p.n5149 0.006
R24688 vp_p.n5147 vp_p.n5146 0.006
R24689 vp_p.n5136 vp_p.n5135 0.006
R24690 vp_p.n5133 vp_p.n5132 0.006
R24691 vp_p.n5122 vp_p.n5121 0.006
R24692 vp_p.n5119 vp_p.n5118 0.006
R24693 vp_p.n5108 vp_p.n5107 0.006
R24694 vp_p.n5105 vp_p.n5104 0.006
R24695 vp_p.n5094 vp_p.n5093 0.006
R24696 vp_p.n5091 vp_p.n5090 0.006
R24697 vp_p.n5080 vp_p.n5079 0.006
R24698 vp_p.n5077 vp_p.n5076 0.006
R24699 vp_p.n5066 vp_p.n5065 0.006
R24700 vp_p.n5063 vp_p.n5062 0.006
R24701 vp_p.n5052 vp_p.n5051 0.006
R24702 vp_p.n5049 vp_p.n5048 0.006
R24703 vp_p.n5038 vp_p.n5037 0.006
R24704 vp_p.n5035 vp_p.n5034 0.006
R24705 vp_p.n5024 vp_p.n5023 0.006
R24706 vp_p.n5021 vp_p.n5020 0.006
R24707 vp_p.n5010 vp_p.n5009 0.006
R24708 vp_p.n5007 vp_p.n5006 0.006
R24709 vp_p.n4996 vp_p.n4995 0.006
R24710 vp_p.n4993 vp_p.n4992 0.006
R24711 vp_p.n4982 vp_p.n4981 0.006
R24712 vp_p.n4979 vp_p.n4978 0.006
R24713 vp_p.n4968 vp_p.n4967 0.006
R24714 vp_p.n4965 vp_p.n4964 0.006
R24715 vp_p.n4954 vp_p.n4953 0.006
R24716 vp_p.n4951 vp_p.n4950 0.006
R24717 vp_p.n4940 vp_p.n4939 0.006
R24718 vp_p.n4937 vp_p.n4936 0.006
R24719 vp_p.n4926 vp_p.n4925 0.006
R24720 vp_p.n4923 vp_p.n4922 0.006
R24721 vp_p.n4912 vp_p.n4911 0.006
R24722 vp_p.n4909 vp_p.n4908 0.006
R24723 vp_p.n4898 vp_p.n4897 0.006
R24724 vp_p.n4895 vp_p.n4894 0.006
R24725 vp_p.n4884 vp_p.n4883 0.006
R24726 vp_p.n4881 vp_p.n4880 0.006
R24727 vp_p.n4870 vp_p.n4869 0.006
R24728 vp_p.n4867 vp_p.n4866 0.006
R24729 vp_p.n4856 vp_p.n4855 0.006
R24730 vp_p.n4853 vp_p.n4852 0.006
R24731 vp_p.n4842 vp_p.n4841 0.006
R24732 vp_p.n4839 vp_p.n4838 0.006
R24733 vp_p.n4828 vp_p.n4827 0.006
R24734 vp_p.n4825 vp_p.n4824 0.006
R24735 vp_p.n4814 vp_p.n4813 0.006
R24736 vp_p.n4811 vp_p.n4810 0.006
R24737 vp_p.n4800 vp_p.n4799 0.006
R24738 vp_p.n4797 vp_p.n4796 0.006
R24739 vp_p.n4786 vp_p.n4785 0.006
R24740 vp_p.n4783 vp_p.n4782 0.006
R24741 vp_p.n4772 vp_p.n4771 0.006
R24742 vp_p.n4769 vp_p.n4768 0.006
R24743 vp_p.n4758 vp_p.n4757 0.006
R24744 vp_p.n4755 vp_p.n4754 0.006
R24745 vp_p.n4744 vp_p.n4743 0.006
R24746 vp_p.n5752 vp_p.n5751 0.006
R24747 vp_p.n4330 vp_p.n4329 0.006
R24748 vp_p.n2901 vp_p.n2900 0.006
R24749 vp_p.n1471 vp_p.n1470 0.006
R24750 vp_p.n10213 vp_p.n10212 0.006
R24751 vp_p.n11646 vp_p.n11645 0.006
R24752 vp_p.n13080 vp_p.n13079 0.006
R24753 vp_p.n14449 vp_p.n14448 0.006
R24754 vp_p.n15882 vp_p.n15881 0.006
R24755 vp_p.n17314 vp_p.n17313 0.006
R24756 vp_p.n18745 vp_p.n18744 0.006
R24757 vp_p.n20175 vp_p.n20174 0.006
R24758 vp_p.n21604 vp_p.n21603 0.006
R24759 vp_p.n23032 vp_p.n23031 0.006
R24760 vp_p.n23436 vp_p.n23435 0.006
R24761 vp_p.n23441 vp_p.n23440 0.006
R24762 vp_p.n23452 vp_p.n23446 0.006
R24763 vp_p.n23456 vp_p.n23455 0.006
R24764 vp_p.n23466 vp_p.n23460 0.006
R24765 vp_p.n23470 vp_p.n23469 0.006
R24766 vp_p.n23480 vp_p.n23474 0.006
R24767 vp_p.n23484 vp_p.n23483 0.006
R24768 vp_p.n23494 vp_p.n23488 0.006
R24769 vp_p.n23498 vp_p.n23497 0.006
R24770 vp_p.n23508 vp_p.n23502 0.006
R24771 vp_p.n23512 vp_p.n23511 0.006
R24772 vp_p.n23522 vp_p.n23516 0.006
R24773 vp_p.n23526 vp_p.n23525 0.006
R24774 vp_p.n23536 vp_p.n23530 0.006
R24775 vp_p.n23540 vp_p.n23539 0.006
R24776 vp_p.n23550 vp_p.n23544 0.006
R24777 vp_p.n23554 vp_p.n23553 0.006
R24778 vp_p.n23564 vp_p.n23558 0.006
R24779 vp_p.n23568 vp_p.n23567 0.006
R24780 vp_p.n23578 vp_p.n23572 0.006
R24781 vp_p.n23582 vp_p.n23581 0.006
R24782 vp_p.n23592 vp_p.n23586 0.006
R24783 vp_p.n23596 vp_p.n23595 0.006
R24784 vp_p.n23606 vp_p.n23600 0.006
R24785 vp_p.n23610 vp_p.n23609 0.006
R24786 vp_p.n23620 vp_p.n23614 0.006
R24787 vp_p.n23624 vp_p.n23623 0.006
R24788 vp_p.n23634 vp_p.n23628 0.006
R24789 vp_p.n23638 vp_p.n23637 0.006
R24790 vp_p.n23648 vp_p.n23642 0.006
R24791 vp_p.n23652 vp_p.n23651 0.006
R24792 vp_p.n23662 vp_p.n23656 0.006
R24793 vp_p.n23666 vp_p.n23665 0.006
R24794 vp_p.n23676 vp_p.n23670 0.006
R24795 vp_p.n23680 vp_p.n23679 0.006
R24796 vp_p.n23690 vp_p.n23684 0.006
R24797 vp_p.n23694 vp_p.n23693 0.006
R24798 vp_p.n23704 vp_p.n23698 0.006
R24799 vp_p.n23708 vp_p.n23707 0.006
R24800 vp_p.n23718 vp_p.n23712 0.006
R24801 vp_p.n23722 vp_p.n23721 0.006
R24802 vp_p.n23732 vp_p.n23726 0.006
R24803 vp_p.n23736 vp_p.n23735 0.006
R24804 vp_p.n23746 vp_p.n23740 0.006
R24805 vp_p.n23750 vp_p.n23749 0.006
R24806 vp_p.n23760 vp_p.n23754 0.006
R24807 vp_p.n23764 vp_p.n23763 0.006
R24808 vp_p.n23774 vp_p.n23768 0.006
R24809 vp_p.n23778 vp_p.n23777 0.006
R24810 vp_p.n23788 vp_p.n23782 0.006
R24811 vp_p.n23792 vp_p.n23791 0.006
R24812 vp_p.n23802 vp_p.n23796 0.006
R24813 vp_p.n23806 vp_p.n23805 0.006
R24814 vp_p.n23816 vp_p.n23810 0.006
R24815 vp_p.n23820 vp_p.n23819 0.006
R24816 vp_p.n23830 vp_p.n23824 0.006
R24817 vp_p.n23834 vp_p.n23833 0.006
R24818 vp_p.n23844 vp_p.n23838 0.006
R24819 vp_p.n23848 vp_p.n23847 0.006
R24820 vp_p.n23858 vp_p.n23852 0.006
R24821 vp_p.n23862 vp_p.n23861 0.006
R24822 vp_p.n23872 vp_p.n23866 0.006
R24823 vp_p.n23876 vp_p.n23875 0.006
R24824 vp_p.n23886 vp_p.n23880 0.006
R24825 vp_p.n23890 vp_p.n23889 0.006
R24826 vp_p.n23900 vp_p.n23894 0.006
R24827 vp_p.n23904 vp_p.n23903 0.006
R24828 vp_p.n23914 vp_p.n23908 0.006
R24829 vp_p.n23918 vp_p.n23917 0.006
R24830 vp_p.n23928 vp_p.n23922 0.006
R24831 vp_p.n23932 vp_p.n23931 0.006
R24832 vp_p.n23942 vp_p.n23936 0.006
R24833 vp_p.n23946 vp_p.n23945 0.006
R24834 vp_p.n23956 vp_p.n23950 0.006
R24835 vp_p.n23960 vp_p.n23959 0.006
R24836 vp_p.n23970 vp_p.n23964 0.006
R24837 vp_p.n23974 vp_p.n23973 0.006
R24838 vp_p.n23984 vp_p.n23978 0.006
R24839 vp_p.n23988 vp_p.n23987 0.006
R24840 vp_p.n23998 vp_p.n23992 0.006
R24841 vp_p.n24002 vp_p.n24001 0.006
R24842 vp_p.n24012 vp_p.n24006 0.006
R24843 vp_p.n24016 vp_p.n24015 0.006
R24844 vp_p.n24026 vp_p.n24020 0.006
R24845 vp_p.n24030 vp_p.n24029 0.006
R24846 vp_p.n24040 vp_p.n24034 0.006
R24847 vp_p.n24044 vp_p.n24043 0.006
R24848 vp_p.n24054 vp_p.n24048 0.006
R24849 vp_p.n24058 vp_p.n24057 0.006
R24850 vp_p.n24068 vp_p.n24062 0.006
R24851 vp_p.n24072 vp_p.n24071 0.006
R24852 vp_p.n24082 vp_p.n24076 0.006
R24853 vp_p.n24086 vp_p.n24085 0.006
R24854 vp_p.n24096 vp_p.n24090 0.006
R24855 vp_p.n24100 vp_p.n24099 0.006
R24856 vp_p.n24110 vp_p.n24104 0.006
R24857 vp_p.n24114 vp_p.n24113 0.006
R24858 vp_p.n24124 vp_p.n24118 0.006
R24859 vp_p.n24128 vp_p.n24127 0.006
R24860 vp_p.n24138 vp_p.n24132 0.006
R24861 vp_p.n24142 vp_p.n24141 0.006
R24862 vp_p.n24152 vp_p.n24146 0.006
R24863 vp_p.n24156 vp_p.n24155 0.006
R24864 vp_p.n24166 vp_p.n24160 0.006
R24865 vp_p.n24170 vp_p.n24169 0.006
R24866 vp_p.n24180 vp_p.n24174 0.006
R24867 vp_p.n24184 vp_p.n24183 0.006
R24868 vp_p.n24194 vp_p.n24188 0.006
R24869 vp_p.n24198 vp_p.n24197 0.006
R24870 vp_p.n24208 vp_p.n24202 0.006
R24871 vp_p.n24212 vp_p.n24211 0.006
R24872 vp_p.n24222 vp_p.n24216 0.006
R24873 vp_p.n24226 vp_p.n24225 0.006
R24874 vp_p.n24236 vp_p.n24230 0.006
R24875 vp_p.n24240 vp_p.n24239 0.006
R24876 vp_p.n24250 vp_p.n24244 0.006
R24877 vp_p.n24254 vp_p.n24253 0.006
R24878 vp_p.n24264 vp_p.n24258 0.006
R24879 vp_p.n24268 vp_p.n24267 0.006
R24880 vp_p.n24278 vp_p.n24272 0.006
R24881 vp_p.n24282 vp_p.n24281 0.006
R24882 vp_p.n24292 vp_p.n24286 0.006
R24883 vp_p.n24296 vp_p.n24295 0.006
R24884 vp_p.n24306 vp_p.n24300 0.006
R24885 vp_p.n24310 vp_p.n24309 0.006
R24886 vp_p.n24320 vp_p.n24314 0.006
R24887 vp_p.n24324 vp_p.n24323 0.006
R24888 vp_p.n24334 vp_p.n24328 0.006
R24889 vp_p.n24338 vp_p.n24337 0.006
R24890 vp_p.n24348 vp_p.n24342 0.006
R24891 vp_p.n24352 vp_p.n24351 0.006
R24892 vp_p.n24362 vp_p.n24356 0.006
R24893 vp_p.n24366 vp_p.n24365 0.006
R24894 vp_p.n24376 vp_p.n24370 0.006
R24895 vp_p.n24380 vp_p.n24379 0.006
R24896 vp_p.n24390 vp_p.n24384 0.006
R24897 vp_p.n24394 vp_p.n24393 0.006
R24898 vp_p.n24404 vp_p.n24398 0.006
R24899 vp_p.n24408 vp_p.n24407 0.006
R24900 vp_p.n24418 vp_p.n24412 0.006
R24901 vp_p.n24422 vp_p.n24421 0.006
R24902 vp_p.n24432 vp_p.n24426 0.006
R24903 vp_p.n24436 vp_p.n24435 0.006
R24904 vp_p.n24446 vp_p.n24440 0.006
R24905 vp_p.n24450 vp_p.n24449 0.006
R24906 vp_p.n24454 vp_p.n24453 0.006
R24907 vp_p.n24464 vp_p.n24458 0.006
R24908 vp_p.n24468 vp_p.n24467 0.006
R24909 vp_p.n24473 vp_p.n24472 0.006
R24910 vp_p.n24455 vp_p.n24454 0.006
R24911 vp_p.n24451 vp_p.n24450 0.006
R24912 vp_p.n24440 vp_p.n24439 0.006
R24913 vp_p.n24437 vp_p.n24436 0.006
R24914 vp_p.n24426 vp_p.n24425 0.006
R24915 vp_p.n24423 vp_p.n24422 0.006
R24916 vp_p.n24412 vp_p.n24411 0.006
R24917 vp_p.n24409 vp_p.n24408 0.006
R24918 vp_p.n24398 vp_p.n24397 0.006
R24919 vp_p.n24395 vp_p.n24394 0.006
R24920 vp_p.n24384 vp_p.n24383 0.006
R24921 vp_p.n24381 vp_p.n24380 0.006
R24922 vp_p.n24370 vp_p.n24369 0.006
R24923 vp_p.n24367 vp_p.n24366 0.006
R24924 vp_p.n24356 vp_p.n24355 0.006
R24925 vp_p.n24353 vp_p.n24352 0.006
R24926 vp_p.n24342 vp_p.n24341 0.006
R24927 vp_p.n24339 vp_p.n24338 0.006
R24928 vp_p.n24328 vp_p.n24327 0.006
R24929 vp_p.n24325 vp_p.n24324 0.006
R24930 vp_p.n24314 vp_p.n24313 0.006
R24931 vp_p.n24311 vp_p.n24310 0.006
R24932 vp_p.n24300 vp_p.n24299 0.006
R24933 vp_p.n24297 vp_p.n24296 0.006
R24934 vp_p.n24286 vp_p.n24285 0.006
R24935 vp_p.n24283 vp_p.n24282 0.006
R24936 vp_p.n24272 vp_p.n24271 0.006
R24937 vp_p.n24269 vp_p.n24268 0.006
R24938 vp_p.n24258 vp_p.n24257 0.006
R24939 vp_p.n24255 vp_p.n24254 0.006
R24940 vp_p.n24244 vp_p.n24243 0.006
R24941 vp_p.n24241 vp_p.n24240 0.006
R24942 vp_p.n24230 vp_p.n24229 0.006
R24943 vp_p.n24227 vp_p.n24226 0.006
R24944 vp_p.n24216 vp_p.n24215 0.006
R24945 vp_p.n24213 vp_p.n24212 0.006
R24946 vp_p.n24202 vp_p.n24201 0.006
R24947 vp_p.n24199 vp_p.n24198 0.006
R24948 vp_p.n24188 vp_p.n24187 0.006
R24949 vp_p.n24185 vp_p.n24184 0.006
R24950 vp_p.n24174 vp_p.n24173 0.006
R24951 vp_p.n24171 vp_p.n24170 0.006
R24952 vp_p.n24160 vp_p.n24159 0.006
R24953 vp_p.n24157 vp_p.n24156 0.006
R24954 vp_p.n24146 vp_p.n24145 0.006
R24955 vp_p.n24143 vp_p.n24142 0.006
R24956 vp_p.n24132 vp_p.n24131 0.006
R24957 vp_p.n24129 vp_p.n24128 0.006
R24958 vp_p.n24118 vp_p.n24117 0.006
R24959 vp_p.n24115 vp_p.n24114 0.006
R24960 vp_p.n24104 vp_p.n24103 0.006
R24961 vp_p.n24101 vp_p.n24100 0.006
R24962 vp_p.n24090 vp_p.n24089 0.006
R24963 vp_p.n24087 vp_p.n24086 0.006
R24964 vp_p.n24076 vp_p.n24075 0.006
R24965 vp_p.n24073 vp_p.n24072 0.006
R24966 vp_p.n24062 vp_p.n24061 0.006
R24967 vp_p.n24059 vp_p.n24058 0.006
R24968 vp_p.n24048 vp_p.n24047 0.006
R24969 vp_p.n24045 vp_p.n24044 0.006
R24970 vp_p.n24034 vp_p.n24033 0.006
R24971 vp_p.n24031 vp_p.n24030 0.006
R24972 vp_p.n24020 vp_p.n24019 0.006
R24973 vp_p.n24017 vp_p.n24016 0.006
R24974 vp_p.n24006 vp_p.n24005 0.006
R24975 vp_p.n24003 vp_p.n24002 0.006
R24976 vp_p.n23992 vp_p.n23991 0.006
R24977 vp_p.n23989 vp_p.n23988 0.006
R24978 vp_p.n23978 vp_p.n23977 0.006
R24979 vp_p.n23975 vp_p.n23974 0.006
R24980 vp_p.n23964 vp_p.n23963 0.006
R24981 vp_p.n23961 vp_p.n23960 0.006
R24982 vp_p.n23950 vp_p.n23949 0.006
R24983 vp_p.n23947 vp_p.n23946 0.006
R24984 vp_p.n23936 vp_p.n23935 0.006
R24985 vp_p.n23933 vp_p.n23932 0.006
R24986 vp_p.n23922 vp_p.n23921 0.006
R24987 vp_p.n23919 vp_p.n23918 0.006
R24988 vp_p.n23908 vp_p.n23907 0.006
R24989 vp_p.n23905 vp_p.n23904 0.006
R24990 vp_p.n23894 vp_p.n23893 0.006
R24991 vp_p.n23891 vp_p.n23890 0.006
R24992 vp_p.n23880 vp_p.n23879 0.006
R24993 vp_p.n23877 vp_p.n23876 0.006
R24994 vp_p.n23866 vp_p.n23865 0.006
R24995 vp_p.n23863 vp_p.n23862 0.006
R24996 vp_p.n23852 vp_p.n23851 0.006
R24997 vp_p.n23849 vp_p.n23848 0.006
R24998 vp_p.n23838 vp_p.n23837 0.006
R24999 vp_p.n23835 vp_p.n23834 0.006
R25000 vp_p.n23824 vp_p.n23823 0.006
R25001 vp_p.n23821 vp_p.n23820 0.006
R25002 vp_p.n23810 vp_p.n23809 0.006
R25003 vp_p.n23807 vp_p.n23806 0.006
R25004 vp_p.n23796 vp_p.n23795 0.006
R25005 vp_p.n23793 vp_p.n23792 0.006
R25006 vp_p.n23782 vp_p.n23781 0.006
R25007 vp_p.n23779 vp_p.n23778 0.006
R25008 vp_p.n23768 vp_p.n23767 0.006
R25009 vp_p.n23765 vp_p.n23764 0.006
R25010 vp_p.n23754 vp_p.n23753 0.006
R25011 vp_p.n23751 vp_p.n23750 0.006
R25012 vp_p.n23740 vp_p.n23739 0.006
R25013 vp_p.n23737 vp_p.n23736 0.006
R25014 vp_p.n23726 vp_p.n23725 0.006
R25015 vp_p.n23723 vp_p.n23722 0.006
R25016 vp_p.n23712 vp_p.n23711 0.006
R25017 vp_p.n23709 vp_p.n23708 0.006
R25018 vp_p.n23698 vp_p.n23697 0.006
R25019 vp_p.n23695 vp_p.n23694 0.006
R25020 vp_p.n23684 vp_p.n23683 0.006
R25021 vp_p.n23681 vp_p.n23680 0.006
R25022 vp_p.n23670 vp_p.n23669 0.006
R25023 vp_p.n23667 vp_p.n23666 0.006
R25024 vp_p.n23656 vp_p.n23655 0.006
R25025 vp_p.n23653 vp_p.n23652 0.006
R25026 vp_p.n23642 vp_p.n23641 0.006
R25027 vp_p.n23639 vp_p.n23638 0.006
R25028 vp_p.n23628 vp_p.n23627 0.006
R25029 vp_p.n23625 vp_p.n23624 0.006
R25030 vp_p.n23614 vp_p.n23613 0.006
R25031 vp_p.n23611 vp_p.n23610 0.006
R25032 vp_p.n23600 vp_p.n23599 0.006
R25033 vp_p.n23597 vp_p.n23596 0.006
R25034 vp_p.n23586 vp_p.n23585 0.006
R25035 vp_p.n23583 vp_p.n23582 0.006
R25036 vp_p.n23572 vp_p.n23571 0.006
R25037 vp_p.n23569 vp_p.n23568 0.006
R25038 vp_p.n23558 vp_p.n23557 0.006
R25039 vp_p.n23555 vp_p.n23554 0.006
R25040 vp_p.n23544 vp_p.n23543 0.006
R25041 vp_p.n23541 vp_p.n23540 0.006
R25042 vp_p.n23530 vp_p.n23529 0.006
R25043 vp_p.n23527 vp_p.n23526 0.006
R25044 vp_p.n23516 vp_p.n23515 0.006
R25045 vp_p.n23513 vp_p.n23512 0.006
R25046 vp_p.n23502 vp_p.n23501 0.006
R25047 vp_p.n23499 vp_p.n23498 0.006
R25048 vp_p.n23488 vp_p.n23487 0.006
R25049 vp_p.n23485 vp_p.n23484 0.006
R25050 vp_p.n23474 vp_p.n23473 0.006
R25051 vp_p.n23471 vp_p.n23470 0.006
R25052 vp_p.n23460 vp_p.n23459 0.006
R25053 vp_p.n23457 vp_p.n23456 0.006
R25054 vp_p.n23446 vp_p.n23445 0.006
R25055 vp_p.n24458 vp_p.n24457 0.006
R25056 vp_p.n23037 vp_p.n23036 0.006
R25057 vp_p.n21609 vp_p.n21608 0.006
R25058 vp_p.n20180 vp_p.n20179 0.006
R25059 vp_p.n18750 vp_p.n18749 0.006
R25060 vp_p.n17319 vp_p.n17318 0.006
R25061 vp_p.n15887 vp_p.n15886 0.006
R25062 vp_p.n14454 vp_p.n14453 0.006
R25063 vp_p.n13085 vp_p.n13084 0.006
R25064 vp_p.n11651 vp_p.n11650 0.006
R25065 vp_p.n10218 vp_p.n10217 0.006
R25066 vp_p.n1476 vp_p.n1475 0.006
R25067 vp_p.n2906 vp_p.n2905 0.006
R25068 vp_p.n4335 vp_p.n4334 0.006
R25069 vp_p.n5763 vp_p.n5762 0.006
R25070 vp_p.n6157 vp_p.n6156 0.006
R25071 vp_p.n6162 vp_p.n6161 0.006
R25072 vp_p.n6173 vp_p.n6167 0.006
R25073 vp_p.n6177 vp_p.n6176 0.006
R25074 vp_p.n6187 vp_p.n6181 0.006
R25075 vp_p.n6191 vp_p.n6190 0.006
R25076 vp_p.n6201 vp_p.n6195 0.006
R25077 vp_p.n6205 vp_p.n6204 0.006
R25078 vp_p.n6215 vp_p.n6209 0.006
R25079 vp_p.n6219 vp_p.n6218 0.006
R25080 vp_p.n6229 vp_p.n6223 0.006
R25081 vp_p.n6233 vp_p.n6232 0.006
R25082 vp_p.n6243 vp_p.n6237 0.006
R25083 vp_p.n6247 vp_p.n6246 0.006
R25084 vp_p.n6257 vp_p.n6251 0.006
R25085 vp_p.n6261 vp_p.n6260 0.006
R25086 vp_p.n6271 vp_p.n6265 0.006
R25087 vp_p.n6275 vp_p.n6274 0.006
R25088 vp_p.n6285 vp_p.n6279 0.006
R25089 vp_p.n6289 vp_p.n6288 0.006
R25090 vp_p.n6299 vp_p.n6293 0.006
R25091 vp_p.n6303 vp_p.n6302 0.006
R25092 vp_p.n6313 vp_p.n6307 0.006
R25093 vp_p.n6317 vp_p.n6316 0.006
R25094 vp_p.n6327 vp_p.n6321 0.006
R25095 vp_p.n6331 vp_p.n6330 0.006
R25096 vp_p.n6341 vp_p.n6335 0.006
R25097 vp_p.n6345 vp_p.n6344 0.006
R25098 vp_p.n6355 vp_p.n6349 0.006
R25099 vp_p.n6359 vp_p.n6358 0.006
R25100 vp_p.n6369 vp_p.n6363 0.006
R25101 vp_p.n6373 vp_p.n6372 0.006
R25102 vp_p.n6383 vp_p.n6377 0.006
R25103 vp_p.n6387 vp_p.n6386 0.006
R25104 vp_p.n6397 vp_p.n6391 0.006
R25105 vp_p.n6401 vp_p.n6400 0.006
R25106 vp_p.n6411 vp_p.n6405 0.006
R25107 vp_p.n6415 vp_p.n6414 0.006
R25108 vp_p.n6425 vp_p.n6419 0.006
R25109 vp_p.n6429 vp_p.n6428 0.006
R25110 vp_p.n6439 vp_p.n6433 0.006
R25111 vp_p.n6443 vp_p.n6442 0.006
R25112 vp_p.n6453 vp_p.n6447 0.006
R25113 vp_p.n6457 vp_p.n6456 0.006
R25114 vp_p.n6467 vp_p.n6461 0.006
R25115 vp_p.n6471 vp_p.n6470 0.006
R25116 vp_p.n6481 vp_p.n6475 0.006
R25117 vp_p.n6485 vp_p.n6484 0.006
R25118 vp_p.n6495 vp_p.n6489 0.006
R25119 vp_p.n6499 vp_p.n6498 0.006
R25120 vp_p.n6509 vp_p.n6503 0.006
R25121 vp_p.n6513 vp_p.n6512 0.006
R25122 vp_p.n6523 vp_p.n6517 0.006
R25123 vp_p.n6527 vp_p.n6526 0.006
R25124 vp_p.n6537 vp_p.n6531 0.006
R25125 vp_p.n6541 vp_p.n6540 0.006
R25126 vp_p.n6551 vp_p.n6545 0.006
R25127 vp_p.n6555 vp_p.n6554 0.006
R25128 vp_p.n6565 vp_p.n6559 0.006
R25129 vp_p.n6569 vp_p.n6568 0.006
R25130 vp_p.n6579 vp_p.n6573 0.006
R25131 vp_p.n6583 vp_p.n6582 0.006
R25132 vp_p.n6593 vp_p.n6587 0.006
R25133 vp_p.n6597 vp_p.n6596 0.006
R25134 vp_p.n6607 vp_p.n6601 0.006
R25135 vp_p.n6611 vp_p.n6610 0.006
R25136 vp_p.n6621 vp_p.n6615 0.006
R25137 vp_p.n6625 vp_p.n6624 0.006
R25138 vp_p.n6635 vp_p.n6629 0.006
R25139 vp_p.n6639 vp_p.n6638 0.006
R25140 vp_p.n6649 vp_p.n6643 0.006
R25141 vp_p.n6653 vp_p.n6652 0.006
R25142 vp_p.n6663 vp_p.n6657 0.006
R25143 vp_p.n6667 vp_p.n6666 0.006
R25144 vp_p.n6677 vp_p.n6671 0.006
R25145 vp_p.n6681 vp_p.n6680 0.006
R25146 vp_p.n6691 vp_p.n6685 0.006
R25147 vp_p.n6695 vp_p.n6694 0.006
R25148 vp_p.n6705 vp_p.n6699 0.006
R25149 vp_p.n6709 vp_p.n6708 0.006
R25150 vp_p.n6719 vp_p.n6713 0.006
R25151 vp_p.n6723 vp_p.n6722 0.006
R25152 vp_p.n6733 vp_p.n6727 0.006
R25153 vp_p.n6737 vp_p.n6736 0.006
R25154 vp_p.n6747 vp_p.n6741 0.006
R25155 vp_p.n6751 vp_p.n6750 0.006
R25156 vp_p.n6761 vp_p.n6755 0.006
R25157 vp_p.n6765 vp_p.n6764 0.006
R25158 vp_p.n6775 vp_p.n6769 0.006
R25159 vp_p.n6779 vp_p.n6778 0.006
R25160 vp_p.n6789 vp_p.n6783 0.006
R25161 vp_p.n6793 vp_p.n6792 0.006
R25162 vp_p.n6803 vp_p.n6797 0.006
R25163 vp_p.n6807 vp_p.n6806 0.006
R25164 vp_p.n6817 vp_p.n6811 0.006
R25165 vp_p.n6821 vp_p.n6820 0.006
R25166 vp_p.n6831 vp_p.n6825 0.006
R25167 vp_p.n6835 vp_p.n6834 0.006
R25168 vp_p.n6845 vp_p.n6839 0.006
R25169 vp_p.n6849 vp_p.n6848 0.006
R25170 vp_p.n6859 vp_p.n6853 0.006
R25171 vp_p.n6863 vp_p.n6862 0.006
R25172 vp_p.n6873 vp_p.n6867 0.006
R25173 vp_p.n6877 vp_p.n6876 0.006
R25174 vp_p.n6887 vp_p.n6881 0.006
R25175 vp_p.n6891 vp_p.n6890 0.006
R25176 vp_p.n6901 vp_p.n6895 0.006
R25177 vp_p.n6905 vp_p.n6904 0.006
R25178 vp_p.n6915 vp_p.n6909 0.006
R25179 vp_p.n6919 vp_p.n6918 0.006
R25180 vp_p.n6929 vp_p.n6923 0.006
R25181 vp_p.n6933 vp_p.n6932 0.006
R25182 vp_p.n6943 vp_p.n6937 0.006
R25183 vp_p.n6947 vp_p.n6946 0.006
R25184 vp_p.n6957 vp_p.n6951 0.006
R25185 vp_p.n6961 vp_p.n6960 0.006
R25186 vp_p.n6971 vp_p.n6965 0.006
R25187 vp_p.n6975 vp_p.n6974 0.006
R25188 vp_p.n6985 vp_p.n6979 0.006
R25189 vp_p.n6989 vp_p.n6988 0.006
R25190 vp_p.n6999 vp_p.n6993 0.006
R25191 vp_p.n7003 vp_p.n7002 0.006
R25192 vp_p.n7013 vp_p.n7007 0.006
R25193 vp_p.n7017 vp_p.n7016 0.006
R25194 vp_p.n7027 vp_p.n7021 0.006
R25195 vp_p.n7031 vp_p.n7030 0.006
R25196 vp_p.n7041 vp_p.n7035 0.006
R25197 vp_p.n7045 vp_p.n7044 0.006
R25198 vp_p.n7055 vp_p.n7049 0.006
R25199 vp_p.n7059 vp_p.n7058 0.006
R25200 vp_p.n7069 vp_p.n7063 0.006
R25201 vp_p.n7073 vp_p.n7072 0.006
R25202 vp_p.n7083 vp_p.n7077 0.006
R25203 vp_p.n7087 vp_p.n7086 0.006
R25204 vp_p.n7097 vp_p.n7091 0.006
R25205 vp_p.n7101 vp_p.n7100 0.006
R25206 vp_p.n7111 vp_p.n7105 0.006
R25207 vp_p.n7115 vp_p.n7114 0.006
R25208 vp_p.n7125 vp_p.n7119 0.006
R25209 vp_p.n7129 vp_p.n7128 0.006
R25210 vp_p.n7139 vp_p.n7133 0.006
R25211 vp_p.n7143 vp_p.n7142 0.006
R25212 vp_p.n7153 vp_p.n7147 0.006
R25213 vp_p.n7157 vp_p.n7156 0.006
R25214 vp_p.n7167 vp_p.n7161 0.006
R25215 vp_p.n7171 vp_p.n7170 0.006
R25216 vp_p.n7181 vp_p.n7175 0.006
R25217 vp_p.n7185 vp_p.n7184 0.006
R25218 vp_p.n7195 vp_p.n7189 0.006
R25219 vp_p.n7199 vp_p.n7198 0.006
R25220 vp_p.n7186 vp_p.n7185 0.006
R25221 vp_p.n7175 vp_p.n7174 0.006
R25222 vp_p.n7172 vp_p.n7171 0.006
R25223 vp_p.n7161 vp_p.n7160 0.006
R25224 vp_p.n7158 vp_p.n7157 0.006
R25225 vp_p.n7147 vp_p.n7146 0.006
R25226 vp_p.n7144 vp_p.n7143 0.006
R25227 vp_p.n7133 vp_p.n7132 0.006
R25228 vp_p.n7130 vp_p.n7129 0.006
R25229 vp_p.n7119 vp_p.n7118 0.006
R25230 vp_p.n7116 vp_p.n7115 0.006
R25231 vp_p.n7105 vp_p.n7104 0.006
R25232 vp_p.n7102 vp_p.n7101 0.006
R25233 vp_p.n7091 vp_p.n7090 0.006
R25234 vp_p.n7088 vp_p.n7087 0.006
R25235 vp_p.n7077 vp_p.n7076 0.006
R25236 vp_p.n7074 vp_p.n7073 0.006
R25237 vp_p.n7063 vp_p.n7062 0.006
R25238 vp_p.n7060 vp_p.n7059 0.006
R25239 vp_p.n7049 vp_p.n7048 0.006
R25240 vp_p.n7046 vp_p.n7045 0.006
R25241 vp_p.n7035 vp_p.n7034 0.006
R25242 vp_p.n7032 vp_p.n7031 0.006
R25243 vp_p.n7021 vp_p.n7020 0.006
R25244 vp_p.n7018 vp_p.n7017 0.006
R25245 vp_p.n7007 vp_p.n7006 0.006
R25246 vp_p.n7004 vp_p.n7003 0.006
R25247 vp_p.n6993 vp_p.n6992 0.006
R25248 vp_p.n6990 vp_p.n6989 0.006
R25249 vp_p.n6979 vp_p.n6978 0.006
R25250 vp_p.n6976 vp_p.n6975 0.006
R25251 vp_p.n6965 vp_p.n6964 0.006
R25252 vp_p.n6962 vp_p.n6961 0.006
R25253 vp_p.n6951 vp_p.n6950 0.006
R25254 vp_p.n6948 vp_p.n6947 0.006
R25255 vp_p.n6937 vp_p.n6936 0.006
R25256 vp_p.n6934 vp_p.n6933 0.006
R25257 vp_p.n6923 vp_p.n6922 0.006
R25258 vp_p.n6920 vp_p.n6919 0.006
R25259 vp_p.n6909 vp_p.n6908 0.006
R25260 vp_p.n6906 vp_p.n6905 0.006
R25261 vp_p.n6895 vp_p.n6894 0.006
R25262 vp_p.n6892 vp_p.n6891 0.006
R25263 vp_p.n6881 vp_p.n6880 0.006
R25264 vp_p.n6878 vp_p.n6877 0.006
R25265 vp_p.n6867 vp_p.n6866 0.006
R25266 vp_p.n6864 vp_p.n6863 0.006
R25267 vp_p.n6853 vp_p.n6852 0.006
R25268 vp_p.n6850 vp_p.n6849 0.006
R25269 vp_p.n6839 vp_p.n6838 0.006
R25270 vp_p.n6836 vp_p.n6835 0.006
R25271 vp_p.n6825 vp_p.n6824 0.006
R25272 vp_p.n6822 vp_p.n6821 0.006
R25273 vp_p.n6811 vp_p.n6810 0.006
R25274 vp_p.n6808 vp_p.n6807 0.006
R25275 vp_p.n6797 vp_p.n6796 0.006
R25276 vp_p.n6794 vp_p.n6793 0.006
R25277 vp_p.n6783 vp_p.n6782 0.006
R25278 vp_p.n6780 vp_p.n6779 0.006
R25279 vp_p.n6769 vp_p.n6768 0.006
R25280 vp_p.n6766 vp_p.n6765 0.006
R25281 vp_p.n6755 vp_p.n6754 0.006
R25282 vp_p.n6752 vp_p.n6751 0.006
R25283 vp_p.n6741 vp_p.n6740 0.006
R25284 vp_p.n6738 vp_p.n6737 0.006
R25285 vp_p.n6727 vp_p.n6726 0.006
R25286 vp_p.n6724 vp_p.n6723 0.006
R25287 vp_p.n6713 vp_p.n6712 0.006
R25288 vp_p.n6710 vp_p.n6709 0.006
R25289 vp_p.n6699 vp_p.n6698 0.006
R25290 vp_p.n6696 vp_p.n6695 0.006
R25291 vp_p.n6685 vp_p.n6684 0.006
R25292 vp_p.n6682 vp_p.n6681 0.006
R25293 vp_p.n6671 vp_p.n6670 0.006
R25294 vp_p.n6668 vp_p.n6667 0.006
R25295 vp_p.n6657 vp_p.n6656 0.006
R25296 vp_p.n6654 vp_p.n6653 0.006
R25297 vp_p.n6643 vp_p.n6642 0.006
R25298 vp_p.n6640 vp_p.n6639 0.006
R25299 vp_p.n6629 vp_p.n6628 0.006
R25300 vp_p.n6626 vp_p.n6625 0.006
R25301 vp_p.n6615 vp_p.n6614 0.006
R25302 vp_p.n6612 vp_p.n6611 0.006
R25303 vp_p.n6601 vp_p.n6600 0.006
R25304 vp_p.n6598 vp_p.n6597 0.006
R25305 vp_p.n6587 vp_p.n6586 0.006
R25306 vp_p.n6584 vp_p.n6583 0.006
R25307 vp_p.n6573 vp_p.n6572 0.006
R25308 vp_p.n6570 vp_p.n6569 0.006
R25309 vp_p.n6559 vp_p.n6558 0.006
R25310 vp_p.n6556 vp_p.n6555 0.006
R25311 vp_p.n6545 vp_p.n6544 0.006
R25312 vp_p.n6542 vp_p.n6541 0.006
R25313 vp_p.n6531 vp_p.n6530 0.006
R25314 vp_p.n6528 vp_p.n6527 0.006
R25315 vp_p.n6517 vp_p.n6516 0.006
R25316 vp_p.n6514 vp_p.n6513 0.006
R25317 vp_p.n6503 vp_p.n6502 0.006
R25318 vp_p.n6500 vp_p.n6499 0.006
R25319 vp_p.n6489 vp_p.n6488 0.006
R25320 vp_p.n6486 vp_p.n6485 0.006
R25321 vp_p.n6475 vp_p.n6474 0.006
R25322 vp_p.n6472 vp_p.n6471 0.006
R25323 vp_p.n6461 vp_p.n6460 0.006
R25324 vp_p.n6458 vp_p.n6457 0.006
R25325 vp_p.n6447 vp_p.n6446 0.006
R25326 vp_p.n6444 vp_p.n6443 0.006
R25327 vp_p.n6433 vp_p.n6432 0.006
R25328 vp_p.n6430 vp_p.n6429 0.006
R25329 vp_p.n6419 vp_p.n6418 0.006
R25330 vp_p.n6416 vp_p.n6415 0.006
R25331 vp_p.n6405 vp_p.n6404 0.006
R25332 vp_p.n6402 vp_p.n6401 0.006
R25333 vp_p.n6391 vp_p.n6390 0.006
R25334 vp_p.n6388 vp_p.n6387 0.006
R25335 vp_p.n6377 vp_p.n6376 0.006
R25336 vp_p.n6374 vp_p.n6373 0.006
R25337 vp_p.n6363 vp_p.n6362 0.006
R25338 vp_p.n6360 vp_p.n6359 0.006
R25339 vp_p.n6349 vp_p.n6348 0.006
R25340 vp_p.n6346 vp_p.n6345 0.006
R25341 vp_p.n6335 vp_p.n6334 0.006
R25342 vp_p.n6332 vp_p.n6331 0.006
R25343 vp_p.n6321 vp_p.n6320 0.006
R25344 vp_p.n6318 vp_p.n6317 0.006
R25345 vp_p.n6307 vp_p.n6306 0.006
R25346 vp_p.n6304 vp_p.n6303 0.006
R25347 vp_p.n6293 vp_p.n6292 0.006
R25348 vp_p.n6290 vp_p.n6289 0.006
R25349 vp_p.n6279 vp_p.n6278 0.006
R25350 vp_p.n6276 vp_p.n6275 0.006
R25351 vp_p.n6265 vp_p.n6264 0.006
R25352 vp_p.n6262 vp_p.n6261 0.006
R25353 vp_p.n6251 vp_p.n6250 0.006
R25354 vp_p.n6248 vp_p.n6247 0.006
R25355 vp_p.n6237 vp_p.n6236 0.006
R25356 vp_p.n6234 vp_p.n6233 0.006
R25357 vp_p.n6223 vp_p.n6222 0.006
R25358 vp_p.n6220 vp_p.n6219 0.006
R25359 vp_p.n6209 vp_p.n6208 0.006
R25360 vp_p.n6206 vp_p.n6205 0.006
R25361 vp_p.n6195 vp_p.n6194 0.006
R25362 vp_p.n6192 vp_p.n6191 0.006
R25363 vp_p.n6181 vp_p.n6180 0.006
R25364 vp_p.n6178 vp_p.n6177 0.006
R25365 vp_p.n6167 vp_p.n6166 0.006
R25366 vp_p.n7189 vp_p.n7188 0.006
R25367 vp_p.n5768 vp_p.n5767 0.006
R25368 vp_p.n4340 vp_p.n4339 0.006
R25369 vp_p.n2911 vp_p.n2910 0.006
R25370 vp_p.n1481 vp_p.n1480 0.006
R25371 vp_p.n10223 vp_p.n10222 0.006
R25372 vp_p.n11656 vp_p.n11655 0.006
R25373 vp_p.n13090 vp_p.n13089 0.006
R25374 vp_p.n14459 vp_p.n14458 0.006
R25375 vp_p.n15892 vp_p.n15891 0.006
R25376 vp_p.n17324 vp_p.n17323 0.006
R25377 vp_p.n18755 vp_p.n18754 0.006
R25378 vp_p.n20185 vp_p.n20184 0.006
R25379 vp_p.n21614 vp_p.n21613 0.006
R25380 vp_p.n23042 vp_p.n23041 0.006
R25381 vp_p.n24469 vp_p.n24468 0.006
R25382 vp_p.n24858 vp_p.n24857 0.006
R25383 vp_p.n24863 vp_p.n24862 0.006
R25384 vp_p.n24874 vp_p.n24868 0.006
R25385 vp_p.n24878 vp_p.n24877 0.006
R25386 vp_p.n24888 vp_p.n24882 0.006
R25387 vp_p.n24892 vp_p.n24891 0.006
R25388 vp_p.n24902 vp_p.n24896 0.006
R25389 vp_p.n24906 vp_p.n24905 0.006
R25390 vp_p.n24916 vp_p.n24910 0.006
R25391 vp_p.n24920 vp_p.n24919 0.006
R25392 vp_p.n24930 vp_p.n24924 0.006
R25393 vp_p.n24934 vp_p.n24933 0.006
R25394 vp_p.n24944 vp_p.n24938 0.006
R25395 vp_p.n24948 vp_p.n24947 0.006
R25396 vp_p.n24958 vp_p.n24952 0.006
R25397 vp_p.n24962 vp_p.n24961 0.006
R25398 vp_p.n24972 vp_p.n24966 0.006
R25399 vp_p.n24976 vp_p.n24975 0.006
R25400 vp_p.n24986 vp_p.n24980 0.006
R25401 vp_p.n24990 vp_p.n24989 0.006
R25402 vp_p.n25000 vp_p.n24994 0.006
R25403 vp_p.n25004 vp_p.n25003 0.006
R25404 vp_p.n25014 vp_p.n25008 0.006
R25405 vp_p.n25018 vp_p.n25017 0.006
R25406 vp_p.n25028 vp_p.n25022 0.006
R25407 vp_p.n25032 vp_p.n25031 0.006
R25408 vp_p.n25042 vp_p.n25036 0.006
R25409 vp_p.n25046 vp_p.n25045 0.006
R25410 vp_p.n25056 vp_p.n25050 0.006
R25411 vp_p.n25060 vp_p.n25059 0.006
R25412 vp_p.n25070 vp_p.n25064 0.006
R25413 vp_p.n25074 vp_p.n25073 0.006
R25414 vp_p.n25084 vp_p.n25078 0.006
R25415 vp_p.n25088 vp_p.n25087 0.006
R25416 vp_p.n25098 vp_p.n25092 0.006
R25417 vp_p.n25102 vp_p.n25101 0.006
R25418 vp_p.n25112 vp_p.n25106 0.006
R25419 vp_p.n25116 vp_p.n25115 0.006
R25420 vp_p.n25126 vp_p.n25120 0.006
R25421 vp_p.n25130 vp_p.n25129 0.006
R25422 vp_p.n25140 vp_p.n25134 0.006
R25423 vp_p.n25144 vp_p.n25143 0.006
R25424 vp_p.n25154 vp_p.n25148 0.006
R25425 vp_p.n25158 vp_p.n25157 0.006
R25426 vp_p.n25168 vp_p.n25162 0.006
R25427 vp_p.n25172 vp_p.n25171 0.006
R25428 vp_p.n25182 vp_p.n25176 0.006
R25429 vp_p.n25186 vp_p.n25185 0.006
R25430 vp_p.n25196 vp_p.n25190 0.006
R25431 vp_p.n25200 vp_p.n25199 0.006
R25432 vp_p.n25210 vp_p.n25204 0.006
R25433 vp_p.n25214 vp_p.n25213 0.006
R25434 vp_p.n25224 vp_p.n25218 0.006
R25435 vp_p.n25228 vp_p.n25227 0.006
R25436 vp_p.n25238 vp_p.n25232 0.006
R25437 vp_p.n25242 vp_p.n25241 0.006
R25438 vp_p.n25252 vp_p.n25246 0.006
R25439 vp_p.n25256 vp_p.n25255 0.006
R25440 vp_p.n25266 vp_p.n25260 0.006
R25441 vp_p.n25270 vp_p.n25269 0.006
R25442 vp_p.n25280 vp_p.n25274 0.006
R25443 vp_p.n25284 vp_p.n25283 0.006
R25444 vp_p.n25294 vp_p.n25288 0.006
R25445 vp_p.n25298 vp_p.n25297 0.006
R25446 vp_p.n25308 vp_p.n25302 0.006
R25447 vp_p.n25312 vp_p.n25311 0.006
R25448 vp_p.n25322 vp_p.n25316 0.006
R25449 vp_p.n25326 vp_p.n25325 0.006
R25450 vp_p.n25336 vp_p.n25330 0.006
R25451 vp_p.n25340 vp_p.n25339 0.006
R25452 vp_p.n25350 vp_p.n25344 0.006
R25453 vp_p.n25354 vp_p.n25353 0.006
R25454 vp_p.n25364 vp_p.n25358 0.006
R25455 vp_p.n25368 vp_p.n25367 0.006
R25456 vp_p.n25378 vp_p.n25372 0.006
R25457 vp_p.n25382 vp_p.n25381 0.006
R25458 vp_p.n25392 vp_p.n25386 0.006
R25459 vp_p.n25396 vp_p.n25395 0.006
R25460 vp_p.n25406 vp_p.n25400 0.006
R25461 vp_p.n25410 vp_p.n25409 0.006
R25462 vp_p.n25420 vp_p.n25414 0.006
R25463 vp_p.n25424 vp_p.n25423 0.006
R25464 vp_p.n25434 vp_p.n25428 0.006
R25465 vp_p.n25438 vp_p.n25437 0.006
R25466 vp_p.n25448 vp_p.n25442 0.006
R25467 vp_p.n25452 vp_p.n25451 0.006
R25468 vp_p.n25462 vp_p.n25456 0.006
R25469 vp_p.n25466 vp_p.n25465 0.006
R25470 vp_p.n25476 vp_p.n25470 0.006
R25471 vp_p.n25480 vp_p.n25479 0.006
R25472 vp_p.n25490 vp_p.n25484 0.006
R25473 vp_p.n25494 vp_p.n25493 0.006
R25474 vp_p.n25504 vp_p.n25498 0.006
R25475 vp_p.n25508 vp_p.n25507 0.006
R25476 vp_p.n25518 vp_p.n25512 0.006
R25477 vp_p.n25522 vp_p.n25521 0.006
R25478 vp_p.n25532 vp_p.n25526 0.006
R25479 vp_p.n25536 vp_p.n25535 0.006
R25480 vp_p.n25546 vp_p.n25540 0.006
R25481 vp_p.n25550 vp_p.n25549 0.006
R25482 vp_p.n25560 vp_p.n25554 0.006
R25483 vp_p.n25564 vp_p.n25563 0.006
R25484 vp_p.n25574 vp_p.n25568 0.006
R25485 vp_p.n25578 vp_p.n25577 0.006
R25486 vp_p.n25588 vp_p.n25582 0.006
R25487 vp_p.n25592 vp_p.n25591 0.006
R25488 vp_p.n25602 vp_p.n25596 0.006
R25489 vp_p.n25606 vp_p.n25605 0.006
R25490 vp_p.n25616 vp_p.n25610 0.006
R25491 vp_p.n25620 vp_p.n25619 0.006
R25492 vp_p.n25630 vp_p.n25624 0.006
R25493 vp_p.n25634 vp_p.n25633 0.006
R25494 vp_p.n25644 vp_p.n25638 0.006
R25495 vp_p.n25648 vp_p.n25647 0.006
R25496 vp_p.n25658 vp_p.n25652 0.006
R25497 vp_p.n25662 vp_p.n25661 0.006
R25498 vp_p.n25672 vp_p.n25666 0.006
R25499 vp_p.n25676 vp_p.n25675 0.006
R25500 vp_p.n25686 vp_p.n25680 0.006
R25501 vp_p.n25690 vp_p.n25689 0.006
R25502 vp_p.n25700 vp_p.n25694 0.006
R25503 vp_p.n25704 vp_p.n25703 0.006
R25504 vp_p.n25714 vp_p.n25708 0.006
R25505 vp_p.n25718 vp_p.n25717 0.006
R25506 vp_p.n25728 vp_p.n25722 0.006
R25507 vp_p.n25732 vp_p.n25731 0.006
R25508 vp_p.n25742 vp_p.n25736 0.006
R25509 vp_p.n25746 vp_p.n25745 0.006
R25510 vp_p.n25756 vp_p.n25750 0.006
R25511 vp_p.n25760 vp_p.n25759 0.006
R25512 vp_p.n25770 vp_p.n25764 0.006
R25513 vp_p.n25774 vp_p.n25773 0.006
R25514 vp_p.n25784 vp_p.n25778 0.006
R25515 vp_p.n25788 vp_p.n25787 0.006
R25516 vp_p.n25798 vp_p.n25792 0.006
R25517 vp_p.n25802 vp_p.n25801 0.006
R25518 vp_p.n25812 vp_p.n25806 0.006
R25519 vp_p.n25816 vp_p.n25815 0.006
R25520 vp_p.n25826 vp_p.n25820 0.006
R25521 vp_p.n25830 vp_p.n25829 0.006
R25522 vp_p.n25840 vp_p.n25834 0.006
R25523 vp_p.n25844 vp_p.n25843 0.006
R25524 vp_p.n25854 vp_p.n25848 0.006
R25525 vp_p.n25858 vp_p.n25857 0.006
R25526 vp_p.n25868 vp_p.n25862 0.006
R25527 vp_p.n25872 vp_p.n25871 0.006
R25528 vp_p.n25882 vp_p.n25876 0.006
R25529 vp_p.n25886 vp_p.n25885 0.006
R25530 vp_p.n25890 vp_p.n25889 0.006
R25531 vp_p.n25900 vp_p.n25894 0.006
R25532 vp_p.n25891 vp_p.n25890 0.006
R25533 vp_p.n25887 vp_p.n25886 0.006
R25534 vp_p.n25876 vp_p.n25875 0.006
R25535 vp_p.n25873 vp_p.n25872 0.006
R25536 vp_p.n25862 vp_p.n25861 0.006
R25537 vp_p.n25859 vp_p.n25858 0.006
R25538 vp_p.n25848 vp_p.n25847 0.006
R25539 vp_p.n25845 vp_p.n25844 0.006
R25540 vp_p.n25834 vp_p.n25833 0.006
R25541 vp_p.n25831 vp_p.n25830 0.006
R25542 vp_p.n25820 vp_p.n25819 0.006
R25543 vp_p.n25817 vp_p.n25816 0.006
R25544 vp_p.n25806 vp_p.n25805 0.006
R25545 vp_p.n25803 vp_p.n25802 0.006
R25546 vp_p.n25792 vp_p.n25791 0.006
R25547 vp_p.n25789 vp_p.n25788 0.006
R25548 vp_p.n25778 vp_p.n25777 0.006
R25549 vp_p.n25775 vp_p.n25774 0.006
R25550 vp_p.n25764 vp_p.n25763 0.006
R25551 vp_p.n25761 vp_p.n25760 0.006
R25552 vp_p.n25750 vp_p.n25749 0.006
R25553 vp_p.n25747 vp_p.n25746 0.006
R25554 vp_p.n25736 vp_p.n25735 0.006
R25555 vp_p.n25733 vp_p.n25732 0.006
R25556 vp_p.n25722 vp_p.n25721 0.006
R25557 vp_p.n25719 vp_p.n25718 0.006
R25558 vp_p.n25708 vp_p.n25707 0.006
R25559 vp_p.n25705 vp_p.n25704 0.006
R25560 vp_p.n25694 vp_p.n25693 0.006
R25561 vp_p.n25691 vp_p.n25690 0.006
R25562 vp_p.n25680 vp_p.n25679 0.006
R25563 vp_p.n25677 vp_p.n25676 0.006
R25564 vp_p.n25666 vp_p.n25665 0.006
R25565 vp_p.n25663 vp_p.n25662 0.006
R25566 vp_p.n25652 vp_p.n25651 0.006
R25567 vp_p.n25649 vp_p.n25648 0.006
R25568 vp_p.n25638 vp_p.n25637 0.006
R25569 vp_p.n25635 vp_p.n25634 0.006
R25570 vp_p.n25624 vp_p.n25623 0.006
R25571 vp_p.n25621 vp_p.n25620 0.006
R25572 vp_p.n25610 vp_p.n25609 0.006
R25573 vp_p.n25607 vp_p.n25606 0.006
R25574 vp_p.n25596 vp_p.n25595 0.006
R25575 vp_p.n25593 vp_p.n25592 0.006
R25576 vp_p.n25582 vp_p.n25581 0.006
R25577 vp_p.n25579 vp_p.n25578 0.006
R25578 vp_p.n25568 vp_p.n25567 0.006
R25579 vp_p.n25565 vp_p.n25564 0.006
R25580 vp_p.n25554 vp_p.n25553 0.006
R25581 vp_p.n25551 vp_p.n25550 0.006
R25582 vp_p.n25540 vp_p.n25539 0.006
R25583 vp_p.n25537 vp_p.n25536 0.006
R25584 vp_p.n25526 vp_p.n25525 0.006
R25585 vp_p.n25523 vp_p.n25522 0.006
R25586 vp_p.n25512 vp_p.n25511 0.006
R25587 vp_p.n25509 vp_p.n25508 0.006
R25588 vp_p.n25498 vp_p.n25497 0.006
R25589 vp_p.n25495 vp_p.n25494 0.006
R25590 vp_p.n25484 vp_p.n25483 0.006
R25591 vp_p.n25481 vp_p.n25480 0.006
R25592 vp_p.n25470 vp_p.n25469 0.006
R25593 vp_p.n25467 vp_p.n25466 0.006
R25594 vp_p.n25456 vp_p.n25455 0.006
R25595 vp_p.n25453 vp_p.n25452 0.006
R25596 vp_p.n25442 vp_p.n25441 0.006
R25597 vp_p.n25439 vp_p.n25438 0.006
R25598 vp_p.n25428 vp_p.n25427 0.006
R25599 vp_p.n25425 vp_p.n25424 0.006
R25600 vp_p.n25414 vp_p.n25413 0.006
R25601 vp_p.n25411 vp_p.n25410 0.006
R25602 vp_p.n25400 vp_p.n25399 0.006
R25603 vp_p.n25397 vp_p.n25396 0.006
R25604 vp_p.n25386 vp_p.n25385 0.006
R25605 vp_p.n25383 vp_p.n25382 0.006
R25606 vp_p.n25372 vp_p.n25371 0.006
R25607 vp_p.n25369 vp_p.n25368 0.006
R25608 vp_p.n25358 vp_p.n25357 0.006
R25609 vp_p.n25355 vp_p.n25354 0.006
R25610 vp_p.n25344 vp_p.n25343 0.006
R25611 vp_p.n25341 vp_p.n25340 0.006
R25612 vp_p.n25330 vp_p.n25329 0.006
R25613 vp_p.n25327 vp_p.n25326 0.006
R25614 vp_p.n25316 vp_p.n25315 0.006
R25615 vp_p.n25313 vp_p.n25312 0.006
R25616 vp_p.n25302 vp_p.n25301 0.006
R25617 vp_p.n25299 vp_p.n25298 0.006
R25618 vp_p.n25288 vp_p.n25287 0.006
R25619 vp_p.n25285 vp_p.n25284 0.006
R25620 vp_p.n25274 vp_p.n25273 0.006
R25621 vp_p.n25271 vp_p.n25270 0.006
R25622 vp_p.n25260 vp_p.n25259 0.006
R25623 vp_p.n25257 vp_p.n25256 0.006
R25624 vp_p.n25246 vp_p.n25245 0.006
R25625 vp_p.n25243 vp_p.n25242 0.006
R25626 vp_p.n25232 vp_p.n25231 0.006
R25627 vp_p.n25229 vp_p.n25228 0.006
R25628 vp_p.n25218 vp_p.n25217 0.006
R25629 vp_p.n25215 vp_p.n25214 0.006
R25630 vp_p.n25204 vp_p.n25203 0.006
R25631 vp_p.n25201 vp_p.n25200 0.006
R25632 vp_p.n25190 vp_p.n25189 0.006
R25633 vp_p.n25187 vp_p.n25186 0.006
R25634 vp_p.n25176 vp_p.n25175 0.006
R25635 vp_p.n25173 vp_p.n25172 0.006
R25636 vp_p.n25162 vp_p.n25161 0.006
R25637 vp_p.n25159 vp_p.n25158 0.006
R25638 vp_p.n25148 vp_p.n25147 0.006
R25639 vp_p.n25145 vp_p.n25144 0.006
R25640 vp_p.n25134 vp_p.n25133 0.006
R25641 vp_p.n25131 vp_p.n25130 0.006
R25642 vp_p.n25120 vp_p.n25119 0.006
R25643 vp_p.n25117 vp_p.n25116 0.006
R25644 vp_p.n25106 vp_p.n25105 0.006
R25645 vp_p.n25103 vp_p.n25102 0.006
R25646 vp_p.n25092 vp_p.n25091 0.006
R25647 vp_p.n25089 vp_p.n25088 0.006
R25648 vp_p.n25078 vp_p.n25077 0.006
R25649 vp_p.n25075 vp_p.n25074 0.006
R25650 vp_p.n25064 vp_p.n25063 0.006
R25651 vp_p.n25061 vp_p.n25060 0.006
R25652 vp_p.n25050 vp_p.n25049 0.006
R25653 vp_p.n25047 vp_p.n25046 0.006
R25654 vp_p.n25036 vp_p.n25035 0.006
R25655 vp_p.n25033 vp_p.n25032 0.006
R25656 vp_p.n25022 vp_p.n25021 0.006
R25657 vp_p.n25019 vp_p.n25018 0.006
R25658 vp_p.n25008 vp_p.n25007 0.006
R25659 vp_p.n25005 vp_p.n25004 0.006
R25660 vp_p.n24994 vp_p.n24993 0.006
R25661 vp_p.n24991 vp_p.n24990 0.006
R25662 vp_p.n24980 vp_p.n24979 0.006
R25663 vp_p.n24977 vp_p.n24976 0.006
R25664 vp_p.n24966 vp_p.n24965 0.006
R25665 vp_p.n24963 vp_p.n24962 0.006
R25666 vp_p.n24952 vp_p.n24951 0.006
R25667 vp_p.n24949 vp_p.n24948 0.006
R25668 vp_p.n24938 vp_p.n24937 0.006
R25669 vp_p.n24935 vp_p.n24934 0.006
R25670 vp_p.n24924 vp_p.n24923 0.006
R25671 vp_p.n24921 vp_p.n24920 0.006
R25672 vp_p.n24910 vp_p.n24909 0.006
R25673 vp_p.n24907 vp_p.n24906 0.006
R25674 vp_p.n24896 vp_p.n24895 0.006
R25675 vp_p.n24893 vp_p.n24892 0.006
R25676 vp_p.n24882 vp_p.n24881 0.006
R25677 vp_p.n24879 vp_p.n24878 0.006
R25678 vp_p.n24868 vp_p.n24867 0.006
R25679 vp_p.n25894 vp_p.n25893 0.006
R25680 vp_p.n24474 vp_p.n24473 0.006
R25681 vp_p.n23047 vp_p.n23046 0.006
R25682 vp_p.n21619 vp_p.n21618 0.006
R25683 vp_p.n20190 vp_p.n20189 0.006
R25684 vp_p.n18760 vp_p.n18759 0.006
R25685 vp_p.n17329 vp_p.n17328 0.006
R25686 vp_p.n15897 vp_p.n15896 0.006
R25687 vp_p.n14464 vp_p.n14463 0.006
R25688 vp_p.n13095 vp_p.n13094 0.006
R25689 vp_p.n11661 vp_p.n11660 0.006
R25690 vp_p.n10228 vp_p.n10227 0.006
R25691 vp_p.n1486 vp_p.n1485 0.006
R25692 vp_p.n2916 vp_p.n2915 0.006
R25693 vp_p.n4345 vp_p.n4344 0.006
R25694 vp_p.n5773 vp_p.n5772 0.006
R25695 vp_p.n7200 vp_p.n7199 0.006
R25696 vp_p.n7574 vp_p.n7573 0.006
R25697 vp_p.n7585 vp_p.n7579 0.006
R25698 vp_p.n7595 vp_p.n7589 0.006
R25699 vp_p.n7599 vp_p.n7598 0.006
R25700 vp_p.n7609 vp_p.n7603 0.006
R25701 vp_p.n7613 vp_p.n7612 0.006
R25702 vp_p.n7623 vp_p.n7617 0.006
R25703 vp_p.n7627 vp_p.n7626 0.006
R25704 vp_p.n7637 vp_p.n7631 0.006
R25705 vp_p.n7641 vp_p.n7640 0.006
R25706 vp_p.n7651 vp_p.n7645 0.006
R25707 vp_p.n7655 vp_p.n7654 0.006
R25708 vp_p.n7665 vp_p.n7659 0.006
R25709 vp_p.n7669 vp_p.n7668 0.006
R25710 vp_p.n7679 vp_p.n7673 0.006
R25711 vp_p.n7683 vp_p.n7682 0.006
R25712 vp_p.n7693 vp_p.n7687 0.006
R25713 vp_p.n7697 vp_p.n7696 0.006
R25714 vp_p.n7707 vp_p.n7701 0.006
R25715 vp_p.n7711 vp_p.n7710 0.006
R25716 vp_p.n7721 vp_p.n7715 0.006
R25717 vp_p.n7725 vp_p.n7724 0.006
R25718 vp_p.n7735 vp_p.n7729 0.006
R25719 vp_p.n7739 vp_p.n7738 0.006
R25720 vp_p.n7749 vp_p.n7743 0.006
R25721 vp_p.n7753 vp_p.n7752 0.006
R25722 vp_p.n7763 vp_p.n7757 0.006
R25723 vp_p.n7767 vp_p.n7766 0.006
R25724 vp_p.n7777 vp_p.n7771 0.006
R25725 vp_p.n7781 vp_p.n7780 0.006
R25726 vp_p.n7791 vp_p.n7785 0.006
R25727 vp_p.n7795 vp_p.n7794 0.006
R25728 vp_p.n7805 vp_p.n7799 0.006
R25729 vp_p.n7809 vp_p.n7808 0.006
R25730 vp_p.n7819 vp_p.n7813 0.006
R25731 vp_p.n7823 vp_p.n7822 0.006
R25732 vp_p.n7833 vp_p.n7827 0.006
R25733 vp_p.n7837 vp_p.n7836 0.006
R25734 vp_p.n7847 vp_p.n7841 0.006
R25735 vp_p.n7851 vp_p.n7850 0.006
R25736 vp_p.n7861 vp_p.n7855 0.006
R25737 vp_p.n7865 vp_p.n7864 0.006
R25738 vp_p.n7875 vp_p.n7869 0.006
R25739 vp_p.n7879 vp_p.n7878 0.006
R25740 vp_p.n7889 vp_p.n7883 0.006
R25741 vp_p.n7893 vp_p.n7892 0.006
R25742 vp_p.n7903 vp_p.n7897 0.006
R25743 vp_p.n7907 vp_p.n7906 0.006
R25744 vp_p.n7917 vp_p.n7911 0.006
R25745 vp_p.n7921 vp_p.n7920 0.006
R25746 vp_p.n7931 vp_p.n7925 0.006
R25747 vp_p.n7935 vp_p.n7934 0.006
R25748 vp_p.n7945 vp_p.n7939 0.006
R25749 vp_p.n7949 vp_p.n7948 0.006
R25750 vp_p.n7959 vp_p.n7953 0.006
R25751 vp_p.n7963 vp_p.n7962 0.006
R25752 vp_p.n7973 vp_p.n7967 0.006
R25753 vp_p.n7977 vp_p.n7976 0.006
R25754 vp_p.n7987 vp_p.n7981 0.006
R25755 vp_p.n7991 vp_p.n7990 0.006
R25756 vp_p.n8001 vp_p.n7995 0.006
R25757 vp_p.n8005 vp_p.n8004 0.006
R25758 vp_p.n8015 vp_p.n8009 0.006
R25759 vp_p.n8019 vp_p.n8018 0.006
R25760 vp_p.n8029 vp_p.n8023 0.006
R25761 vp_p.n8033 vp_p.n8032 0.006
R25762 vp_p.n8043 vp_p.n8037 0.006
R25763 vp_p.n8047 vp_p.n8046 0.006
R25764 vp_p.n8057 vp_p.n8051 0.006
R25765 vp_p.n8061 vp_p.n8060 0.006
R25766 vp_p.n8071 vp_p.n8065 0.006
R25767 vp_p.n8075 vp_p.n8074 0.006
R25768 vp_p.n8085 vp_p.n8079 0.006
R25769 vp_p.n8089 vp_p.n8088 0.006
R25770 vp_p.n8099 vp_p.n8093 0.006
R25771 vp_p.n8103 vp_p.n8102 0.006
R25772 vp_p.n8113 vp_p.n8107 0.006
R25773 vp_p.n8117 vp_p.n8116 0.006
R25774 vp_p.n8127 vp_p.n8121 0.006
R25775 vp_p.n8131 vp_p.n8130 0.006
R25776 vp_p.n8141 vp_p.n8135 0.006
R25777 vp_p.n8145 vp_p.n8144 0.006
R25778 vp_p.n8155 vp_p.n8149 0.006
R25779 vp_p.n8159 vp_p.n8158 0.006
R25780 vp_p.n8169 vp_p.n8163 0.006
R25781 vp_p.n8173 vp_p.n8172 0.006
R25782 vp_p.n8183 vp_p.n8177 0.006
R25783 vp_p.n8187 vp_p.n8186 0.006
R25784 vp_p.n8197 vp_p.n8191 0.006
R25785 vp_p.n8201 vp_p.n8200 0.006
R25786 vp_p.n8211 vp_p.n8205 0.006
R25787 vp_p.n8215 vp_p.n8214 0.006
R25788 vp_p.n8225 vp_p.n8219 0.006
R25789 vp_p.n8229 vp_p.n8228 0.006
R25790 vp_p.n8239 vp_p.n8233 0.006
R25791 vp_p.n8243 vp_p.n8242 0.006
R25792 vp_p.n8253 vp_p.n8247 0.006
R25793 vp_p.n8257 vp_p.n8256 0.006
R25794 vp_p.n8267 vp_p.n8261 0.006
R25795 vp_p.n8271 vp_p.n8270 0.006
R25796 vp_p.n8281 vp_p.n8275 0.006
R25797 vp_p.n8285 vp_p.n8284 0.006
R25798 vp_p.n8295 vp_p.n8289 0.006
R25799 vp_p.n8299 vp_p.n8298 0.006
R25800 vp_p.n8309 vp_p.n8303 0.006
R25801 vp_p.n8313 vp_p.n8312 0.006
R25802 vp_p.n8323 vp_p.n8317 0.006
R25803 vp_p.n8327 vp_p.n8326 0.006
R25804 vp_p.n8337 vp_p.n8331 0.006
R25805 vp_p.n8341 vp_p.n8340 0.006
R25806 vp_p.n8351 vp_p.n8345 0.006
R25807 vp_p.n8355 vp_p.n8354 0.006
R25808 vp_p.n8365 vp_p.n8359 0.006
R25809 vp_p.n8369 vp_p.n8368 0.006
R25810 vp_p.n8379 vp_p.n8373 0.006
R25811 vp_p.n8383 vp_p.n8382 0.006
R25812 vp_p.n8393 vp_p.n8387 0.006
R25813 vp_p.n8397 vp_p.n8396 0.006
R25814 vp_p.n8407 vp_p.n8401 0.006
R25815 vp_p.n8411 vp_p.n8410 0.006
R25816 vp_p.n8421 vp_p.n8415 0.006
R25817 vp_p.n8425 vp_p.n8424 0.006
R25818 vp_p.n8435 vp_p.n8429 0.006
R25819 vp_p.n8439 vp_p.n8438 0.006
R25820 vp_p.n8449 vp_p.n8443 0.006
R25821 vp_p.n8453 vp_p.n8452 0.006
R25822 vp_p.n8463 vp_p.n8457 0.006
R25823 vp_p.n8467 vp_p.n8466 0.006
R25824 vp_p.n8477 vp_p.n8471 0.006
R25825 vp_p.n8481 vp_p.n8480 0.006
R25826 vp_p.n8491 vp_p.n8485 0.006
R25827 vp_p.n8495 vp_p.n8494 0.006
R25828 vp_p.n8505 vp_p.n8499 0.006
R25829 vp_p.n8509 vp_p.n8508 0.006
R25830 vp_p.n8519 vp_p.n8513 0.006
R25831 vp_p.n8523 vp_p.n8522 0.006
R25832 vp_p.n8533 vp_p.n8527 0.006
R25833 vp_p.n8537 vp_p.n8536 0.006
R25834 vp_p.n8547 vp_p.n8541 0.006
R25835 vp_p.n8551 vp_p.n8550 0.006
R25836 vp_p.n8561 vp_p.n8555 0.006
R25837 vp_p.n8565 vp_p.n8564 0.006
R25838 vp_p.n8575 vp_p.n8569 0.006
R25839 vp_p.n8579 vp_p.n8578 0.006
R25840 vp_p.n8589 vp_p.n8583 0.006
R25841 vp_p.n8593 vp_p.n8592 0.006
R25842 vp_p.n8603 vp_p.n8597 0.006
R25843 vp_p.n8607 vp_p.n8606 0.006
R25844 vp_p.n8617 vp_p.n8611 0.006
R25845 vp_p.n7589 vp_p.n7588 0.006
R25846 vp_p.n7600 vp_p.n7599 0.006
R25847 vp_p.n7603 vp_p.n7602 0.006
R25848 vp_p.n7614 vp_p.n7613 0.006
R25849 vp_p.n7617 vp_p.n7616 0.006
R25850 vp_p.n7628 vp_p.n7627 0.006
R25851 vp_p.n7631 vp_p.n7630 0.006
R25852 vp_p.n7642 vp_p.n7641 0.006
R25853 vp_p.n7645 vp_p.n7644 0.006
R25854 vp_p.n7656 vp_p.n7655 0.006
R25855 vp_p.n7659 vp_p.n7658 0.006
R25856 vp_p.n7670 vp_p.n7669 0.006
R25857 vp_p.n7673 vp_p.n7672 0.006
R25858 vp_p.n7684 vp_p.n7683 0.006
R25859 vp_p.n7687 vp_p.n7686 0.006
R25860 vp_p.n7698 vp_p.n7697 0.006
R25861 vp_p.n7701 vp_p.n7700 0.006
R25862 vp_p.n7712 vp_p.n7711 0.006
R25863 vp_p.n7715 vp_p.n7714 0.006
R25864 vp_p.n7726 vp_p.n7725 0.006
R25865 vp_p.n7729 vp_p.n7728 0.006
R25866 vp_p.n7740 vp_p.n7739 0.006
R25867 vp_p.n7743 vp_p.n7742 0.006
R25868 vp_p.n7754 vp_p.n7753 0.006
R25869 vp_p.n7757 vp_p.n7756 0.006
R25870 vp_p.n7768 vp_p.n7767 0.006
R25871 vp_p.n7771 vp_p.n7770 0.006
R25872 vp_p.n7782 vp_p.n7781 0.006
R25873 vp_p.n7785 vp_p.n7784 0.006
R25874 vp_p.n7796 vp_p.n7795 0.006
R25875 vp_p.n7799 vp_p.n7798 0.006
R25876 vp_p.n7810 vp_p.n7809 0.006
R25877 vp_p.n7813 vp_p.n7812 0.006
R25878 vp_p.n7824 vp_p.n7823 0.006
R25879 vp_p.n7827 vp_p.n7826 0.006
R25880 vp_p.n7838 vp_p.n7837 0.006
R25881 vp_p.n7841 vp_p.n7840 0.006
R25882 vp_p.n7852 vp_p.n7851 0.006
R25883 vp_p.n7855 vp_p.n7854 0.006
R25884 vp_p.n7866 vp_p.n7865 0.006
R25885 vp_p.n7869 vp_p.n7868 0.006
R25886 vp_p.n7880 vp_p.n7879 0.006
R25887 vp_p.n7883 vp_p.n7882 0.006
R25888 vp_p.n7894 vp_p.n7893 0.006
R25889 vp_p.n7897 vp_p.n7896 0.006
R25890 vp_p.n7908 vp_p.n7907 0.006
R25891 vp_p.n7911 vp_p.n7910 0.006
R25892 vp_p.n7922 vp_p.n7921 0.006
R25893 vp_p.n7925 vp_p.n7924 0.006
R25894 vp_p.n7936 vp_p.n7935 0.006
R25895 vp_p.n7939 vp_p.n7938 0.006
R25896 vp_p.n7950 vp_p.n7949 0.006
R25897 vp_p.n7953 vp_p.n7952 0.006
R25898 vp_p.n7964 vp_p.n7963 0.006
R25899 vp_p.n7967 vp_p.n7966 0.006
R25900 vp_p.n7978 vp_p.n7977 0.006
R25901 vp_p.n7981 vp_p.n7980 0.006
R25902 vp_p.n7992 vp_p.n7991 0.006
R25903 vp_p.n7995 vp_p.n7994 0.006
R25904 vp_p.n8006 vp_p.n8005 0.006
R25905 vp_p.n8009 vp_p.n8008 0.006
R25906 vp_p.n8020 vp_p.n8019 0.006
R25907 vp_p.n8023 vp_p.n8022 0.006
R25908 vp_p.n8034 vp_p.n8033 0.006
R25909 vp_p.n8037 vp_p.n8036 0.006
R25910 vp_p.n8048 vp_p.n8047 0.006
R25911 vp_p.n8051 vp_p.n8050 0.006
R25912 vp_p.n8062 vp_p.n8061 0.006
R25913 vp_p.n8065 vp_p.n8064 0.006
R25914 vp_p.n8076 vp_p.n8075 0.006
R25915 vp_p.n8079 vp_p.n8078 0.006
R25916 vp_p.n8090 vp_p.n8089 0.006
R25917 vp_p.n8093 vp_p.n8092 0.006
R25918 vp_p.n8104 vp_p.n8103 0.006
R25919 vp_p.n8107 vp_p.n8106 0.006
R25920 vp_p.n8118 vp_p.n8117 0.006
R25921 vp_p.n8121 vp_p.n8120 0.006
R25922 vp_p.n8132 vp_p.n8131 0.006
R25923 vp_p.n8135 vp_p.n8134 0.006
R25924 vp_p.n8146 vp_p.n8145 0.006
R25925 vp_p.n8149 vp_p.n8148 0.006
R25926 vp_p.n8160 vp_p.n8159 0.006
R25927 vp_p.n8163 vp_p.n8162 0.006
R25928 vp_p.n8174 vp_p.n8173 0.006
R25929 vp_p.n8177 vp_p.n8176 0.006
R25930 vp_p.n8188 vp_p.n8187 0.006
R25931 vp_p.n8191 vp_p.n8190 0.006
R25932 vp_p.n8202 vp_p.n8201 0.006
R25933 vp_p.n8205 vp_p.n8204 0.006
R25934 vp_p.n8216 vp_p.n8215 0.006
R25935 vp_p.n8219 vp_p.n8218 0.006
R25936 vp_p.n8230 vp_p.n8229 0.006
R25937 vp_p.n8233 vp_p.n8232 0.006
R25938 vp_p.n8244 vp_p.n8243 0.006
R25939 vp_p.n8247 vp_p.n8246 0.006
R25940 vp_p.n8258 vp_p.n8257 0.006
R25941 vp_p.n8261 vp_p.n8260 0.006
R25942 vp_p.n8272 vp_p.n8271 0.006
R25943 vp_p.n8275 vp_p.n8274 0.006
R25944 vp_p.n8286 vp_p.n8285 0.006
R25945 vp_p.n8289 vp_p.n8288 0.006
R25946 vp_p.n8300 vp_p.n8299 0.006
R25947 vp_p.n8303 vp_p.n8302 0.006
R25948 vp_p.n8314 vp_p.n8313 0.006
R25949 vp_p.n8317 vp_p.n8316 0.006
R25950 vp_p.n8328 vp_p.n8327 0.006
R25951 vp_p.n8331 vp_p.n8330 0.006
R25952 vp_p.n8342 vp_p.n8341 0.006
R25953 vp_p.n8345 vp_p.n8344 0.006
R25954 vp_p.n8356 vp_p.n8355 0.006
R25955 vp_p.n8359 vp_p.n8358 0.006
R25956 vp_p.n8370 vp_p.n8369 0.006
R25957 vp_p.n8373 vp_p.n8372 0.006
R25958 vp_p.n8384 vp_p.n8383 0.006
R25959 vp_p.n8387 vp_p.n8386 0.006
R25960 vp_p.n8398 vp_p.n8397 0.006
R25961 vp_p.n8401 vp_p.n8400 0.006
R25962 vp_p.n8412 vp_p.n8411 0.006
R25963 vp_p.n8415 vp_p.n8414 0.006
R25964 vp_p.n8426 vp_p.n8425 0.006
R25965 vp_p.n8429 vp_p.n8428 0.006
R25966 vp_p.n8440 vp_p.n8439 0.006
R25967 vp_p.n8443 vp_p.n8442 0.006
R25968 vp_p.n8454 vp_p.n8453 0.006
R25969 vp_p.n8457 vp_p.n8456 0.006
R25970 vp_p.n8468 vp_p.n8467 0.006
R25971 vp_p.n8471 vp_p.n8470 0.006
R25972 vp_p.n8482 vp_p.n8481 0.006
R25973 vp_p.n8485 vp_p.n8484 0.006
R25974 vp_p.n8496 vp_p.n8495 0.006
R25975 vp_p.n8499 vp_p.n8498 0.006
R25976 vp_p.n8510 vp_p.n8509 0.006
R25977 vp_p.n8513 vp_p.n8512 0.006
R25978 vp_p.n8524 vp_p.n8523 0.006
R25979 vp_p.n8527 vp_p.n8526 0.006
R25980 vp_p.n8538 vp_p.n8537 0.006
R25981 vp_p.n8541 vp_p.n8540 0.006
R25982 vp_p.n8552 vp_p.n8551 0.006
R25983 vp_p.n8555 vp_p.n8554 0.006
R25984 vp_p.n8566 vp_p.n8565 0.006
R25985 vp_p.n8569 vp_p.n8568 0.006
R25986 vp_p.n8580 vp_p.n8579 0.006
R25987 vp_p.n8583 vp_p.n8582 0.006
R25988 vp_p.n8594 vp_p.n8593 0.006
R25989 vp_p.n8597 vp_p.n8596 0.006
R25990 vp_p.n8608 vp_p.n8607 0.006
R25991 vp_p.n8611 vp_p.n8610 0.006
R25992 vp_p.n7579 vp_p.n7578 0.006
R25993 vp_p.n6163 vp_p.n6162 0.006
R25994 vp_p.n4740 vp_p.n4739 0.006
R25995 vp_p.n3316 vp_p.n3315 0.006
R25996 vp_p.n1891 vp_p.n1890 0.006
R25997 vp_p.n465 vp_p.n464 0.006
R25998 vp_p.n9211 vp_p.n9210 0.006
R25999 vp_p.n10648 vp_p.n10647 0.006
R26000 vp_p.n12086 vp_p.n12085 0.006
R26001 vp_p.n13850 vp_p.n13849 0.006
R26002 vp_p.n14889 vp_p.n14888 0.006
R26003 vp_p.n16317 vp_p.n16316 0.006
R26004 vp_p.n17744 vp_p.n17743 0.006
R26005 vp_p.n19170 vp_p.n19169 0.006
R26006 vp_p.n20595 vp_p.n20594 0.006
R26007 vp_p.n22019 vp_p.n22018 0.006
R26008 vp_p.n23442 vp_p.n23441 0.006
R26009 vp_p.n24864 vp_p.n24863 0.006
R26010 vp_p.n26285 vp_p.n26279 0.006
R26011 vp_p.n26289 vp_p.n26288 0.006
R26012 vp_p.n26299 vp_p.n26293 0.006
R26013 vp_p.n26303 vp_p.n26302 0.006
R26014 vp_p.n26313 vp_p.n26307 0.006
R26015 vp_p.n26317 vp_p.n26316 0.006
R26016 vp_p.n26327 vp_p.n26321 0.006
R26017 vp_p.n26331 vp_p.n26330 0.006
R26018 vp_p.n26341 vp_p.n26335 0.006
R26019 vp_p.n26345 vp_p.n26344 0.006
R26020 vp_p.n26355 vp_p.n26349 0.006
R26021 vp_p.n26359 vp_p.n26358 0.006
R26022 vp_p.n26369 vp_p.n26363 0.006
R26023 vp_p.n26373 vp_p.n26372 0.006
R26024 vp_p.n26383 vp_p.n26377 0.006
R26025 vp_p.n26387 vp_p.n26386 0.006
R26026 vp_p.n26397 vp_p.n26391 0.006
R26027 vp_p.n26401 vp_p.n26400 0.006
R26028 vp_p.n26411 vp_p.n26405 0.006
R26029 vp_p.n26415 vp_p.n26414 0.006
R26030 vp_p.n26425 vp_p.n26419 0.006
R26031 vp_p.n26429 vp_p.n26428 0.006
R26032 vp_p.n26439 vp_p.n26433 0.006
R26033 vp_p.n26443 vp_p.n26442 0.006
R26034 vp_p.n26453 vp_p.n26447 0.006
R26035 vp_p.n26457 vp_p.n26456 0.006
R26036 vp_p.n26467 vp_p.n26461 0.006
R26037 vp_p.n26471 vp_p.n26470 0.006
R26038 vp_p.n26481 vp_p.n26475 0.006
R26039 vp_p.n26485 vp_p.n26484 0.006
R26040 vp_p.n26495 vp_p.n26489 0.006
R26041 vp_p.n26499 vp_p.n26498 0.006
R26042 vp_p.n26509 vp_p.n26503 0.006
R26043 vp_p.n26513 vp_p.n26512 0.006
R26044 vp_p.n26523 vp_p.n26517 0.006
R26045 vp_p.n26527 vp_p.n26526 0.006
R26046 vp_p.n26537 vp_p.n26531 0.006
R26047 vp_p.n26541 vp_p.n26540 0.006
R26048 vp_p.n26551 vp_p.n26545 0.006
R26049 vp_p.n26555 vp_p.n26554 0.006
R26050 vp_p.n26565 vp_p.n26559 0.006
R26051 vp_p.n26569 vp_p.n26568 0.006
R26052 vp_p.n26579 vp_p.n26573 0.006
R26053 vp_p.n26583 vp_p.n26582 0.006
R26054 vp_p.n26593 vp_p.n26587 0.006
R26055 vp_p.n26597 vp_p.n26596 0.006
R26056 vp_p.n26607 vp_p.n26601 0.006
R26057 vp_p.n26611 vp_p.n26610 0.006
R26058 vp_p.n26621 vp_p.n26615 0.006
R26059 vp_p.n26625 vp_p.n26624 0.006
R26060 vp_p.n26635 vp_p.n26629 0.006
R26061 vp_p.n26639 vp_p.n26638 0.006
R26062 vp_p.n26649 vp_p.n26643 0.006
R26063 vp_p.n26653 vp_p.n26652 0.006
R26064 vp_p.n26663 vp_p.n26657 0.006
R26065 vp_p.n26667 vp_p.n26666 0.006
R26066 vp_p.n26677 vp_p.n26671 0.006
R26067 vp_p.n26681 vp_p.n26680 0.006
R26068 vp_p.n26691 vp_p.n26685 0.006
R26069 vp_p.n26695 vp_p.n26694 0.006
R26070 vp_p.n26705 vp_p.n26699 0.006
R26071 vp_p.n26709 vp_p.n26708 0.006
R26072 vp_p.n26719 vp_p.n26713 0.006
R26073 vp_p.n26723 vp_p.n26722 0.006
R26074 vp_p.n26733 vp_p.n26727 0.006
R26075 vp_p.n26737 vp_p.n26736 0.006
R26076 vp_p.n26747 vp_p.n26741 0.006
R26077 vp_p.n26751 vp_p.n26750 0.006
R26078 vp_p.n26761 vp_p.n26755 0.006
R26079 vp_p.n26765 vp_p.n26764 0.006
R26080 vp_p.n26775 vp_p.n26769 0.006
R26081 vp_p.n26779 vp_p.n26778 0.006
R26082 vp_p.n26789 vp_p.n26783 0.006
R26083 vp_p.n26793 vp_p.n26792 0.006
R26084 vp_p.n26803 vp_p.n26797 0.006
R26085 vp_p.n26807 vp_p.n26806 0.006
R26086 vp_p.n26817 vp_p.n26811 0.006
R26087 vp_p.n26821 vp_p.n26820 0.006
R26088 vp_p.n26831 vp_p.n26825 0.006
R26089 vp_p.n26835 vp_p.n26834 0.006
R26090 vp_p.n26845 vp_p.n26839 0.006
R26091 vp_p.n26849 vp_p.n26848 0.006
R26092 vp_p.n26859 vp_p.n26853 0.006
R26093 vp_p.n26863 vp_p.n26862 0.006
R26094 vp_p.n26873 vp_p.n26867 0.006
R26095 vp_p.n26877 vp_p.n26876 0.006
R26096 vp_p.n26887 vp_p.n26881 0.006
R26097 vp_p.n26891 vp_p.n26890 0.006
R26098 vp_p.n26901 vp_p.n26895 0.006
R26099 vp_p.n26905 vp_p.n26904 0.006
R26100 vp_p.n26915 vp_p.n26909 0.006
R26101 vp_p.n26919 vp_p.n26918 0.006
R26102 vp_p.n26929 vp_p.n26923 0.006
R26103 vp_p.n26933 vp_p.n26932 0.006
R26104 vp_p.n26943 vp_p.n26937 0.006
R26105 vp_p.n26947 vp_p.n26946 0.006
R26106 vp_p.n26957 vp_p.n26951 0.006
R26107 vp_p.n26961 vp_p.n26960 0.006
R26108 vp_p.n26971 vp_p.n26965 0.006
R26109 vp_p.n26975 vp_p.n26974 0.006
R26110 vp_p.n26985 vp_p.n26979 0.006
R26111 vp_p.n26989 vp_p.n26988 0.006
R26112 vp_p.n26999 vp_p.n26993 0.006
R26113 vp_p.n27003 vp_p.n27002 0.006
R26114 vp_p.n27013 vp_p.n27007 0.006
R26115 vp_p.n27017 vp_p.n27016 0.006
R26116 vp_p.n27027 vp_p.n27021 0.006
R26117 vp_p.n27031 vp_p.n27030 0.006
R26118 vp_p.n27041 vp_p.n27035 0.006
R26119 vp_p.n27045 vp_p.n27044 0.006
R26120 vp_p.n27055 vp_p.n27049 0.006
R26121 vp_p.n27059 vp_p.n27058 0.006
R26122 vp_p.n27069 vp_p.n27063 0.006
R26123 vp_p.n27073 vp_p.n27072 0.006
R26124 vp_p.n27083 vp_p.n27077 0.006
R26125 vp_p.n27087 vp_p.n27086 0.006
R26126 vp_p.n27097 vp_p.n27091 0.006
R26127 vp_p.n27101 vp_p.n27100 0.006
R26128 vp_p.n27111 vp_p.n27105 0.006
R26129 vp_p.n27115 vp_p.n27114 0.006
R26130 vp_p.n27125 vp_p.n27119 0.006
R26131 vp_p.n27129 vp_p.n27128 0.006
R26132 vp_p.n27139 vp_p.n27133 0.006
R26133 vp_p.n27143 vp_p.n27142 0.006
R26134 vp_p.n27153 vp_p.n27147 0.006
R26135 vp_p.n27157 vp_p.n27156 0.006
R26136 vp_p.n27167 vp_p.n27161 0.006
R26137 vp_p.n27171 vp_p.n27170 0.006
R26138 vp_p.n27181 vp_p.n27175 0.006
R26139 vp_p.n27185 vp_p.n27184 0.006
R26140 vp_p.n27195 vp_p.n27189 0.006
R26141 vp_p.n27199 vp_p.n27198 0.006
R26142 vp_p.n27209 vp_p.n27203 0.006
R26143 vp_p.n27213 vp_p.n27212 0.006
R26144 vp_p.n27223 vp_p.n27217 0.006
R26145 vp_p.n27227 vp_p.n27226 0.006
R26146 vp_p.n27237 vp_p.n27231 0.006
R26147 vp_p.n27241 vp_p.n27240 0.006
R26148 vp_p.n27251 vp_p.n27245 0.006
R26149 vp_p.n27255 vp_p.n27254 0.006
R26150 vp_p.n27265 vp_p.n27259 0.006
R26151 vp_p.n27269 vp_p.n27268 0.006
R26152 vp_p.n27279 vp_p.n27273 0.006
R26153 vp_p.n27283 vp_p.n27282 0.006
R26154 vp_p.n27293 vp_p.n27287 0.006
R26155 vp_p.n27297 vp_p.n27296 0.006
R26156 vp_p.n27307 vp_p.n27301 0.006
R26157 vp_p.n27311 vp_p.n27310 0.006
R26158 vp_p.n27321 vp_p.n27315 0.006
R26159 vp_p.n27325 vp_p.n27324 0.006
R26160 vp_p.n26290 vp_p.n26289 0.006
R26161 vp_p.n26293 vp_p.n26292 0.006
R26162 vp_p.n26304 vp_p.n26303 0.006
R26163 vp_p.n26307 vp_p.n26306 0.006
R26164 vp_p.n26318 vp_p.n26317 0.006
R26165 vp_p.n26321 vp_p.n26320 0.006
R26166 vp_p.n26332 vp_p.n26331 0.006
R26167 vp_p.n26335 vp_p.n26334 0.006
R26168 vp_p.n26346 vp_p.n26345 0.006
R26169 vp_p.n26349 vp_p.n26348 0.006
R26170 vp_p.n26360 vp_p.n26359 0.006
R26171 vp_p.n26363 vp_p.n26362 0.006
R26172 vp_p.n26374 vp_p.n26373 0.006
R26173 vp_p.n26377 vp_p.n26376 0.006
R26174 vp_p.n26388 vp_p.n26387 0.006
R26175 vp_p.n26391 vp_p.n26390 0.006
R26176 vp_p.n26402 vp_p.n26401 0.006
R26177 vp_p.n26405 vp_p.n26404 0.006
R26178 vp_p.n26416 vp_p.n26415 0.006
R26179 vp_p.n26419 vp_p.n26418 0.006
R26180 vp_p.n26430 vp_p.n26429 0.006
R26181 vp_p.n26433 vp_p.n26432 0.006
R26182 vp_p.n26444 vp_p.n26443 0.006
R26183 vp_p.n26447 vp_p.n26446 0.006
R26184 vp_p.n26458 vp_p.n26457 0.006
R26185 vp_p.n26461 vp_p.n26460 0.006
R26186 vp_p.n26472 vp_p.n26471 0.006
R26187 vp_p.n26475 vp_p.n26474 0.006
R26188 vp_p.n26486 vp_p.n26485 0.006
R26189 vp_p.n26489 vp_p.n26488 0.006
R26190 vp_p.n26500 vp_p.n26499 0.006
R26191 vp_p.n26503 vp_p.n26502 0.006
R26192 vp_p.n26514 vp_p.n26513 0.006
R26193 vp_p.n26517 vp_p.n26516 0.006
R26194 vp_p.n26528 vp_p.n26527 0.006
R26195 vp_p.n26531 vp_p.n26530 0.006
R26196 vp_p.n26542 vp_p.n26541 0.006
R26197 vp_p.n26545 vp_p.n26544 0.006
R26198 vp_p.n26556 vp_p.n26555 0.006
R26199 vp_p.n26559 vp_p.n26558 0.006
R26200 vp_p.n26570 vp_p.n26569 0.006
R26201 vp_p.n26573 vp_p.n26572 0.006
R26202 vp_p.n26584 vp_p.n26583 0.006
R26203 vp_p.n26587 vp_p.n26586 0.006
R26204 vp_p.n26598 vp_p.n26597 0.006
R26205 vp_p.n26601 vp_p.n26600 0.006
R26206 vp_p.n26612 vp_p.n26611 0.006
R26207 vp_p.n26615 vp_p.n26614 0.006
R26208 vp_p.n26626 vp_p.n26625 0.006
R26209 vp_p.n26629 vp_p.n26628 0.006
R26210 vp_p.n26640 vp_p.n26639 0.006
R26211 vp_p.n26643 vp_p.n26642 0.006
R26212 vp_p.n26654 vp_p.n26653 0.006
R26213 vp_p.n26657 vp_p.n26656 0.006
R26214 vp_p.n26668 vp_p.n26667 0.006
R26215 vp_p.n26671 vp_p.n26670 0.006
R26216 vp_p.n26682 vp_p.n26681 0.006
R26217 vp_p.n26685 vp_p.n26684 0.006
R26218 vp_p.n26696 vp_p.n26695 0.006
R26219 vp_p.n26699 vp_p.n26698 0.006
R26220 vp_p.n26710 vp_p.n26709 0.006
R26221 vp_p.n26713 vp_p.n26712 0.006
R26222 vp_p.n26724 vp_p.n26723 0.006
R26223 vp_p.n26727 vp_p.n26726 0.006
R26224 vp_p.n26738 vp_p.n26737 0.006
R26225 vp_p.n26741 vp_p.n26740 0.006
R26226 vp_p.n26752 vp_p.n26751 0.006
R26227 vp_p.n26755 vp_p.n26754 0.006
R26228 vp_p.n26766 vp_p.n26765 0.006
R26229 vp_p.n26769 vp_p.n26768 0.006
R26230 vp_p.n26780 vp_p.n26779 0.006
R26231 vp_p.n26783 vp_p.n26782 0.006
R26232 vp_p.n26794 vp_p.n26793 0.006
R26233 vp_p.n26797 vp_p.n26796 0.006
R26234 vp_p.n26808 vp_p.n26807 0.006
R26235 vp_p.n26811 vp_p.n26810 0.006
R26236 vp_p.n26822 vp_p.n26821 0.006
R26237 vp_p.n26825 vp_p.n26824 0.006
R26238 vp_p.n26836 vp_p.n26835 0.006
R26239 vp_p.n26839 vp_p.n26838 0.006
R26240 vp_p.n26850 vp_p.n26849 0.006
R26241 vp_p.n26853 vp_p.n26852 0.006
R26242 vp_p.n26864 vp_p.n26863 0.006
R26243 vp_p.n26867 vp_p.n26866 0.006
R26244 vp_p.n26878 vp_p.n26877 0.006
R26245 vp_p.n26881 vp_p.n26880 0.006
R26246 vp_p.n26892 vp_p.n26891 0.006
R26247 vp_p.n26895 vp_p.n26894 0.006
R26248 vp_p.n26906 vp_p.n26905 0.006
R26249 vp_p.n26909 vp_p.n26908 0.006
R26250 vp_p.n26920 vp_p.n26919 0.006
R26251 vp_p.n26923 vp_p.n26922 0.006
R26252 vp_p.n26934 vp_p.n26933 0.006
R26253 vp_p.n26937 vp_p.n26936 0.006
R26254 vp_p.n26948 vp_p.n26947 0.006
R26255 vp_p.n26951 vp_p.n26950 0.006
R26256 vp_p.n26962 vp_p.n26961 0.006
R26257 vp_p.n26965 vp_p.n26964 0.006
R26258 vp_p.n26976 vp_p.n26975 0.006
R26259 vp_p.n26979 vp_p.n26978 0.006
R26260 vp_p.n26990 vp_p.n26989 0.006
R26261 vp_p.n26993 vp_p.n26992 0.006
R26262 vp_p.n27004 vp_p.n27003 0.006
R26263 vp_p.n27007 vp_p.n27006 0.006
R26264 vp_p.n27018 vp_p.n27017 0.006
R26265 vp_p.n27021 vp_p.n27020 0.006
R26266 vp_p.n27032 vp_p.n27031 0.006
R26267 vp_p.n27035 vp_p.n27034 0.006
R26268 vp_p.n27046 vp_p.n27045 0.006
R26269 vp_p.n27049 vp_p.n27048 0.006
R26270 vp_p.n27060 vp_p.n27059 0.006
R26271 vp_p.n27063 vp_p.n27062 0.006
R26272 vp_p.n27074 vp_p.n27073 0.006
R26273 vp_p.n27077 vp_p.n27076 0.006
R26274 vp_p.n27088 vp_p.n27087 0.006
R26275 vp_p.n27091 vp_p.n27090 0.006
R26276 vp_p.n27102 vp_p.n27101 0.006
R26277 vp_p.n27105 vp_p.n27104 0.006
R26278 vp_p.n27116 vp_p.n27115 0.006
R26279 vp_p.n27119 vp_p.n27118 0.006
R26280 vp_p.n27130 vp_p.n27129 0.006
R26281 vp_p.n27133 vp_p.n27132 0.006
R26282 vp_p.n27144 vp_p.n27143 0.006
R26283 vp_p.n27147 vp_p.n27146 0.006
R26284 vp_p.n27158 vp_p.n27157 0.006
R26285 vp_p.n27161 vp_p.n27160 0.006
R26286 vp_p.n27172 vp_p.n27171 0.006
R26287 vp_p.n27175 vp_p.n27174 0.006
R26288 vp_p.n27186 vp_p.n27185 0.006
R26289 vp_p.n27189 vp_p.n27188 0.006
R26290 vp_p.n27200 vp_p.n27199 0.006
R26291 vp_p.n27203 vp_p.n27202 0.006
R26292 vp_p.n27214 vp_p.n27213 0.006
R26293 vp_p.n27217 vp_p.n27216 0.006
R26294 vp_p.n27228 vp_p.n27227 0.006
R26295 vp_p.n27231 vp_p.n27230 0.006
R26296 vp_p.n27242 vp_p.n27241 0.006
R26297 vp_p.n27245 vp_p.n27244 0.006
R26298 vp_p.n27256 vp_p.n27255 0.006
R26299 vp_p.n27259 vp_p.n27258 0.006
R26300 vp_p.n27270 vp_p.n27269 0.006
R26301 vp_p.n27273 vp_p.n27272 0.006
R26302 vp_p.n27284 vp_p.n27283 0.006
R26303 vp_p.n27287 vp_p.n27286 0.006
R26304 vp_p.n27298 vp_p.n27297 0.006
R26305 vp_p.n27301 vp_p.n27300 0.006
R26306 vp_p.n27312 vp_p.n27311 0.006
R26307 vp_p.n27315 vp_p.n27314 0.006
R26308 vp_p.n27326 vp_p.n27325 0.006
R26309 vp_p.n26279 vp_p.n26278 0.006
R26310 vp_p.n24859 vp_p.n24858 0.006
R26311 vp_p.n23437 vp_p.n23436 0.006
R26312 vp_p.n22014 vp_p.n22013 0.006
R26313 vp_p.n20590 vp_p.n20589 0.006
R26314 vp_p.n19165 vp_p.n19164 0.006
R26315 vp_p.n17739 vp_p.n17738 0.006
R26316 vp_p.n16312 vp_p.n16311 0.006
R26317 vp_p.n14884 vp_p.n14883 0.006
R26318 vp_p.n13845 vp_p.n13844 0.006
R26319 vp_p.n12081 vp_p.n12080 0.006
R26320 vp_p.n10643 vp_p.n10642 0.006
R26321 vp_p.n9206 vp_p.n9205 0.006
R26322 vp_p.n460 vp_p.n459 0.006
R26323 vp_p.n1886 vp_p.n1885 0.006
R26324 vp_p.n3311 vp_p.n3310 0.006
R26325 vp_p.n4735 vp_p.n4734 0.006
R26326 vp_p.n6158 vp_p.n6157 0.006
R26327 vp_p.n7575 vp_p.n7574 0.006
R26328 vp_p.n8621 vp_p.n8620 0.006
R26329 vp_p.n13007 vp_p.n13006 0.005
R26330 vp_p.n12993 vp_p.n12992 0.005
R26331 vp_p.n12979 vp_p.n12978 0.005
R26332 vp_p.n12965 vp_p.n12964 0.005
R26333 vp_p.n12951 vp_p.n12950 0.005
R26334 vp_p.n12937 vp_p.n12936 0.005
R26335 vp_p.n12923 vp_p.n12922 0.005
R26336 vp_p.n12909 vp_p.n12908 0.005
R26337 vp_p.n12895 vp_p.n12894 0.005
R26338 vp_p.n12881 vp_p.n12880 0.005
R26339 vp_p.n12867 vp_p.n12866 0.005
R26340 vp_p.n12853 vp_p.n12852 0.005
R26341 vp_p.n12839 vp_p.n12838 0.005
R26342 vp_p.n12825 vp_p.n12824 0.005
R26343 vp_p.n12811 vp_p.n12810 0.005
R26344 vp_p.n12797 vp_p.n12796 0.005
R26345 vp_p.n12783 vp_p.n12782 0.005
R26346 vp_p.n12769 vp_p.n12768 0.005
R26347 vp_p.n12755 vp_p.n12754 0.005
R26348 vp_p.n12741 vp_p.n12740 0.005
R26349 vp_p.n12727 vp_p.n12726 0.005
R26350 vp_p.n12713 vp_p.n12712 0.005
R26351 vp_p.n12699 vp_p.n12698 0.005
R26352 vp_p.n12685 vp_p.n12684 0.005
R26353 vp_p.n12671 vp_p.n12670 0.005
R26354 vp_p.n12657 vp_p.n12656 0.005
R26355 vp_p.n12643 vp_p.n12642 0.005
R26356 vp_p.n12629 vp_p.n12628 0.005
R26357 vp_p.n12615 vp_p.n12614 0.005
R26358 vp_p.n12601 vp_p.n12600 0.005
R26359 vp_p.n12587 vp_p.n12586 0.005
R26360 vp_p.n12573 vp_p.n12572 0.005
R26361 vp_p.n12559 vp_p.n12558 0.005
R26362 vp_p.n12545 vp_p.n12544 0.005
R26363 vp_p.n12531 vp_p.n12530 0.005
R26364 vp_p.n12517 vp_p.n12516 0.005
R26365 vp_p.n12503 vp_p.n12502 0.005
R26366 vp_p.n12489 vp_p.n12488 0.005
R26367 vp_p.n12475 vp_p.n12474 0.005
R26368 vp_p.n12461 vp_p.n12460 0.005
R26369 vp_p.n12447 vp_p.n12446 0.005
R26370 vp_p.n12433 vp_p.n12432 0.005
R26371 vp_p.n12419 vp_p.n12418 0.005
R26372 vp_p.n12405 vp_p.n12404 0.005
R26373 vp_p.n12391 vp_p.n12390 0.005
R26374 vp_p.n12377 vp_p.n12376 0.005
R26375 vp_p.n12363 vp_p.n12362 0.005
R26376 vp_p.n12349 vp_p.n12348 0.005
R26377 vp_p.n12335 vp_p.n12334 0.005
R26378 vp_p.n12321 vp_p.n12320 0.005
R26379 vp_p.n12307 vp_p.n12306 0.005
R26380 vp_p.n12293 vp_p.n12292 0.005
R26381 vp_p.n12279 vp_p.n12278 0.005
R26382 vp_p.n12265 vp_p.n12264 0.005
R26383 vp_p.n12251 vp_p.n12250 0.005
R26384 vp_p.n12237 vp_p.n12236 0.005
R26385 vp_p.n12223 vp_p.n12222 0.005
R26386 vp_p.n12209 vp_p.n12208 0.005
R26387 vp_p.n12195 vp_p.n12194 0.005
R26388 vp_p.n12181 vp_p.n12180 0.005
R26389 vp_p.n12167 vp_p.n12166 0.005
R26390 vp_p.n12153 vp_p.n12152 0.005
R26391 vp_p.n12139 vp_p.n12138 0.005
R26392 vp_p.n12125 vp_p.n12124 0.005
R26393 vp_p.n12111 vp_p.n12110 0.005
R26394 vp_p.n12097 vp_p.n12096 0.005
R26395 vp_p.n15810 vp_p.n15809 0.005
R26396 vp_p.n15796 vp_p.n15795 0.005
R26397 vp_p.n15782 vp_p.n15781 0.005
R26398 vp_p.n15768 vp_p.n15767 0.005
R26399 vp_p.n15754 vp_p.n15753 0.005
R26400 vp_p.n15740 vp_p.n15739 0.005
R26401 vp_p.n15726 vp_p.n15725 0.005
R26402 vp_p.n15712 vp_p.n15711 0.005
R26403 vp_p.n15698 vp_p.n15697 0.005
R26404 vp_p.n15684 vp_p.n15683 0.005
R26405 vp_p.n15670 vp_p.n15669 0.005
R26406 vp_p.n15656 vp_p.n15655 0.005
R26407 vp_p.n15642 vp_p.n15641 0.005
R26408 vp_p.n15628 vp_p.n15627 0.005
R26409 vp_p.n15614 vp_p.n15613 0.005
R26410 vp_p.n15600 vp_p.n15599 0.005
R26411 vp_p.n15586 vp_p.n15585 0.005
R26412 vp_p.n15572 vp_p.n15571 0.005
R26413 vp_p.n15558 vp_p.n15557 0.005
R26414 vp_p.n15544 vp_p.n15543 0.005
R26415 vp_p.n15530 vp_p.n15529 0.005
R26416 vp_p.n15516 vp_p.n15515 0.005
R26417 vp_p.n15502 vp_p.n15501 0.005
R26418 vp_p.n15488 vp_p.n15487 0.005
R26419 vp_p.n15474 vp_p.n15473 0.005
R26420 vp_p.n15460 vp_p.n15459 0.005
R26421 vp_p.n15446 vp_p.n15445 0.005
R26422 vp_p.n15432 vp_p.n15431 0.005
R26423 vp_p.n15418 vp_p.n15417 0.005
R26424 vp_p.n15404 vp_p.n15403 0.005
R26425 vp_p.n15390 vp_p.n15389 0.005
R26426 vp_p.n15376 vp_p.n15375 0.005
R26427 vp_p.n15362 vp_p.n15361 0.005
R26428 vp_p.n15348 vp_p.n15347 0.005
R26429 vp_p.n15334 vp_p.n15333 0.005
R26430 vp_p.n15320 vp_p.n15319 0.005
R26431 vp_p.n15306 vp_p.n15305 0.005
R26432 vp_p.n15292 vp_p.n15291 0.005
R26433 vp_p.n15278 vp_p.n15277 0.005
R26434 vp_p.n15264 vp_p.n15263 0.005
R26435 vp_p.n15250 vp_p.n15249 0.005
R26436 vp_p.n15236 vp_p.n15235 0.005
R26437 vp_p.n15222 vp_p.n15221 0.005
R26438 vp_p.n15208 vp_p.n15207 0.005
R26439 vp_p.n15194 vp_p.n15193 0.005
R26440 vp_p.n15180 vp_p.n15179 0.005
R26441 vp_p.n15166 vp_p.n15165 0.005
R26442 vp_p.n15152 vp_p.n15151 0.005
R26443 vp_p.n15138 vp_p.n15137 0.005
R26444 vp_p.n15124 vp_p.n15123 0.005
R26445 vp_p.n15110 vp_p.n15109 0.005
R26446 vp_p.n15096 vp_p.n15095 0.005
R26447 vp_p.n15082 vp_p.n15081 0.005
R26448 vp_p.n15068 vp_p.n15067 0.005
R26449 vp_p.n15054 vp_p.n15053 0.005
R26450 vp_p.n15040 vp_p.n15039 0.005
R26451 vp_p.n15026 vp_p.n15025 0.005
R26452 vp_p.n15012 vp_p.n15011 0.005
R26453 vp_p.n14998 vp_p.n14997 0.005
R26454 vp_p.n14984 vp_p.n14983 0.005
R26455 vp_p.n14970 vp_p.n14969 0.005
R26456 vp_p.n14956 vp_p.n14955 0.005
R26457 vp_p.n14942 vp_p.n14941 0.005
R26458 vp_p.n14928 vp_p.n14927 0.005
R26459 vp_p.n14914 vp_p.n14913 0.005
R26460 vp_p.n14900 vp_p.n14899 0.005
R26461 vp_p.n11583 vp_p.n11582 0.005
R26462 vp_p.n11569 vp_p.n11568 0.005
R26463 vp_p.n11555 vp_p.n11554 0.005
R26464 vp_p.n11541 vp_p.n11540 0.005
R26465 vp_p.n11527 vp_p.n11526 0.005
R26466 vp_p.n11513 vp_p.n11512 0.005
R26467 vp_p.n11499 vp_p.n11498 0.005
R26468 vp_p.n11485 vp_p.n11484 0.005
R26469 vp_p.n11471 vp_p.n11470 0.005
R26470 vp_p.n11457 vp_p.n11456 0.005
R26471 vp_p.n11443 vp_p.n11442 0.005
R26472 vp_p.n11429 vp_p.n11428 0.005
R26473 vp_p.n11415 vp_p.n11414 0.005
R26474 vp_p.n11401 vp_p.n11400 0.005
R26475 vp_p.n11387 vp_p.n11386 0.005
R26476 vp_p.n11373 vp_p.n11372 0.005
R26477 vp_p.n11359 vp_p.n11358 0.005
R26478 vp_p.n11345 vp_p.n11344 0.005
R26479 vp_p.n11331 vp_p.n11330 0.005
R26480 vp_p.n11317 vp_p.n11316 0.005
R26481 vp_p.n11303 vp_p.n11302 0.005
R26482 vp_p.n11289 vp_p.n11288 0.005
R26483 vp_p.n11275 vp_p.n11274 0.005
R26484 vp_p.n11261 vp_p.n11260 0.005
R26485 vp_p.n11247 vp_p.n11246 0.005
R26486 vp_p.n11233 vp_p.n11232 0.005
R26487 vp_p.n11219 vp_p.n11218 0.005
R26488 vp_p.n11205 vp_p.n11204 0.005
R26489 vp_p.n11191 vp_p.n11190 0.005
R26490 vp_p.n11177 vp_p.n11176 0.005
R26491 vp_p.n11163 vp_p.n11162 0.005
R26492 vp_p.n11149 vp_p.n11148 0.005
R26493 vp_p.n11135 vp_p.n11134 0.005
R26494 vp_p.n11121 vp_p.n11120 0.005
R26495 vp_p.n11107 vp_p.n11106 0.005
R26496 vp_p.n11093 vp_p.n11092 0.005
R26497 vp_p.n11079 vp_p.n11078 0.005
R26498 vp_p.n11065 vp_p.n11064 0.005
R26499 vp_p.n11051 vp_p.n11050 0.005
R26500 vp_p.n11037 vp_p.n11036 0.005
R26501 vp_p.n11023 vp_p.n11022 0.005
R26502 vp_p.n11009 vp_p.n11008 0.005
R26503 vp_p.n10995 vp_p.n10994 0.005
R26504 vp_p.n10981 vp_p.n10980 0.005
R26505 vp_p.n10967 vp_p.n10966 0.005
R26506 vp_p.n10953 vp_p.n10952 0.005
R26507 vp_p.n10939 vp_p.n10938 0.005
R26508 vp_p.n10925 vp_p.n10924 0.005
R26509 vp_p.n10911 vp_p.n10910 0.005
R26510 vp_p.n10897 vp_p.n10896 0.005
R26511 vp_p.n10883 vp_p.n10882 0.005
R26512 vp_p.n10869 vp_p.n10868 0.005
R26513 vp_p.n10855 vp_p.n10854 0.005
R26514 vp_p.n10841 vp_p.n10840 0.005
R26515 vp_p.n10827 vp_p.n10826 0.005
R26516 vp_p.n10813 vp_p.n10812 0.005
R26517 vp_p.n10799 vp_p.n10798 0.005
R26518 vp_p.n10785 vp_p.n10784 0.005
R26519 vp_p.n10771 vp_p.n10770 0.005
R26520 vp_p.n10757 vp_p.n10756 0.005
R26521 vp_p.n10743 vp_p.n10742 0.005
R26522 vp_p.n10729 vp_p.n10728 0.005
R26523 vp_p.n10715 vp_p.n10714 0.005
R26524 vp_p.n10701 vp_p.n10700 0.005
R26525 vp_p.n10687 vp_p.n10686 0.005
R26526 vp_p.n10673 vp_p.n10672 0.005
R26527 vp_p.n10659 vp_p.n10658 0.005
R26528 vp_p.n17252 vp_p.n17251 0.005
R26529 vp_p.n17238 vp_p.n17237 0.005
R26530 vp_p.n17224 vp_p.n17223 0.005
R26531 vp_p.n17210 vp_p.n17209 0.005
R26532 vp_p.n17196 vp_p.n17195 0.005
R26533 vp_p.n17182 vp_p.n17181 0.005
R26534 vp_p.n17168 vp_p.n17167 0.005
R26535 vp_p.n17154 vp_p.n17153 0.005
R26536 vp_p.n17140 vp_p.n17139 0.005
R26537 vp_p.n17126 vp_p.n17125 0.005
R26538 vp_p.n17112 vp_p.n17111 0.005
R26539 vp_p.n17098 vp_p.n17097 0.005
R26540 vp_p.n17084 vp_p.n17083 0.005
R26541 vp_p.n17070 vp_p.n17069 0.005
R26542 vp_p.n17056 vp_p.n17055 0.005
R26543 vp_p.n17042 vp_p.n17041 0.005
R26544 vp_p.n17028 vp_p.n17027 0.005
R26545 vp_p.n17014 vp_p.n17013 0.005
R26546 vp_p.n17000 vp_p.n16999 0.005
R26547 vp_p.n16986 vp_p.n16985 0.005
R26548 vp_p.n16972 vp_p.n16971 0.005
R26549 vp_p.n16958 vp_p.n16957 0.005
R26550 vp_p.n16944 vp_p.n16943 0.005
R26551 vp_p.n16930 vp_p.n16929 0.005
R26552 vp_p.n16916 vp_p.n16915 0.005
R26553 vp_p.n16902 vp_p.n16901 0.005
R26554 vp_p.n16888 vp_p.n16887 0.005
R26555 vp_p.n16874 vp_p.n16873 0.005
R26556 vp_p.n16860 vp_p.n16859 0.005
R26557 vp_p.n16846 vp_p.n16845 0.005
R26558 vp_p.n16832 vp_p.n16831 0.005
R26559 vp_p.n16818 vp_p.n16817 0.005
R26560 vp_p.n16804 vp_p.n16803 0.005
R26561 vp_p.n16790 vp_p.n16789 0.005
R26562 vp_p.n16776 vp_p.n16775 0.005
R26563 vp_p.n16762 vp_p.n16761 0.005
R26564 vp_p.n16748 vp_p.n16747 0.005
R26565 vp_p.n16734 vp_p.n16733 0.005
R26566 vp_p.n16720 vp_p.n16719 0.005
R26567 vp_p.n16706 vp_p.n16705 0.005
R26568 vp_p.n16692 vp_p.n16691 0.005
R26569 vp_p.n16678 vp_p.n16677 0.005
R26570 vp_p.n16664 vp_p.n16663 0.005
R26571 vp_p.n16650 vp_p.n16649 0.005
R26572 vp_p.n16636 vp_p.n16635 0.005
R26573 vp_p.n16622 vp_p.n16621 0.005
R26574 vp_p.n16608 vp_p.n16607 0.005
R26575 vp_p.n16594 vp_p.n16593 0.005
R26576 vp_p.n16580 vp_p.n16579 0.005
R26577 vp_p.n16566 vp_p.n16565 0.005
R26578 vp_p.n16552 vp_p.n16551 0.005
R26579 vp_p.n16538 vp_p.n16537 0.005
R26580 vp_p.n16524 vp_p.n16523 0.005
R26581 vp_p.n16510 vp_p.n16509 0.005
R26582 vp_p.n16496 vp_p.n16495 0.005
R26583 vp_p.n16482 vp_p.n16481 0.005
R26584 vp_p.n16468 vp_p.n16467 0.005
R26585 vp_p.n16454 vp_p.n16453 0.005
R26586 vp_p.n16440 vp_p.n16439 0.005
R26587 vp_p.n16426 vp_p.n16425 0.005
R26588 vp_p.n16412 vp_p.n16411 0.005
R26589 vp_p.n16398 vp_p.n16397 0.005
R26590 vp_p.n16384 vp_p.n16383 0.005
R26591 vp_p.n16370 vp_p.n16369 0.005
R26592 vp_p.n16356 vp_p.n16355 0.005
R26593 vp_p.n16342 vp_p.n16341 0.005
R26594 vp_p.n16328 vp_p.n16327 0.005
R26595 vp_p.n10160 vp_p.n10159 0.005
R26596 vp_p.n10146 vp_p.n10145 0.005
R26597 vp_p.n10132 vp_p.n10131 0.005
R26598 vp_p.n10118 vp_p.n10117 0.005
R26599 vp_p.n10104 vp_p.n10103 0.005
R26600 vp_p.n10090 vp_p.n10089 0.005
R26601 vp_p.n10076 vp_p.n10075 0.005
R26602 vp_p.n10062 vp_p.n10061 0.005
R26603 vp_p.n10048 vp_p.n10047 0.005
R26604 vp_p.n10034 vp_p.n10033 0.005
R26605 vp_p.n10020 vp_p.n10019 0.005
R26606 vp_p.n10006 vp_p.n10005 0.005
R26607 vp_p.n9992 vp_p.n9991 0.005
R26608 vp_p.n9978 vp_p.n9977 0.005
R26609 vp_p.n9964 vp_p.n9963 0.005
R26610 vp_p.n9950 vp_p.n9949 0.005
R26611 vp_p.n9936 vp_p.n9935 0.005
R26612 vp_p.n9922 vp_p.n9921 0.005
R26613 vp_p.n9908 vp_p.n9907 0.005
R26614 vp_p.n9894 vp_p.n9893 0.005
R26615 vp_p.n9880 vp_p.n9879 0.005
R26616 vp_p.n9866 vp_p.n9865 0.005
R26617 vp_p.n9852 vp_p.n9851 0.005
R26618 vp_p.n9838 vp_p.n9837 0.005
R26619 vp_p.n9824 vp_p.n9823 0.005
R26620 vp_p.n9810 vp_p.n9809 0.005
R26621 vp_p.n9796 vp_p.n9795 0.005
R26622 vp_p.n9782 vp_p.n9781 0.005
R26623 vp_p.n9768 vp_p.n9767 0.005
R26624 vp_p.n9754 vp_p.n9753 0.005
R26625 vp_p.n9740 vp_p.n9739 0.005
R26626 vp_p.n9726 vp_p.n9725 0.005
R26627 vp_p.n9712 vp_p.n9711 0.005
R26628 vp_p.n9698 vp_p.n9697 0.005
R26629 vp_p.n9684 vp_p.n9683 0.005
R26630 vp_p.n9670 vp_p.n9669 0.005
R26631 vp_p.n9656 vp_p.n9655 0.005
R26632 vp_p.n9642 vp_p.n9641 0.005
R26633 vp_p.n9628 vp_p.n9627 0.005
R26634 vp_p.n9614 vp_p.n9613 0.005
R26635 vp_p.n9600 vp_p.n9599 0.005
R26636 vp_p.n9586 vp_p.n9585 0.005
R26637 vp_p.n9572 vp_p.n9571 0.005
R26638 vp_p.n9558 vp_p.n9557 0.005
R26639 vp_p.n9544 vp_p.n9543 0.005
R26640 vp_p.n9530 vp_p.n9529 0.005
R26641 vp_p.n9516 vp_p.n9515 0.005
R26642 vp_p.n9502 vp_p.n9501 0.005
R26643 vp_p.n9488 vp_p.n9487 0.005
R26644 vp_p.n9474 vp_p.n9473 0.005
R26645 vp_p.n9460 vp_p.n9459 0.005
R26646 vp_p.n9446 vp_p.n9445 0.005
R26647 vp_p.n9432 vp_p.n9431 0.005
R26648 vp_p.n9418 vp_p.n9417 0.005
R26649 vp_p.n9404 vp_p.n9403 0.005
R26650 vp_p.n9390 vp_p.n9389 0.005
R26651 vp_p.n9376 vp_p.n9375 0.005
R26652 vp_p.n9362 vp_p.n9361 0.005
R26653 vp_p.n9348 vp_p.n9347 0.005
R26654 vp_p.n9334 vp_p.n9333 0.005
R26655 vp_p.n9320 vp_p.n9319 0.005
R26656 vp_p.n9306 vp_p.n9305 0.005
R26657 vp_p.n9292 vp_p.n9291 0.005
R26658 vp_p.n9278 vp_p.n9277 0.005
R26659 vp_p.n9264 vp_p.n9263 0.005
R26660 vp_p.n9250 vp_p.n9249 0.005
R26661 vp_p.n9236 vp_p.n9235 0.005
R26662 vp_p.n9222 vp_p.n9221 0.005
R26663 vp_p.n18693 vp_p.n18692 0.005
R26664 vp_p.n18679 vp_p.n18678 0.005
R26665 vp_p.n18665 vp_p.n18664 0.005
R26666 vp_p.n18651 vp_p.n18650 0.005
R26667 vp_p.n18637 vp_p.n18636 0.005
R26668 vp_p.n18623 vp_p.n18622 0.005
R26669 vp_p.n18609 vp_p.n18608 0.005
R26670 vp_p.n18595 vp_p.n18594 0.005
R26671 vp_p.n18581 vp_p.n18580 0.005
R26672 vp_p.n18567 vp_p.n18566 0.005
R26673 vp_p.n18553 vp_p.n18552 0.005
R26674 vp_p.n18539 vp_p.n18538 0.005
R26675 vp_p.n18525 vp_p.n18524 0.005
R26676 vp_p.n18511 vp_p.n18510 0.005
R26677 vp_p.n18497 vp_p.n18496 0.005
R26678 vp_p.n18483 vp_p.n18482 0.005
R26679 vp_p.n18469 vp_p.n18468 0.005
R26680 vp_p.n18455 vp_p.n18454 0.005
R26681 vp_p.n18441 vp_p.n18440 0.005
R26682 vp_p.n18427 vp_p.n18426 0.005
R26683 vp_p.n18413 vp_p.n18412 0.005
R26684 vp_p.n18399 vp_p.n18398 0.005
R26685 vp_p.n18385 vp_p.n18384 0.005
R26686 vp_p.n18371 vp_p.n18370 0.005
R26687 vp_p.n18357 vp_p.n18356 0.005
R26688 vp_p.n18343 vp_p.n18342 0.005
R26689 vp_p.n18329 vp_p.n18328 0.005
R26690 vp_p.n18315 vp_p.n18314 0.005
R26691 vp_p.n18301 vp_p.n18300 0.005
R26692 vp_p.n18287 vp_p.n18286 0.005
R26693 vp_p.n18273 vp_p.n18272 0.005
R26694 vp_p.n18259 vp_p.n18258 0.005
R26695 vp_p.n18245 vp_p.n18244 0.005
R26696 vp_p.n18231 vp_p.n18230 0.005
R26697 vp_p.n18217 vp_p.n18216 0.005
R26698 vp_p.n18203 vp_p.n18202 0.005
R26699 vp_p.n18189 vp_p.n18188 0.005
R26700 vp_p.n18175 vp_p.n18174 0.005
R26701 vp_p.n18161 vp_p.n18160 0.005
R26702 vp_p.n18147 vp_p.n18146 0.005
R26703 vp_p.n18133 vp_p.n18132 0.005
R26704 vp_p.n18119 vp_p.n18118 0.005
R26705 vp_p.n18105 vp_p.n18104 0.005
R26706 vp_p.n18091 vp_p.n18090 0.005
R26707 vp_p.n18077 vp_p.n18076 0.005
R26708 vp_p.n18063 vp_p.n18062 0.005
R26709 vp_p.n18049 vp_p.n18048 0.005
R26710 vp_p.n18035 vp_p.n18034 0.005
R26711 vp_p.n18021 vp_p.n18020 0.005
R26712 vp_p.n18007 vp_p.n18006 0.005
R26713 vp_p.n17993 vp_p.n17992 0.005
R26714 vp_p.n17979 vp_p.n17978 0.005
R26715 vp_p.n17965 vp_p.n17964 0.005
R26716 vp_p.n17951 vp_p.n17950 0.005
R26717 vp_p.n17937 vp_p.n17936 0.005
R26718 vp_p.n17923 vp_p.n17922 0.005
R26719 vp_p.n17909 vp_p.n17908 0.005
R26720 vp_p.n17895 vp_p.n17894 0.005
R26721 vp_p.n17881 vp_p.n17880 0.005
R26722 vp_p.n17867 vp_p.n17866 0.005
R26723 vp_p.n17853 vp_p.n17852 0.005
R26724 vp_p.n17839 vp_p.n17838 0.005
R26725 vp_p.n17825 vp_p.n17824 0.005
R26726 vp_p.n17811 vp_p.n17810 0.005
R26727 vp_p.n17797 vp_p.n17796 0.005
R26728 vp_p.n17783 vp_p.n17782 0.005
R26729 vp_p.n17769 vp_p.n17768 0.005
R26730 vp_p.n17755 vp_p.n17754 0.005
R26731 vp_p.n1428 vp_p.n1427 0.005
R26732 vp_p.n1414 vp_p.n1413 0.005
R26733 vp_p.n1400 vp_p.n1399 0.005
R26734 vp_p.n1386 vp_p.n1385 0.005
R26735 vp_p.n1372 vp_p.n1371 0.005
R26736 vp_p.n1358 vp_p.n1357 0.005
R26737 vp_p.n1344 vp_p.n1343 0.005
R26738 vp_p.n1330 vp_p.n1329 0.005
R26739 vp_p.n1316 vp_p.n1315 0.005
R26740 vp_p.n1302 vp_p.n1301 0.005
R26741 vp_p.n1288 vp_p.n1287 0.005
R26742 vp_p.n1274 vp_p.n1273 0.005
R26743 vp_p.n1260 vp_p.n1259 0.005
R26744 vp_p.n1246 vp_p.n1245 0.005
R26745 vp_p.n1232 vp_p.n1231 0.005
R26746 vp_p.n1218 vp_p.n1217 0.005
R26747 vp_p.n1204 vp_p.n1203 0.005
R26748 vp_p.n1190 vp_p.n1189 0.005
R26749 vp_p.n1176 vp_p.n1175 0.005
R26750 vp_p.n1162 vp_p.n1161 0.005
R26751 vp_p.n1148 vp_p.n1147 0.005
R26752 vp_p.n1134 vp_p.n1133 0.005
R26753 vp_p.n1120 vp_p.n1119 0.005
R26754 vp_p.n1106 vp_p.n1105 0.005
R26755 vp_p.n1092 vp_p.n1091 0.005
R26756 vp_p.n1078 vp_p.n1077 0.005
R26757 vp_p.n1064 vp_p.n1063 0.005
R26758 vp_p.n1050 vp_p.n1049 0.005
R26759 vp_p.n1036 vp_p.n1035 0.005
R26760 vp_p.n1022 vp_p.n1021 0.005
R26761 vp_p.n1008 vp_p.n1007 0.005
R26762 vp_p.n994 vp_p.n993 0.005
R26763 vp_p.n980 vp_p.n979 0.005
R26764 vp_p.n966 vp_p.n965 0.005
R26765 vp_p.n952 vp_p.n951 0.005
R26766 vp_p.n938 vp_p.n937 0.005
R26767 vp_p.n924 vp_p.n923 0.005
R26768 vp_p.n910 vp_p.n909 0.005
R26769 vp_p.n896 vp_p.n895 0.005
R26770 vp_p.n882 vp_p.n881 0.005
R26771 vp_p.n868 vp_p.n867 0.005
R26772 vp_p.n854 vp_p.n853 0.005
R26773 vp_p.n840 vp_p.n839 0.005
R26774 vp_p.n826 vp_p.n825 0.005
R26775 vp_p.n812 vp_p.n811 0.005
R26776 vp_p.n798 vp_p.n797 0.005
R26777 vp_p.n784 vp_p.n783 0.005
R26778 vp_p.n770 vp_p.n769 0.005
R26779 vp_p.n756 vp_p.n755 0.005
R26780 vp_p.n742 vp_p.n741 0.005
R26781 vp_p.n728 vp_p.n727 0.005
R26782 vp_p.n714 vp_p.n713 0.005
R26783 vp_p.n700 vp_p.n699 0.005
R26784 vp_p.n686 vp_p.n685 0.005
R26785 vp_p.n672 vp_p.n671 0.005
R26786 vp_p.n658 vp_p.n657 0.005
R26787 vp_p.n644 vp_p.n643 0.005
R26788 vp_p.n630 vp_p.n629 0.005
R26789 vp_p.n616 vp_p.n615 0.005
R26790 vp_p.n602 vp_p.n601 0.005
R26791 vp_p.n588 vp_p.n587 0.005
R26792 vp_p.n574 vp_p.n573 0.005
R26793 vp_p.n560 vp_p.n559 0.005
R26794 vp_p.n546 vp_p.n545 0.005
R26795 vp_p.n532 vp_p.n531 0.005
R26796 vp_p.n518 vp_p.n517 0.005
R26797 vp_p.n504 vp_p.n503 0.005
R26798 vp_p.n490 vp_p.n489 0.005
R26799 vp_p.n476 vp_p.n475 0.005
R26800 vp_p.n20133 vp_p.n20132 0.005
R26801 vp_p.n20119 vp_p.n20118 0.005
R26802 vp_p.n20105 vp_p.n20104 0.005
R26803 vp_p.n20091 vp_p.n20090 0.005
R26804 vp_p.n20077 vp_p.n20076 0.005
R26805 vp_p.n20063 vp_p.n20062 0.005
R26806 vp_p.n20049 vp_p.n20048 0.005
R26807 vp_p.n20035 vp_p.n20034 0.005
R26808 vp_p.n20021 vp_p.n20020 0.005
R26809 vp_p.n20007 vp_p.n20006 0.005
R26810 vp_p.n19993 vp_p.n19992 0.005
R26811 vp_p.n19979 vp_p.n19978 0.005
R26812 vp_p.n19965 vp_p.n19964 0.005
R26813 vp_p.n19951 vp_p.n19950 0.005
R26814 vp_p.n19937 vp_p.n19936 0.005
R26815 vp_p.n19923 vp_p.n19922 0.005
R26816 vp_p.n19909 vp_p.n19908 0.005
R26817 vp_p.n19895 vp_p.n19894 0.005
R26818 vp_p.n19881 vp_p.n19880 0.005
R26819 vp_p.n19867 vp_p.n19866 0.005
R26820 vp_p.n19853 vp_p.n19852 0.005
R26821 vp_p.n19839 vp_p.n19838 0.005
R26822 vp_p.n19825 vp_p.n19824 0.005
R26823 vp_p.n19811 vp_p.n19810 0.005
R26824 vp_p.n19797 vp_p.n19796 0.005
R26825 vp_p.n19783 vp_p.n19782 0.005
R26826 vp_p.n19769 vp_p.n19768 0.005
R26827 vp_p.n19755 vp_p.n19754 0.005
R26828 vp_p.n19741 vp_p.n19740 0.005
R26829 vp_p.n19727 vp_p.n19726 0.005
R26830 vp_p.n19713 vp_p.n19712 0.005
R26831 vp_p.n19699 vp_p.n19698 0.005
R26832 vp_p.n19685 vp_p.n19684 0.005
R26833 vp_p.n19671 vp_p.n19670 0.005
R26834 vp_p.n19657 vp_p.n19656 0.005
R26835 vp_p.n19643 vp_p.n19642 0.005
R26836 vp_p.n19629 vp_p.n19628 0.005
R26837 vp_p.n19615 vp_p.n19614 0.005
R26838 vp_p.n19601 vp_p.n19600 0.005
R26839 vp_p.n19587 vp_p.n19586 0.005
R26840 vp_p.n19573 vp_p.n19572 0.005
R26841 vp_p.n19559 vp_p.n19558 0.005
R26842 vp_p.n19545 vp_p.n19544 0.005
R26843 vp_p.n19531 vp_p.n19530 0.005
R26844 vp_p.n19517 vp_p.n19516 0.005
R26845 vp_p.n19503 vp_p.n19502 0.005
R26846 vp_p.n19489 vp_p.n19488 0.005
R26847 vp_p.n19475 vp_p.n19474 0.005
R26848 vp_p.n19461 vp_p.n19460 0.005
R26849 vp_p.n19447 vp_p.n19446 0.005
R26850 vp_p.n19433 vp_p.n19432 0.005
R26851 vp_p.n19419 vp_p.n19418 0.005
R26852 vp_p.n19405 vp_p.n19404 0.005
R26853 vp_p.n19391 vp_p.n19390 0.005
R26854 vp_p.n19377 vp_p.n19376 0.005
R26855 vp_p.n19363 vp_p.n19362 0.005
R26856 vp_p.n19349 vp_p.n19348 0.005
R26857 vp_p.n19335 vp_p.n19334 0.005
R26858 vp_p.n19321 vp_p.n19320 0.005
R26859 vp_p.n19307 vp_p.n19306 0.005
R26860 vp_p.n19293 vp_p.n19292 0.005
R26861 vp_p.n19279 vp_p.n19278 0.005
R26862 vp_p.n19265 vp_p.n19264 0.005
R26863 vp_p.n19251 vp_p.n19250 0.005
R26864 vp_p.n19237 vp_p.n19236 0.005
R26865 vp_p.n19223 vp_p.n19222 0.005
R26866 vp_p.n19209 vp_p.n19208 0.005
R26867 vp_p.n19195 vp_p.n19194 0.005
R26868 vp_p.n19181 vp_p.n19180 0.005
R26869 vp_p.n2868 vp_p.n2867 0.005
R26870 vp_p.n2854 vp_p.n2853 0.005
R26871 vp_p.n2840 vp_p.n2839 0.005
R26872 vp_p.n2826 vp_p.n2825 0.005
R26873 vp_p.n2812 vp_p.n2811 0.005
R26874 vp_p.n2798 vp_p.n2797 0.005
R26875 vp_p.n2784 vp_p.n2783 0.005
R26876 vp_p.n2770 vp_p.n2769 0.005
R26877 vp_p.n2756 vp_p.n2755 0.005
R26878 vp_p.n2742 vp_p.n2741 0.005
R26879 vp_p.n2728 vp_p.n2727 0.005
R26880 vp_p.n2714 vp_p.n2713 0.005
R26881 vp_p.n2700 vp_p.n2699 0.005
R26882 vp_p.n2686 vp_p.n2685 0.005
R26883 vp_p.n2672 vp_p.n2671 0.005
R26884 vp_p.n2658 vp_p.n2657 0.005
R26885 vp_p.n2644 vp_p.n2643 0.005
R26886 vp_p.n2630 vp_p.n2629 0.005
R26887 vp_p.n2616 vp_p.n2615 0.005
R26888 vp_p.n2602 vp_p.n2601 0.005
R26889 vp_p.n2588 vp_p.n2587 0.005
R26890 vp_p.n2574 vp_p.n2573 0.005
R26891 vp_p.n2560 vp_p.n2559 0.005
R26892 vp_p.n2546 vp_p.n2545 0.005
R26893 vp_p.n2532 vp_p.n2531 0.005
R26894 vp_p.n2518 vp_p.n2517 0.005
R26895 vp_p.n2504 vp_p.n2503 0.005
R26896 vp_p.n2490 vp_p.n2489 0.005
R26897 vp_p.n2476 vp_p.n2475 0.005
R26898 vp_p.n2462 vp_p.n2461 0.005
R26899 vp_p.n2448 vp_p.n2447 0.005
R26900 vp_p.n2434 vp_p.n2433 0.005
R26901 vp_p.n2420 vp_p.n2419 0.005
R26902 vp_p.n2406 vp_p.n2405 0.005
R26903 vp_p.n2392 vp_p.n2391 0.005
R26904 vp_p.n2378 vp_p.n2377 0.005
R26905 vp_p.n2364 vp_p.n2363 0.005
R26906 vp_p.n2350 vp_p.n2349 0.005
R26907 vp_p.n2336 vp_p.n2335 0.005
R26908 vp_p.n2322 vp_p.n2321 0.005
R26909 vp_p.n2308 vp_p.n2307 0.005
R26910 vp_p.n2294 vp_p.n2293 0.005
R26911 vp_p.n2280 vp_p.n2279 0.005
R26912 vp_p.n2266 vp_p.n2265 0.005
R26913 vp_p.n2252 vp_p.n2251 0.005
R26914 vp_p.n2238 vp_p.n2237 0.005
R26915 vp_p.n2224 vp_p.n2223 0.005
R26916 vp_p.n2210 vp_p.n2209 0.005
R26917 vp_p.n2196 vp_p.n2195 0.005
R26918 vp_p.n2182 vp_p.n2181 0.005
R26919 vp_p.n2168 vp_p.n2167 0.005
R26920 vp_p.n2154 vp_p.n2153 0.005
R26921 vp_p.n2140 vp_p.n2139 0.005
R26922 vp_p.n2126 vp_p.n2125 0.005
R26923 vp_p.n2112 vp_p.n2111 0.005
R26924 vp_p.n2098 vp_p.n2097 0.005
R26925 vp_p.n2084 vp_p.n2083 0.005
R26926 vp_p.n2070 vp_p.n2069 0.005
R26927 vp_p.n2056 vp_p.n2055 0.005
R26928 vp_p.n2042 vp_p.n2041 0.005
R26929 vp_p.n2028 vp_p.n2027 0.005
R26930 vp_p.n2014 vp_p.n2013 0.005
R26931 vp_p.n2000 vp_p.n1999 0.005
R26932 vp_p.n1986 vp_p.n1985 0.005
R26933 vp_p.n1972 vp_p.n1971 0.005
R26934 vp_p.n1958 vp_p.n1957 0.005
R26935 vp_p.n1944 vp_p.n1943 0.005
R26936 vp_p.n1930 vp_p.n1929 0.005
R26937 vp_p.n1916 vp_p.n1915 0.005
R26938 vp_p.n1902 vp_p.n1901 0.005
R26939 vp_p.n21572 vp_p.n21571 0.005
R26940 vp_p.n21558 vp_p.n21557 0.005
R26941 vp_p.n21544 vp_p.n21543 0.005
R26942 vp_p.n21530 vp_p.n21529 0.005
R26943 vp_p.n21516 vp_p.n21515 0.005
R26944 vp_p.n21502 vp_p.n21501 0.005
R26945 vp_p.n21488 vp_p.n21487 0.005
R26946 vp_p.n21474 vp_p.n21473 0.005
R26947 vp_p.n21460 vp_p.n21459 0.005
R26948 vp_p.n21446 vp_p.n21445 0.005
R26949 vp_p.n21432 vp_p.n21431 0.005
R26950 vp_p.n21418 vp_p.n21417 0.005
R26951 vp_p.n21404 vp_p.n21403 0.005
R26952 vp_p.n21390 vp_p.n21389 0.005
R26953 vp_p.n21376 vp_p.n21375 0.005
R26954 vp_p.n21362 vp_p.n21361 0.005
R26955 vp_p.n21348 vp_p.n21347 0.005
R26956 vp_p.n21334 vp_p.n21333 0.005
R26957 vp_p.n21320 vp_p.n21319 0.005
R26958 vp_p.n21306 vp_p.n21305 0.005
R26959 vp_p.n21292 vp_p.n21291 0.005
R26960 vp_p.n21278 vp_p.n21277 0.005
R26961 vp_p.n21264 vp_p.n21263 0.005
R26962 vp_p.n21250 vp_p.n21249 0.005
R26963 vp_p.n21236 vp_p.n21235 0.005
R26964 vp_p.n21222 vp_p.n21221 0.005
R26965 vp_p.n21208 vp_p.n21207 0.005
R26966 vp_p.n21194 vp_p.n21193 0.005
R26967 vp_p.n21180 vp_p.n21179 0.005
R26968 vp_p.n21166 vp_p.n21165 0.005
R26969 vp_p.n21152 vp_p.n21151 0.005
R26970 vp_p.n21138 vp_p.n21137 0.005
R26971 vp_p.n21124 vp_p.n21123 0.005
R26972 vp_p.n21110 vp_p.n21109 0.005
R26973 vp_p.n21096 vp_p.n21095 0.005
R26974 vp_p.n21082 vp_p.n21081 0.005
R26975 vp_p.n21068 vp_p.n21067 0.005
R26976 vp_p.n21054 vp_p.n21053 0.005
R26977 vp_p.n21040 vp_p.n21039 0.005
R26978 vp_p.n21026 vp_p.n21025 0.005
R26979 vp_p.n21012 vp_p.n21011 0.005
R26980 vp_p.n20998 vp_p.n20997 0.005
R26981 vp_p.n20984 vp_p.n20983 0.005
R26982 vp_p.n20970 vp_p.n20969 0.005
R26983 vp_p.n20956 vp_p.n20955 0.005
R26984 vp_p.n20942 vp_p.n20941 0.005
R26985 vp_p.n20928 vp_p.n20927 0.005
R26986 vp_p.n20914 vp_p.n20913 0.005
R26987 vp_p.n20900 vp_p.n20899 0.005
R26988 vp_p.n20886 vp_p.n20885 0.005
R26989 vp_p.n20872 vp_p.n20871 0.005
R26990 vp_p.n20858 vp_p.n20857 0.005
R26991 vp_p.n20844 vp_p.n20843 0.005
R26992 vp_p.n20830 vp_p.n20829 0.005
R26993 vp_p.n20816 vp_p.n20815 0.005
R26994 vp_p.n20802 vp_p.n20801 0.005
R26995 vp_p.n20788 vp_p.n20787 0.005
R26996 vp_p.n20774 vp_p.n20773 0.005
R26997 vp_p.n20760 vp_p.n20759 0.005
R26998 vp_p.n20746 vp_p.n20745 0.005
R26999 vp_p.n20732 vp_p.n20731 0.005
R27000 vp_p.n20718 vp_p.n20717 0.005
R27001 vp_p.n20704 vp_p.n20703 0.005
R27002 vp_p.n20690 vp_p.n20689 0.005
R27003 vp_p.n20676 vp_p.n20675 0.005
R27004 vp_p.n20662 vp_p.n20661 0.005
R27005 vp_p.n20648 vp_p.n20647 0.005
R27006 vp_p.n20634 vp_p.n20633 0.005
R27007 vp_p.n20620 vp_p.n20619 0.005
R27008 vp_p.n20606 vp_p.n20605 0.005
R27009 vp_p.n4307 vp_p.n4306 0.005
R27010 vp_p.n4293 vp_p.n4292 0.005
R27011 vp_p.n4279 vp_p.n4278 0.005
R27012 vp_p.n4265 vp_p.n4264 0.005
R27013 vp_p.n4251 vp_p.n4250 0.005
R27014 vp_p.n4237 vp_p.n4236 0.005
R27015 vp_p.n4223 vp_p.n4222 0.005
R27016 vp_p.n4209 vp_p.n4208 0.005
R27017 vp_p.n4195 vp_p.n4194 0.005
R27018 vp_p.n4181 vp_p.n4180 0.005
R27019 vp_p.n4167 vp_p.n4166 0.005
R27020 vp_p.n4153 vp_p.n4152 0.005
R27021 vp_p.n4139 vp_p.n4138 0.005
R27022 vp_p.n4125 vp_p.n4124 0.005
R27023 vp_p.n4111 vp_p.n4110 0.005
R27024 vp_p.n4097 vp_p.n4096 0.005
R27025 vp_p.n4083 vp_p.n4082 0.005
R27026 vp_p.n4069 vp_p.n4068 0.005
R27027 vp_p.n4055 vp_p.n4054 0.005
R27028 vp_p.n4041 vp_p.n4040 0.005
R27029 vp_p.n4027 vp_p.n4026 0.005
R27030 vp_p.n4013 vp_p.n4012 0.005
R27031 vp_p.n3999 vp_p.n3998 0.005
R27032 vp_p.n3985 vp_p.n3984 0.005
R27033 vp_p.n3971 vp_p.n3970 0.005
R27034 vp_p.n3957 vp_p.n3956 0.005
R27035 vp_p.n3943 vp_p.n3942 0.005
R27036 vp_p.n3929 vp_p.n3928 0.005
R27037 vp_p.n3915 vp_p.n3914 0.005
R27038 vp_p.n3901 vp_p.n3900 0.005
R27039 vp_p.n3887 vp_p.n3886 0.005
R27040 vp_p.n3873 vp_p.n3872 0.005
R27041 vp_p.n3859 vp_p.n3858 0.005
R27042 vp_p.n3845 vp_p.n3844 0.005
R27043 vp_p.n3831 vp_p.n3830 0.005
R27044 vp_p.n3817 vp_p.n3816 0.005
R27045 vp_p.n3803 vp_p.n3802 0.005
R27046 vp_p.n3789 vp_p.n3788 0.005
R27047 vp_p.n3775 vp_p.n3774 0.005
R27048 vp_p.n3761 vp_p.n3760 0.005
R27049 vp_p.n3747 vp_p.n3746 0.005
R27050 vp_p.n3733 vp_p.n3732 0.005
R27051 vp_p.n3719 vp_p.n3718 0.005
R27052 vp_p.n3705 vp_p.n3704 0.005
R27053 vp_p.n3691 vp_p.n3690 0.005
R27054 vp_p.n3677 vp_p.n3676 0.005
R27055 vp_p.n3663 vp_p.n3662 0.005
R27056 vp_p.n3649 vp_p.n3648 0.005
R27057 vp_p.n3635 vp_p.n3634 0.005
R27058 vp_p.n3621 vp_p.n3620 0.005
R27059 vp_p.n3607 vp_p.n3606 0.005
R27060 vp_p.n3593 vp_p.n3592 0.005
R27061 vp_p.n3579 vp_p.n3578 0.005
R27062 vp_p.n3565 vp_p.n3564 0.005
R27063 vp_p.n3551 vp_p.n3550 0.005
R27064 vp_p.n3537 vp_p.n3536 0.005
R27065 vp_p.n3523 vp_p.n3522 0.005
R27066 vp_p.n3509 vp_p.n3508 0.005
R27067 vp_p.n3495 vp_p.n3494 0.005
R27068 vp_p.n3481 vp_p.n3480 0.005
R27069 vp_p.n3467 vp_p.n3466 0.005
R27070 vp_p.n3453 vp_p.n3452 0.005
R27071 vp_p.n3439 vp_p.n3438 0.005
R27072 vp_p.n3425 vp_p.n3424 0.005
R27073 vp_p.n3411 vp_p.n3410 0.005
R27074 vp_p.n3397 vp_p.n3396 0.005
R27075 vp_p.n3383 vp_p.n3382 0.005
R27076 vp_p.n3369 vp_p.n3368 0.005
R27077 vp_p.n3355 vp_p.n3354 0.005
R27078 vp_p.n3341 vp_p.n3340 0.005
R27079 vp_p.n3327 vp_p.n3326 0.005
R27080 vp_p.n23010 vp_p.n23009 0.005
R27081 vp_p.n22996 vp_p.n22995 0.005
R27082 vp_p.n22982 vp_p.n22981 0.005
R27083 vp_p.n22968 vp_p.n22967 0.005
R27084 vp_p.n22954 vp_p.n22953 0.005
R27085 vp_p.n22940 vp_p.n22939 0.005
R27086 vp_p.n22926 vp_p.n22925 0.005
R27087 vp_p.n22912 vp_p.n22911 0.005
R27088 vp_p.n22898 vp_p.n22897 0.005
R27089 vp_p.n22884 vp_p.n22883 0.005
R27090 vp_p.n22870 vp_p.n22869 0.005
R27091 vp_p.n22856 vp_p.n22855 0.005
R27092 vp_p.n22842 vp_p.n22841 0.005
R27093 vp_p.n22828 vp_p.n22827 0.005
R27094 vp_p.n22814 vp_p.n22813 0.005
R27095 vp_p.n22800 vp_p.n22799 0.005
R27096 vp_p.n22786 vp_p.n22785 0.005
R27097 vp_p.n22772 vp_p.n22771 0.005
R27098 vp_p.n22758 vp_p.n22757 0.005
R27099 vp_p.n22744 vp_p.n22743 0.005
R27100 vp_p.n22730 vp_p.n22729 0.005
R27101 vp_p.n22716 vp_p.n22715 0.005
R27102 vp_p.n22702 vp_p.n22701 0.005
R27103 vp_p.n22688 vp_p.n22687 0.005
R27104 vp_p.n22674 vp_p.n22673 0.005
R27105 vp_p.n22660 vp_p.n22659 0.005
R27106 vp_p.n22646 vp_p.n22645 0.005
R27107 vp_p.n22632 vp_p.n22631 0.005
R27108 vp_p.n22618 vp_p.n22617 0.005
R27109 vp_p.n22604 vp_p.n22603 0.005
R27110 vp_p.n22590 vp_p.n22589 0.005
R27111 vp_p.n22576 vp_p.n22575 0.005
R27112 vp_p.n22562 vp_p.n22561 0.005
R27113 vp_p.n22548 vp_p.n22547 0.005
R27114 vp_p.n22534 vp_p.n22533 0.005
R27115 vp_p.n22520 vp_p.n22519 0.005
R27116 vp_p.n22506 vp_p.n22505 0.005
R27117 vp_p.n22492 vp_p.n22491 0.005
R27118 vp_p.n22478 vp_p.n22477 0.005
R27119 vp_p.n22464 vp_p.n22463 0.005
R27120 vp_p.n22450 vp_p.n22449 0.005
R27121 vp_p.n22436 vp_p.n22435 0.005
R27122 vp_p.n22422 vp_p.n22421 0.005
R27123 vp_p.n22408 vp_p.n22407 0.005
R27124 vp_p.n22394 vp_p.n22393 0.005
R27125 vp_p.n22380 vp_p.n22379 0.005
R27126 vp_p.n22366 vp_p.n22365 0.005
R27127 vp_p.n22352 vp_p.n22351 0.005
R27128 vp_p.n22338 vp_p.n22337 0.005
R27129 vp_p.n22324 vp_p.n22323 0.005
R27130 vp_p.n22310 vp_p.n22309 0.005
R27131 vp_p.n22296 vp_p.n22295 0.005
R27132 vp_p.n22282 vp_p.n22281 0.005
R27133 vp_p.n22268 vp_p.n22267 0.005
R27134 vp_p.n22254 vp_p.n22253 0.005
R27135 vp_p.n22240 vp_p.n22239 0.005
R27136 vp_p.n22226 vp_p.n22225 0.005
R27137 vp_p.n22212 vp_p.n22211 0.005
R27138 vp_p.n22198 vp_p.n22197 0.005
R27139 vp_p.n22184 vp_p.n22183 0.005
R27140 vp_p.n22170 vp_p.n22169 0.005
R27141 vp_p.n22156 vp_p.n22155 0.005
R27142 vp_p.n22142 vp_p.n22141 0.005
R27143 vp_p.n22128 vp_p.n22127 0.005
R27144 vp_p.n22114 vp_p.n22113 0.005
R27145 vp_p.n22100 vp_p.n22099 0.005
R27146 vp_p.n22086 vp_p.n22085 0.005
R27147 vp_p.n22072 vp_p.n22071 0.005
R27148 vp_p.n22058 vp_p.n22057 0.005
R27149 vp_p.n22044 vp_p.n22043 0.005
R27150 vp_p.n22030 vp_p.n22029 0.005
R27151 vp_p.n5745 vp_p.n5744 0.005
R27152 vp_p.n5731 vp_p.n5730 0.005
R27153 vp_p.n5717 vp_p.n5716 0.005
R27154 vp_p.n5703 vp_p.n5702 0.005
R27155 vp_p.n5689 vp_p.n5688 0.005
R27156 vp_p.n5675 vp_p.n5674 0.005
R27157 vp_p.n5661 vp_p.n5660 0.005
R27158 vp_p.n5647 vp_p.n5646 0.005
R27159 vp_p.n5633 vp_p.n5632 0.005
R27160 vp_p.n5619 vp_p.n5618 0.005
R27161 vp_p.n5605 vp_p.n5604 0.005
R27162 vp_p.n5591 vp_p.n5590 0.005
R27163 vp_p.n5577 vp_p.n5576 0.005
R27164 vp_p.n5563 vp_p.n5562 0.005
R27165 vp_p.n5549 vp_p.n5548 0.005
R27166 vp_p.n5535 vp_p.n5534 0.005
R27167 vp_p.n5521 vp_p.n5520 0.005
R27168 vp_p.n5507 vp_p.n5506 0.005
R27169 vp_p.n5493 vp_p.n5492 0.005
R27170 vp_p.n5479 vp_p.n5478 0.005
R27171 vp_p.n5465 vp_p.n5464 0.005
R27172 vp_p.n5451 vp_p.n5450 0.005
R27173 vp_p.n5437 vp_p.n5436 0.005
R27174 vp_p.n5423 vp_p.n5422 0.005
R27175 vp_p.n5409 vp_p.n5408 0.005
R27176 vp_p.n5395 vp_p.n5394 0.005
R27177 vp_p.n5381 vp_p.n5380 0.005
R27178 vp_p.n5367 vp_p.n5366 0.005
R27179 vp_p.n5353 vp_p.n5352 0.005
R27180 vp_p.n5339 vp_p.n5338 0.005
R27181 vp_p.n5325 vp_p.n5324 0.005
R27182 vp_p.n5311 vp_p.n5310 0.005
R27183 vp_p.n5297 vp_p.n5296 0.005
R27184 vp_p.n5283 vp_p.n5282 0.005
R27185 vp_p.n5269 vp_p.n5268 0.005
R27186 vp_p.n5255 vp_p.n5254 0.005
R27187 vp_p.n5241 vp_p.n5240 0.005
R27188 vp_p.n5227 vp_p.n5226 0.005
R27189 vp_p.n5213 vp_p.n5212 0.005
R27190 vp_p.n5199 vp_p.n5198 0.005
R27191 vp_p.n5185 vp_p.n5184 0.005
R27192 vp_p.n5171 vp_p.n5170 0.005
R27193 vp_p.n5157 vp_p.n5156 0.005
R27194 vp_p.n5143 vp_p.n5142 0.005
R27195 vp_p.n5129 vp_p.n5128 0.005
R27196 vp_p.n5115 vp_p.n5114 0.005
R27197 vp_p.n5101 vp_p.n5100 0.005
R27198 vp_p.n5087 vp_p.n5086 0.005
R27199 vp_p.n5073 vp_p.n5072 0.005
R27200 vp_p.n5059 vp_p.n5058 0.005
R27201 vp_p.n5045 vp_p.n5044 0.005
R27202 vp_p.n5031 vp_p.n5030 0.005
R27203 vp_p.n5017 vp_p.n5016 0.005
R27204 vp_p.n5003 vp_p.n5002 0.005
R27205 vp_p.n4989 vp_p.n4988 0.005
R27206 vp_p.n4975 vp_p.n4974 0.005
R27207 vp_p.n4961 vp_p.n4960 0.005
R27208 vp_p.n4947 vp_p.n4946 0.005
R27209 vp_p.n4933 vp_p.n4932 0.005
R27210 vp_p.n4919 vp_p.n4918 0.005
R27211 vp_p.n4905 vp_p.n4904 0.005
R27212 vp_p.n4891 vp_p.n4890 0.005
R27213 vp_p.n4877 vp_p.n4876 0.005
R27214 vp_p.n4863 vp_p.n4862 0.005
R27215 vp_p.n4849 vp_p.n4848 0.005
R27216 vp_p.n4835 vp_p.n4834 0.005
R27217 vp_p.n4821 vp_p.n4820 0.005
R27218 vp_p.n4807 vp_p.n4806 0.005
R27219 vp_p.n4793 vp_p.n4792 0.005
R27220 vp_p.n4779 vp_p.n4778 0.005
R27221 vp_p.n4765 vp_p.n4764 0.005
R27222 vp_p.n4751 vp_p.n4750 0.005
R27223 vp_p.n24447 vp_p.n24446 0.005
R27224 vp_p.n24433 vp_p.n24432 0.005
R27225 vp_p.n24419 vp_p.n24418 0.005
R27226 vp_p.n24405 vp_p.n24404 0.005
R27227 vp_p.n24391 vp_p.n24390 0.005
R27228 vp_p.n24377 vp_p.n24376 0.005
R27229 vp_p.n24363 vp_p.n24362 0.005
R27230 vp_p.n24349 vp_p.n24348 0.005
R27231 vp_p.n24335 vp_p.n24334 0.005
R27232 vp_p.n24321 vp_p.n24320 0.005
R27233 vp_p.n24307 vp_p.n24306 0.005
R27234 vp_p.n24293 vp_p.n24292 0.005
R27235 vp_p.n24279 vp_p.n24278 0.005
R27236 vp_p.n24265 vp_p.n24264 0.005
R27237 vp_p.n24251 vp_p.n24250 0.005
R27238 vp_p.n24237 vp_p.n24236 0.005
R27239 vp_p.n24223 vp_p.n24222 0.005
R27240 vp_p.n24209 vp_p.n24208 0.005
R27241 vp_p.n24195 vp_p.n24194 0.005
R27242 vp_p.n24181 vp_p.n24180 0.005
R27243 vp_p.n24167 vp_p.n24166 0.005
R27244 vp_p.n24153 vp_p.n24152 0.005
R27245 vp_p.n24139 vp_p.n24138 0.005
R27246 vp_p.n24125 vp_p.n24124 0.005
R27247 vp_p.n24111 vp_p.n24110 0.005
R27248 vp_p.n24097 vp_p.n24096 0.005
R27249 vp_p.n24083 vp_p.n24082 0.005
R27250 vp_p.n24069 vp_p.n24068 0.005
R27251 vp_p.n24055 vp_p.n24054 0.005
R27252 vp_p.n24041 vp_p.n24040 0.005
R27253 vp_p.n24027 vp_p.n24026 0.005
R27254 vp_p.n24013 vp_p.n24012 0.005
R27255 vp_p.n23999 vp_p.n23998 0.005
R27256 vp_p.n23985 vp_p.n23984 0.005
R27257 vp_p.n23971 vp_p.n23970 0.005
R27258 vp_p.n23957 vp_p.n23956 0.005
R27259 vp_p.n23943 vp_p.n23942 0.005
R27260 vp_p.n23929 vp_p.n23928 0.005
R27261 vp_p.n23915 vp_p.n23914 0.005
R27262 vp_p.n23901 vp_p.n23900 0.005
R27263 vp_p.n23887 vp_p.n23886 0.005
R27264 vp_p.n23873 vp_p.n23872 0.005
R27265 vp_p.n23859 vp_p.n23858 0.005
R27266 vp_p.n23845 vp_p.n23844 0.005
R27267 vp_p.n23831 vp_p.n23830 0.005
R27268 vp_p.n23817 vp_p.n23816 0.005
R27269 vp_p.n23803 vp_p.n23802 0.005
R27270 vp_p.n23789 vp_p.n23788 0.005
R27271 vp_p.n23775 vp_p.n23774 0.005
R27272 vp_p.n23761 vp_p.n23760 0.005
R27273 vp_p.n23747 vp_p.n23746 0.005
R27274 vp_p.n23733 vp_p.n23732 0.005
R27275 vp_p.n23719 vp_p.n23718 0.005
R27276 vp_p.n23705 vp_p.n23704 0.005
R27277 vp_p.n23691 vp_p.n23690 0.005
R27278 vp_p.n23677 vp_p.n23676 0.005
R27279 vp_p.n23663 vp_p.n23662 0.005
R27280 vp_p.n23649 vp_p.n23648 0.005
R27281 vp_p.n23635 vp_p.n23634 0.005
R27282 vp_p.n23621 vp_p.n23620 0.005
R27283 vp_p.n23607 vp_p.n23606 0.005
R27284 vp_p.n23593 vp_p.n23592 0.005
R27285 vp_p.n23579 vp_p.n23578 0.005
R27286 vp_p.n23565 vp_p.n23564 0.005
R27287 vp_p.n23551 vp_p.n23550 0.005
R27288 vp_p.n23537 vp_p.n23536 0.005
R27289 vp_p.n23523 vp_p.n23522 0.005
R27290 vp_p.n23509 vp_p.n23508 0.005
R27291 vp_p.n23495 vp_p.n23494 0.005
R27292 vp_p.n23481 vp_p.n23480 0.005
R27293 vp_p.n23467 vp_p.n23466 0.005
R27294 vp_p.n23453 vp_p.n23452 0.005
R27295 vp_p.n7182 vp_p.n7181 0.005
R27296 vp_p.n7168 vp_p.n7167 0.005
R27297 vp_p.n7154 vp_p.n7153 0.005
R27298 vp_p.n7140 vp_p.n7139 0.005
R27299 vp_p.n7126 vp_p.n7125 0.005
R27300 vp_p.n7112 vp_p.n7111 0.005
R27301 vp_p.n7098 vp_p.n7097 0.005
R27302 vp_p.n7084 vp_p.n7083 0.005
R27303 vp_p.n7070 vp_p.n7069 0.005
R27304 vp_p.n7056 vp_p.n7055 0.005
R27305 vp_p.n7042 vp_p.n7041 0.005
R27306 vp_p.n7028 vp_p.n7027 0.005
R27307 vp_p.n7014 vp_p.n7013 0.005
R27308 vp_p.n7000 vp_p.n6999 0.005
R27309 vp_p.n6986 vp_p.n6985 0.005
R27310 vp_p.n6972 vp_p.n6971 0.005
R27311 vp_p.n6958 vp_p.n6957 0.005
R27312 vp_p.n6944 vp_p.n6943 0.005
R27313 vp_p.n6930 vp_p.n6929 0.005
R27314 vp_p.n6916 vp_p.n6915 0.005
R27315 vp_p.n6902 vp_p.n6901 0.005
R27316 vp_p.n6888 vp_p.n6887 0.005
R27317 vp_p.n6874 vp_p.n6873 0.005
R27318 vp_p.n6860 vp_p.n6859 0.005
R27319 vp_p.n6846 vp_p.n6845 0.005
R27320 vp_p.n6832 vp_p.n6831 0.005
R27321 vp_p.n6818 vp_p.n6817 0.005
R27322 vp_p.n6804 vp_p.n6803 0.005
R27323 vp_p.n6790 vp_p.n6789 0.005
R27324 vp_p.n6776 vp_p.n6775 0.005
R27325 vp_p.n6762 vp_p.n6761 0.005
R27326 vp_p.n6748 vp_p.n6747 0.005
R27327 vp_p.n6734 vp_p.n6733 0.005
R27328 vp_p.n6720 vp_p.n6719 0.005
R27329 vp_p.n6706 vp_p.n6705 0.005
R27330 vp_p.n6692 vp_p.n6691 0.005
R27331 vp_p.n6678 vp_p.n6677 0.005
R27332 vp_p.n6664 vp_p.n6663 0.005
R27333 vp_p.n6650 vp_p.n6649 0.005
R27334 vp_p.n6636 vp_p.n6635 0.005
R27335 vp_p.n6622 vp_p.n6621 0.005
R27336 vp_p.n6608 vp_p.n6607 0.005
R27337 vp_p.n6594 vp_p.n6593 0.005
R27338 vp_p.n6580 vp_p.n6579 0.005
R27339 vp_p.n6566 vp_p.n6565 0.005
R27340 vp_p.n6552 vp_p.n6551 0.005
R27341 vp_p.n6538 vp_p.n6537 0.005
R27342 vp_p.n6524 vp_p.n6523 0.005
R27343 vp_p.n6510 vp_p.n6509 0.005
R27344 vp_p.n6496 vp_p.n6495 0.005
R27345 vp_p.n6482 vp_p.n6481 0.005
R27346 vp_p.n6468 vp_p.n6467 0.005
R27347 vp_p.n6454 vp_p.n6453 0.005
R27348 vp_p.n6440 vp_p.n6439 0.005
R27349 vp_p.n6426 vp_p.n6425 0.005
R27350 vp_p.n6412 vp_p.n6411 0.005
R27351 vp_p.n6398 vp_p.n6397 0.005
R27352 vp_p.n6384 vp_p.n6383 0.005
R27353 vp_p.n6370 vp_p.n6369 0.005
R27354 vp_p.n6356 vp_p.n6355 0.005
R27355 vp_p.n6342 vp_p.n6341 0.005
R27356 vp_p.n6328 vp_p.n6327 0.005
R27357 vp_p.n6314 vp_p.n6313 0.005
R27358 vp_p.n6300 vp_p.n6299 0.005
R27359 vp_p.n6286 vp_p.n6285 0.005
R27360 vp_p.n6272 vp_p.n6271 0.005
R27361 vp_p.n6258 vp_p.n6257 0.005
R27362 vp_p.n6244 vp_p.n6243 0.005
R27363 vp_p.n6230 vp_p.n6229 0.005
R27364 vp_p.n6216 vp_p.n6215 0.005
R27365 vp_p.n6202 vp_p.n6201 0.005
R27366 vp_p.n6188 vp_p.n6187 0.005
R27367 vp_p.n6174 vp_p.n6173 0.005
R27368 vp_p.n25883 vp_p.n25882 0.005
R27369 vp_p.n25869 vp_p.n25868 0.005
R27370 vp_p.n25855 vp_p.n25854 0.005
R27371 vp_p.n25841 vp_p.n25840 0.005
R27372 vp_p.n25827 vp_p.n25826 0.005
R27373 vp_p.n25813 vp_p.n25812 0.005
R27374 vp_p.n25799 vp_p.n25798 0.005
R27375 vp_p.n25785 vp_p.n25784 0.005
R27376 vp_p.n25771 vp_p.n25770 0.005
R27377 vp_p.n25757 vp_p.n25756 0.005
R27378 vp_p.n25743 vp_p.n25742 0.005
R27379 vp_p.n25729 vp_p.n25728 0.005
R27380 vp_p.n25715 vp_p.n25714 0.005
R27381 vp_p.n25701 vp_p.n25700 0.005
R27382 vp_p.n25687 vp_p.n25686 0.005
R27383 vp_p.n25673 vp_p.n25672 0.005
R27384 vp_p.n25659 vp_p.n25658 0.005
R27385 vp_p.n25645 vp_p.n25644 0.005
R27386 vp_p.n25631 vp_p.n25630 0.005
R27387 vp_p.n25617 vp_p.n25616 0.005
R27388 vp_p.n25603 vp_p.n25602 0.005
R27389 vp_p.n25589 vp_p.n25588 0.005
R27390 vp_p.n25575 vp_p.n25574 0.005
R27391 vp_p.n25561 vp_p.n25560 0.005
R27392 vp_p.n25547 vp_p.n25546 0.005
R27393 vp_p.n25533 vp_p.n25532 0.005
R27394 vp_p.n25519 vp_p.n25518 0.005
R27395 vp_p.n25505 vp_p.n25504 0.005
R27396 vp_p.n25491 vp_p.n25490 0.005
R27397 vp_p.n25477 vp_p.n25476 0.005
R27398 vp_p.n25463 vp_p.n25462 0.005
R27399 vp_p.n25449 vp_p.n25448 0.005
R27400 vp_p.n25435 vp_p.n25434 0.005
R27401 vp_p.n25421 vp_p.n25420 0.005
R27402 vp_p.n25407 vp_p.n25406 0.005
R27403 vp_p.n25393 vp_p.n25392 0.005
R27404 vp_p.n25379 vp_p.n25378 0.005
R27405 vp_p.n25365 vp_p.n25364 0.005
R27406 vp_p.n25351 vp_p.n25350 0.005
R27407 vp_p.n25337 vp_p.n25336 0.005
R27408 vp_p.n25323 vp_p.n25322 0.005
R27409 vp_p.n25309 vp_p.n25308 0.005
R27410 vp_p.n25295 vp_p.n25294 0.005
R27411 vp_p.n25281 vp_p.n25280 0.005
R27412 vp_p.n25267 vp_p.n25266 0.005
R27413 vp_p.n25253 vp_p.n25252 0.005
R27414 vp_p.n25239 vp_p.n25238 0.005
R27415 vp_p.n25225 vp_p.n25224 0.005
R27416 vp_p.n25211 vp_p.n25210 0.005
R27417 vp_p.n25197 vp_p.n25196 0.005
R27418 vp_p.n25183 vp_p.n25182 0.005
R27419 vp_p.n25169 vp_p.n25168 0.005
R27420 vp_p.n25155 vp_p.n25154 0.005
R27421 vp_p.n25141 vp_p.n25140 0.005
R27422 vp_p.n25127 vp_p.n25126 0.005
R27423 vp_p.n25113 vp_p.n25112 0.005
R27424 vp_p.n25099 vp_p.n25098 0.005
R27425 vp_p.n25085 vp_p.n25084 0.005
R27426 vp_p.n25071 vp_p.n25070 0.005
R27427 vp_p.n25057 vp_p.n25056 0.005
R27428 vp_p.n25043 vp_p.n25042 0.005
R27429 vp_p.n25029 vp_p.n25028 0.005
R27430 vp_p.n25015 vp_p.n25014 0.005
R27431 vp_p.n25001 vp_p.n25000 0.005
R27432 vp_p.n24987 vp_p.n24986 0.005
R27433 vp_p.n24973 vp_p.n24972 0.005
R27434 vp_p.n24959 vp_p.n24958 0.005
R27435 vp_p.n24945 vp_p.n24944 0.005
R27436 vp_p.n24931 vp_p.n24930 0.005
R27437 vp_p.n24917 vp_p.n24916 0.005
R27438 vp_p.n24903 vp_p.n24902 0.005
R27439 vp_p.n24889 vp_p.n24888 0.005
R27440 vp_p.n24875 vp_p.n24874 0.005
R27441 vp_p.n7596 vp_p.n7595 0.005
R27442 vp_p.n7610 vp_p.n7609 0.005
R27443 vp_p.n7624 vp_p.n7623 0.005
R27444 vp_p.n7638 vp_p.n7637 0.005
R27445 vp_p.n7652 vp_p.n7651 0.005
R27446 vp_p.n7666 vp_p.n7665 0.005
R27447 vp_p.n7680 vp_p.n7679 0.005
R27448 vp_p.n7694 vp_p.n7693 0.005
R27449 vp_p.n7708 vp_p.n7707 0.005
R27450 vp_p.n7722 vp_p.n7721 0.005
R27451 vp_p.n7736 vp_p.n7735 0.005
R27452 vp_p.n7750 vp_p.n7749 0.005
R27453 vp_p.n7764 vp_p.n7763 0.005
R27454 vp_p.n7778 vp_p.n7777 0.005
R27455 vp_p.n7792 vp_p.n7791 0.005
R27456 vp_p.n7806 vp_p.n7805 0.005
R27457 vp_p.n7820 vp_p.n7819 0.005
R27458 vp_p.n7834 vp_p.n7833 0.005
R27459 vp_p.n7848 vp_p.n7847 0.005
R27460 vp_p.n7862 vp_p.n7861 0.005
R27461 vp_p.n7876 vp_p.n7875 0.005
R27462 vp_p.n7890 vp_p.n7889 0.005
R27463 vp_p.n7904 vp_p.n7903 0.005
R27464 vp_p.n7918 vp_p.n7917 0.005
R27465 vp_p.n7932 vp_p.n7931 0.005
R27466 vp_p.n7946 vp_p.n7945 0.005
R27467 vp_p.n7960 vp_p.n7959 0.005
R27468 vp_p.n7974 vp_p.n7973 0.005
R27469 vp_p.n7988 vp_p.n7987 0.005
R27470 vp_p.n8002 vp_p.n8001 0.005
R27471 vp_p.n8016 vp_p.n8015 0.005
R27472 vp_p.n8030 vp_p.n8029 0.005
R27473 vp_p.n8044 vp_p.n8043 0.005
R27474 vp_p.n8058 vp_p.n8057 0.005
R27475 vp_p.n8072 vp_p.n8071 0.005
R27476 vp_p.n8086 vp_p.n8085 0.005
R27477 vp_p.n8100 vp_p.n8099 0.005
R27478 vp_p.n8114 vp_p.n8113 0.005
R27479 vp_p.n8128 vp_p.n8127 0.005
R27480 vp_p.n8142 vp_p.n8141 0.005
R27481 vp_p.n8156 vp_p.n8155 0.005
R27482 vp_p.n8170 vp_p.n8169 0.005
R27483 vp_p.n8184 vp_p.n8183 0.005
R27484 vp_p.n8198 vp_p.n8197 0.005
R27485 vp_p.n8212 vp_p.n8211 0.005
R27486 vp_p.n8226 vp_p.n8225 0.005
R27487 vp_p.n8240 vp_p.n8239 0.005
R27488 vp_p.n8254 vp_p.n8253 0.005
R27489 vp_p.n8268 vp_p.n8267 0.005
R27490 vp_p.n8282 vp_p.n8281 0.005
R27491 vp_p.n8296 vp_p.n8295 0.005
R27492 vp_p.n8310 vp_p.n8309 0.005
R27493 vp_p.n8324 vp_p.n8323 0.005
R27494 vp_p.n8338 vp_p.n8337 0.005
R27495 vp_p.n8352 vp_p.n8351 0.005
R27496 vp_p.n8366 vp_p.n8365 0.005
R27497 vp_p.n8380 vp_p.n8379 0.005
R27498 vp_p.n8394 vp_p.n8393 0.005
R27499 vp_p.n8408 vp_p.n8407 0.005
R27500 vp_p.n8422 vp_p.n8421 0.005
R27501 vp_p.n8436 vp_p.n8435 0.005
R27502 vp_p.n8450 vp_p.n8449 0.005
R27503 vp_p.n8464 vp_p.n8463 0.005
R27504 vp_p.n8478 vp_p.n8477 0.005
R27505 vp_p.n8492 vp_p.n8491 0.005
R27506 vp_p.n8506 vp_p.n8505 0.005
R27507 vp_p.n8520 vp_p.n8519 0.005
R27508 vp_p.n8534 vp_p.n8533 0.005
R27509 vp_p.n8548 vp_p.n8547 0.005
R27510 vp_p.n8562 vp_p.n8561 0.005
R27511 vp_p.n8576 vp_p.n8575 0.005
R27512 vp_p.n8590 vp_p.n8589 0.005
R27513 vp_p.n8604 vp_p.n8603 0.005
R27514 vp_p.n8618 vp_p.n8617 0.005
R27515 vp_p.n26300 vp_p.n26299 0.005
R27516 vp_p.n26314 vp_p.n26313 0.005
R27517 vp_p.n26328 vp_p.n26327 0.005
R27518 vp_p.n26342 vp_p.n26341 0.005
R27519 vp_p.n26356 vp_p.n26355 0.005
R27520 vp_p.n26370 vp_p.n26369 0.005
R27521 vp_p.n26384 vp_p.n26383 0.005
R27522 vp_p.n26398 vp_p.n26397 0.005
R27523 vp_p.n26412 vp_p.n26411 0.005
R27524 vp_p.n26426 vp_p.n26425 0.005
R27525 vp_p.n26440 vp_p.n26439 0.005
R27526 vp_p.n26454 vp_p.n26453 0.005
R27527 vp_p.n26468 vp_p.n26467 0.005
R27528 vp_p.n26482 vp_p.n26481 0.005
R27529 vp_p.n26496 vp_p.n26495 0.005
R27530 vp_p.n26510 vp_p.n26509 0.005
R27531 vp_p.n26524 vp_p.n26523 0.005
R27532 vp_p.n26538 vp_p.n26537 0.005
R27533 vp_p.n26552 vp_p.n26551 0.005
R27534 vp_p.n26566 vp_p.n26565 0.005
R27535 vp_p.n26580 vp_p.n26579 0.005
R27536 vp_p.n26594 vp_p.n26593 0.005
R27537 vp_p.n26608 vp_p.n26607 0.005
R27538 vp_p.n26622 vp_p.n26621 0.005
R27539 vp_p.n26636 vp_p.n26635 0.005
R27540 vp_p.n26650 vp_p.n26649 0.005
R27541 vp_p.n26664 vp_p.n26663 0.005
R27542 vp_p.n26678 vp_p.n26677 0.005
R27543 vp_p.n26692 vp_p.n26691 0.005
R27544 vp_p.n26706 vp_p.n26705 0.005
R27545 vp_p.n26720 vp_p.n26719 0.005
R27546 vp_p.n26734 vp_p.n26733 0.005
R27547 vp_p.n26748 vp_p.n26747 0.005
R27548 vp_p.n26762 vp_p.n26761 0.005
R27549 vp_p.n26776 vp_p.n26775 0.005
R27550 vp_p.n26790 vp_p.n26789 0.005
R27551 vp_p.n26804 vp_p.n26803 0.005
R27552 vp_p.n26818 vp_p.n26817 0.005
R27553 vp_p.n26832 vp_p.n26831 0.005
R27554 vp_p.n26846 vp_p.n26845 0.005
R27555 vp_p.n26860 vp_p.n26859 0.005
R27556 vp_p.n26874 vp_p.n26873 0.005
R27557 vp_p.n26888 vp_p.n26887 0.005
R27558 vp_p.n26902 vp_p.n26901 0.005
R27559 vp_p.n26916 vp_p.n26915 0.005
R27560 vp_p.n26930 vp_p.n26929 0.005
R27561 vp_p.n26944 vp_p.n26943 0.005
R27562 vp_p.n26958 vp_p.n26957 0.005
R27563 vp_p.n26972 vp_p.n26971 0.005
R27564 vp_p.n26986 vp_p.n26985 0.005
R27565 vp_p.n27000 vp_p.n26999 0.005
R27566 vp_p.n27014 vp_p.n27013 0.005
R27567 vp_p.n27028 vp_p.n27027 0.005
R27568 vp_p.n27042 vp_p.n27041 0.005
R27569 vp_p.n27056 vp_p.n27055 0.005
R27570 vp_p.n27070 vp_p.n27069 0.005
R27571 vp_p.n27084 vp_p.n27083 0.005
R27572 vp_p.n27098 vp_p.n27097 0.005
R27573 vp_p.n27112 vp_p.n27111 0.005
R27574 vp_p.n27126 vp_p.n27125 0.005
R27575 vp_p.n27140 vp_p.n27139 0.005
R27576 vp_p.n27154 vp_p.n27153 0.005
R27577 vp_p.n27168 vp_p.n27167 0.005
R27578 vp_p.n27182 vp_p.n27181 0.005
R27579 vp_p.n27196 vp_p.n27195 0.005
R27580 vp_p.n27210 vp_p.n27209 0.005
R27581 vp_p.n27224 vp_p.n27223 0.005
R27582 vp_p.n27238 vp_p.n27237 0.005
R27583 vp_p.n27252 vp_p.n27251 0.005
R27584 vp_p.n27266 vp_p.n27265 0.005
R27585 vp_p.n27280 vp_p.n27279 0.005
R27586 vp_p.n27294 vp_p.n27293 0.005
R27587 vp_p.n27308 vp_p.n27307 0.005
R27588 vp_p.n27322 vp_p.n27321 0.005
R27589 vp_p.n14384 vp_p.n14383 0.002
R27590 vp_p.n15827 vp_p.n15826 0.002
R27591 vp_p.n17269 vp_p.n17268 0.002
R27592 vp_p.n18710 vp_p.n18709 0.002
R27593 vp_p.n20150 vp_p.n20149 0.002
R27594 vp_p.n21589 vp_p.n21588 0.002
R27595 vp_p.n23027 vp_p.n23026 0.002
R27596 vp_p.n24464 vp_p.n24463 0.002
R27597 vp_p.n25900 vp_p.n25899 0.002
R27598 vp_p.n7585 vp_p.n7584 0.002
R27599 vp_p.n13020 vp_p.n13019 0.002
R27600 vp_p.n11596 vp_p.n11595 0.002
R27601 vp_p.n10173 vp_p.n10172 0.002
R27602 vp_p.n1441 vp_p.n1440 0.002
R27603 vp_p.n2881 vp_p.n2880 0.002
R27604 vp_p.n4320 vp_p.n4319 0.002
R27605 vp_p.n5758 vp_p.n5757 0.002
R27606 vp_p.n7195 vp_p.n7194 0.002
R27607 vp_p.n26285 vp_p.n26284 0.002
R27608 vp_p.n8608 vp_p.n7207 0.001
R27609 vp_p.n7172 vp_p.n5790 0.001
R27610 vp_p.n8594 vp_p.n7212 0.001
R27611 vp_p.n5735 vp_p.n4372 0.001
R27612 vp_p.n7158 vp_p.n5795 0.001
R27613 vp_p.n8580 vp_p.n7217 0.001
R27614 vp_p.n4297 vp_p.n2953 0.001
R27615 vp_p.n5721 vp_p.n4377 0.001
R27616 vp_p.n7144 vp_p.n5800 0.001
R27617 vp_p.n8566 vp_p.n7222 0.001
R27618 vp_p.n2858 vp_p.n1533 0.001
R27619 vp_p.n4283 vp_p.n2958 0.001
R27620 vp_p.n5707 vp_p.n4382 0.001
R27621 vp_p.n7130 vp_p.n5805 0.001
R27622 vp_p.n8552 vp_p.n7227 0.001
R27623 vp_p.n1418 vp_p.n54 0.001
R27624 vp_p.n2844 vp_p.n1538 0.001
R27625 vp_p.n4269 vp_p.n2963 0.001
R27626 vp_p.n5693 vp_p.n4387 0.001
R27627 vp_p.n7116 vp_p.n5810 0.001
R27628 vp_p.n8538 vp_p.n7232 0.001
R27629 vp_p.n10150 vp_p.n8798 0.001
R27630 vp_p.n1404 vp_p.n59 0.001
R27631 vp_p.n2830 vp_p.n1543 0.001
R27632 vp_p.n4255 vp_p.n2968 0.001
R27633 vp_p.n5679 vp_p.n4392 0.001
R27634 vp_p.n7102 vp_p.n5815 0.001
R27635 vp_p.n8524 vp_p.n7237 0.001
R27636 vp_p.n11573 vp_p.n10305 0.001
R27637 vp_p.n10136 vp_p.n8803 0.001
R27638 vp_p.n1390 vp_p.n64 0.001
R27639 vp_p.n2816 vp_p.n1548 0.001
R27640 vp_p.n4241 vp_p.n2973 0.001
R27641 vp_p.n5665 vp_p.n4397 0.001
R27642 vp_p.n7088 vp_p.n5820 0.001
R27643 vp_p.n8510 vp_p.n7242 0.001
R27644 vp_p.n13855 vp_p.n13832 0.001
R27645 vp_p.n12101 vp_p.n12068 0.001
R27646 vp_p.n10663 vp_p.n10630 0.001
R27647 vp_p.n9226 vp_p.n9128 0.001
R27648 vp_p.n480 vp_p.n389 0.001
R27649 vp_p.n1906 vp_p.n1873 0.001
R27650 vp_p.n3331 vp_p.n3298 0.001
R27651 vp_p.n4755 vp_p.n4722 0.001
R27652 vp_p.n6178 vp_p.n6145 0.001
R27653 vp_p.n7600 vp_p.n7567 0.001
R27654 vp_p.n14904 vp_p.n14871 0.001
R27655 vp_p.n16332 vp_p.n16299 0.001
R27656 vp_p.n17759 vp_p.n17726 0.001
R27657 vp_p.n19185 vp_p.n19152 0.001
R27658 vp_p.n20610 vp_p.n20577 0.001
R27659 vp_p.n22034 vp_p.n22001 0.001
R27660 vp_p.n23457 vp_p.n23424 0.001
R27661 vp_p.n24879 vp_p.n24846 0.001
R27662 vp_p.n26304 vp_p.n26272 0.001
R27663 vp_p.n13859 vp_p.n13827 0.001
R27664 vp_p.n13863 vp_p.n13822 0.001
R27665 vp_p.n12115 vp_p.n12063 0.001
R27666 vp_p.n10677 vp_p.n10625 0.001
R27667 vp_p.n9240 vp_p.n9123 0.001
R27668 vp_p.n494 vp_p.n384 0.001
R27669 vp_p.n1920 vp_p.n1868 0.001
R27670 vp_p.n3345 vp_p.n3293 0.001
R27671 vp_p.n4769 vp_p.n4717 0.001
R27672 vp_p.n6192 vp_p.n6140 0.001
R27673 vp_p.n7614 vp_p.n7562 0.001
R27674 vp_p.n14918 vp_p.n14866 0.001
R27675 vp_p.n16346 vp_p.n16294 0.001
R27676 vp_p.n17773 vp_p.n17721 0.001
R27677 vp_p.n19199 vp_p.n19147 0.001
R27678 vp_p.n20624 vp_p.n20572 0.001
R27679 vp_p.n22048 vp_p.n21996 0.001
R27680 vp_p.n23471 vp_p.n23419 0.001
R27681 vp_p.n24893 vp_p.n24841 0.001
R27682 vp_p.n26318 vp_p.n26267 0.001
R27683 vp_p.n13867 vp_p.n13817 0.001
R27684 vp_p.n13871 vp_p.n13812 0.001
R27685 vp_p.n12129 vp_p.n12058 0.001
R27686 vp_p.n10691 vp_p.n10620 0.001
R27687 vp_p.n9254 vp_p.n9118 0.001
R27688 vp_p.n508 vp_p.n379 0.001
R27689 vp_p.n1934 vp_p.n1863 0.001
R27690 vp_p.n3359 vp_p.n3288 0.001
R27691 vp_p.n4783 vp_p.n4712 0.001
R27692 vp_p.n6206 vp_p.n6135 0.001
R27693 vp_p.n7628 vp_p.n7557 0.001
R27694 vp_p.n14932 vp_p.n14861 0.001
R27695 vp_p.n16360 vp_p.n16289 0.001
R27696 vp_p.n17787 vp_p.n17716 0.001
R27697 vp_p.n19213 vp_p.n19142 0.001
R27698 vp_p.n20638 vp_p.n20567 0.001
R27699 vp_p.n22062 vp_p.n21991 0.001
R27700 vp_p.n23485 vp_p.n23414 0.001
R27701 vp_p.n24907 vp_p.n24836 0.001
R27702 vp_p.n26332 vp_p.n26262 0.001
R27703 vp_p.n13875 vp_p.n13807 0.001
R27704 vp_p.n13879 vp_p.n13802 0.001
R27705 vp_p.n12143 vp_p.n12053 0.001
R27706 vp_p.n10705 vp_p.n10615 0.001
R27707 vp_p.n9268 vp_p.n9113 0.001
R27708 vp_p.n522 vp_p.n374 0.001
R27709 vp_p.n1948 vp_p.n1858 0.001
R27710 vp_p.n3373 vp_p.n3283 0.001
R27711 vp_p.n4797 vp_p.n4707 0.001
R27712 vp_p.n6220 vp_p.n6130 0.001
R27713 vp_p.n7642 vp_p.n7552 0.001
R27714 vp_p.n14946 vp_p.n14856 0.001
R27715 vp_p.n16374 vp_p.n16284 0.001
R27716 vp_p.n17801 vp_p.n17711 0.001
R27717 vp_p.n19227 vp_p.n19137 0.001
R27718 vp_p.n20652 vp_p.n20562 0.001
R27719 vp_p.n22076 vp_p.n21986 0.001
R27720 vp_p.n23499 vp_p.n23409 0.001
R27721 vp_p.n24921 vp_p.n24831 0.001
R27722 vp_p.n26346 vp_p.n26257 0.001
R27723 vp_p.n13883 vp_p.n13797 0.001
R27724 vp_p.n13887 vp_p.n13792 0.001
R27725 vp_p.n12157 vp_p.n12048 0.001
R27726 vp_p.n10719 vp_p.n10610 0.001
R27727 vp_p.n9282 vp_p.n9108 0.001
R27728 vp_p.n536 vp_p.n369 0.001
R27729 vp_p.n1962 vp_p.n1853 0.001
R27730 vp_p.n3387 vp_p.n3278 0.001
R27731 vp_p.n4811 vp_p.n4702 0.001
R27732 vp_p.n6234 vp_p.n6125 0.001
R27733 vp_p.n7656 vp_p.n7547 0.001
R27734 vp_p.n14960 vp_p.n14851 0.001
R27735 vp_p.n16388 vp_p.n16279 0.001
R27736 vp_p.n17815 vp_p.n17706 0.001
R27737 vp_p.n19241 vp_p.n19132 0.001
R27738 vp_p.n20666 vp_p.n20557 0.001
R27739 vp_p.n22090 vp_p.n21981 0.001
R27740 vp_p.n23513 vp_p.n23404 0.001
R27741 vp_p.n24935 vp_p.n24826 0.001
R27742 vp_p.n26360 vp_p.n26252 0.001
R27743 vp_p.n13891 vp_p.n13787 0.001
R27744 vp_p.n13895 vp_p.n13782 0.001
R27745 vp_p.n12171 vp_p.n12043 0.001
R27746 vp_p.n10733 vp_p.n10605 0.001
R27747 vp_p.n9296 vp_p.n9103 0.001
R27748 vp_p.n550 vp_p.n364 0.001
R27749 vp_p.n1976 vp_p.n1848 0.001
R27750 vp_p.n3401 vp_p.n3273 0.001
R27751 vp_p.n4825 vp_p.n4697 0.001
R27752 vp_p.n6248 vp_p.n6120 0.001
R27753 vp_p.n7670 vp_p.n7542 0.001
R27754 vp_p.n14974 vp_p.n14846 0.001
R27755 vp_p.n16402 vp_p.n16274 0.001
R27756 vp_p.n17829 vp_p.n17701 0.001
R27757 vp_p.n19255 vp_p.n19127 0.001
R27758 vp_p.n20680 vp_p.n20552 0.001
R27759 vp_p.n22104 vp_p.n21976 0.001
R27760 vp_p.n23527 vp_p.n23399 0.001
R27761 vp_p.n24949 vp_p.n24821 0.001
R27762 vp_p.n26374 vp_p.n26247 0.001
R27763 vp_p.n13899 vp_p.n13777 0.001
R27764 vp_p.n13903 vp_p.n13772 0.001
R27765 vp_p.n12185 vp_p.n12038 0.001
R27766 vp_p.n10747 vp_p.n10600 0.001
R27767 vp_p.n9310 vp_p.n9098 0.001
R27768 vp_p.n564 vp_p.n359 0.001
R27769 vp_p.n1990 vp_p.n1843 0.001
R27770 vp_p.n3415 vp_p.n3268 0.001
R27771 vp_p.n4839 vp_p.n4692 0.001
R27772 vp_p.n6262 vp_p.n6115 0.001
R27773 vp_p.n7684 vp_p.n7537 0.001
R27774 vp_p.n14988 vp_p.n14841 0.001
R27775 vp_p.n16416 vp_p.n16269 0.001
R27776 vp_p.n17843 vp_p.n17696 0.001
R27777 vp_p.n19269 vp_p.n19122 0.001
R27778 vp_p.n20694 vp_p.n20547 0.001
R27779 vp_p.n22118 vp_p.n21971 0.001
R27780 vp_p.n23541 vp_p.n23394 0.001
R27781 vp_p.n24963 vp_p.n24816 0.001
R27782 vp_p.n26388 vp_p.n26242 0.001
R27783 vp_p.n13907 vp_p.n13767 0.001
R27784 vp_p.n13911 vp_p.n13762 0.001
R27785 vp_p.n12199 vp_p.n12033 0.001
R27786 vp_p.n10761 vp_p.n10595 0.001
R27787 vp_p.n9324 vp_p.n9093 0.001
R27788 vp_p.n578 vp_p.n354 0.001
R27789 vp_p.n2004 vp_p.n1838 0.001
R27790 vp_p.n3429 vp_p.n3263 0.001
R27791 vp_p.n4853 vp_p.n4687 0.001
R27792 vp_p.n6276 vp_p.n6110 0.001
R27793 vp_p.n7698 vp_p.n7532 0.001
R27794 vp_p.n15002 vp_p.n14836 0.001
R27795 vp_p.n16430 vp_p.n16264 0.001
R27796 vp_p.n17857 vp_p.n17691 0.001
R27797 vp_p.n19283 vp_p.n19117 0.001
R27798 vp_p.n20708 vp_p.n20542 0.001
R27799 vp_p.n22132 vp_p.n21966 0.001
R27800 vp_p.n23555 vp_p.n23389 0.001
R27801 vp_p.n24977 vp_p.n24811 0.001
R27802 vp_p.n26402 vp_p.n26237 0.001
R27803 vp_p.n13915 vp_p.n13757 0.001
R27804 vp_p.n13919 vp_p.n13752 0.001
R27805 vp_p.n12213 vp_p.n12028 0.001
R27806 vp_p.n10775 vp_p.n10590 0.001
R27807 vp_p.n9338 vp_p.n9088 0.001
R27808 vp_p.n592 vp_p.n349 0.001
R27809 vp_p.n2018 vp_p.n1833 0.001
R27810 vp_p.n3443 vp_p.n3258 0.001
R27811 vp_p.n4867 vp_p.n4682 0.001
R27812 vp_p.n6290 vp_p.n6105 0.001
R27813 vp_p.n7712 vp_p.n7527 0.001
R27814 vp_p.n15016 vp_p.n14831 0.001
R27815 vp_p.n16444 vp_p.n16259 0.001
R27816 vp_p.n17871 vp_p.n17686 0.001
R27817 vp_p.n19297 vp_p.n19112 0.001
R27818 vp_p.n20722 vp_p.n20537 0.001
R27819 vp_p.n22146 vp_p.n21961 0.001
R27820 vp_p.n23569 vp_p.n23384 0.001
R27821 vp_p.n24991 vp_p.n24806 0.001
R27822 vp_p.n26416 vp_p.n26232 0.001
R27823 vp_p.n13923 vp_p.n13747 0.001
R27824 vp_p.n13927 vp_p.n13742 0.001
R27825 vp_p.n12227 vp_p.n12023 0.001
R27826 vp_p.n10789 vp_p.n10585 0.001
R27827 vp_p.n9352 vp_p.n9083 0.001
R27828 vp_p.n606 vp_p.n344 0.001
R27829 vp_p.n2032 vp_p.n1828 0.001
R27830 vp_p.n3457 vp_p.n3253 0.001
R27831 vp_p.n4881 vp_p.n4677 0.001
R27832 vp_p.n6304 vp_p.n6100 0.001
R27833 vp_p.n7726 vp_p.n7522 0.001
R27834 vp_p.n15030 vp_p.n14826 0.001
R27835 vp_p.n16458 vp_p.n16254 0.001
R27836 vp_p.n17885 vp_p.n17681 0.001
R27837 vp_p.n19311 vp_p.n19107 0.001
R27838 vp_p.n20736 vp_p.n20532 0.001
R27839 vp_p.n22160 vp_p.n21956 0.001
R27840 vp_p.n23583 vp_p.n23379 0.001
R27841 vp_p.n25005 vp_p.n24801 0.001
R27842 vp_p.n26430 vp_p.n26227 0.001
R27843 vp_p.n13931 vp_p.n13737 0.001
R27844 vp_p.n13935 vp_p.n13732 0.001
R27845 vp_p.n12241 vp_p.n12018 0.001
R27846 vp_p.n10803 vp_p.n10580 0.001
R27847 vp_p.n9366 vp_p.n9078 0.001
R27848 vp_p.n620 vp_p.n339 0.001
R27849 vp_p.n2046 vp_p.n1823 0.001
R27850 vp_p.n3471 vp_p.n3248 0.001
R27851 vp_p.n4895 vp_p.n4672 0.001
R27852 vp_p.n6318 vp_p.n6095 0.001
R27853 vp_p.n7740 vp_p.n7517 0.001
R27854 vp_p.n15044 vp_p.n14821 0.001
R27855 vp_p.n16472 vp_p.n16249 0.001
R27856 vp_p.n17899 vp_p.n17676 0.001
R27857 vp_p.n19325 vp_p.n19102 0.001
R27858 vp_p.n20750 vp_p.n20527 0.001
R27859 vp_p.n22174 vp_p.n21951 0.001
R27860 vp_p.n23597 vp_p.n23374 0.001
R27861 vp_p.n25019 vp_p.n24796 0.001
R27862 vp_p.n26444 vp_p.n26222 0.001
R27863 vp_p.n13939 vp_p.n13727 0.001
R27864 vp_p.n13943 vp_p.n13722 0.001
R27865 vp_p.n12255 vp_p.n12013 0.001
R27866 vp_p.n10817 vp_p.n10575 0.001
R27867 vp_p.n9380 vp_p.n9073 0.001
R27868 vp_p.n634 vp_p.n334 0.001
R27869 vp_p.n2060 vp_p.n1818 0.001
R27870 vp_p.n3485 vp_p.n3243 0.001
R27871 vp_p.n4909 vp_p.n4667 0.001
R27872 vp_p.n6332 vp_p.n6090 0.001
R27873 vp_p.n7754 vp_p.n7512 0.001
R27874 vp_p.n15058 vp_p.n14816 0.001
R27875 vp_p.n16486 vp_p.n16244 0.001
R27876 vp_p.n17913 vp_p.n17671 0.001
R27877 vp_p.n19339 vp_p.n19097 0.001
R27878 vp_p.n20764 vp_p.n20522 0.001
R27879 vp_p.n22188 vp_p.n21946 0.001
R27880 vp_p.n23611 vp_p.n23369 0.001
R27881 vp_p.n25033 vp_p.n24791 0.001
R27882 vp_p.n26458 vp_p.n26217 0.001
R27883 vp_p.n13947 vp_p.n13717 0.001
R27884 vp_p.n13951 vp_p.n13712 0.001
R27885 vp_p.n12269 vp_p.n12008 0.001
R27886 vp_p.n10831 vp_p.n10570 0.001
R27887 vp_p.n9394 vp_p.n9068 0.001
R27888 vp_p.n648 vp_p.n329 0.001
R27889 vp_p.n2074 vp_p.n1813 0.001
R27890 vp_p.n3499 vp_p.n3238 0.001
R27891 vp_p.n4923 vp_p.n4662 0.001
R27892 vp_p.n6346 vp_p.n6085 0.001
R27893 vp_p.n7768 vp_p.n7507 0.001
R27894 vp_p.n15072 vp_p.n14811 0.001
R27895 vp_p.n16500 vp_p.n16239 0.001
R27896 vp_p.n17927 vp_p.n17666 0.001
R27897 vp_p.n19353 vp_p.n19092 0.001
R27898 vp_p.n20778 vp_p.n20517 0.001
R27899 vp_p.n22202 vp_p.n21941 0.001
R27900 vp_p.n23625 vp_p.n23364 0.001
R27901 vp_p.n25047 vp_p.n24786 0.001
R27902 vp_p.n26472 vp_p.n26212 0.001
R27903 vp_p.n13955 vp_p.n13707 0.001
R27904 vp_p.n13959 vp_p.n13702 0.001
R27905 vp_p.n12283 vp_p.n12003 0.001
R27906 vp_p.n10845 vp_p.n10565 0.001
R27907 vp_p.n9408 vp_p.n9063 0.001
R27908 vp_p.n662 vp_p.n324 0.001
R27909 vp_p.n2088 vp_p.n1808 0.001
R27910 vp_p.n3513 vp_p.n3233 0.001
R27911 vp_p.n4937 vp_p.n4657 0.001
R27912 vp_p.n6360 vp_p.n6080 0.001
R27913 vp_p.n7782 vp_p.n7502 0.001
R27914 vp_p.n15086 vp_p.n14806 0.001
R27915 vp_p.n16514 vp_p.n16234 0.001
R27916 vp_p.n17941 vp_p.n17661 0.001
R27917 vp_p.n19367 vp_p.n19087 0.001
R27918 vp_p.n20792 vp_p.n20512 0.001
R27919 vp_p.n22216 vp_p.n21936 0.001
R27920 vp_p.n23639 vp_p.n23359 0.001
R27921 vp_p.n25061 vp_p.n24781 0.001
R27922 vp_p.n26486 vp_p.n26207 0.001
R27923 vp_p.n13963 vp_p.n13697 0.001
R27924 vp_p.n13967 vp_p.n13692 0.001
R27925 vp_p.n12297 vp_p.n11998 0.001
R27926 vp_p.n10859 vp_p.n10560 0.001
R27927 vp_p.n9422 vp_p.n9058 0.001
R27928 vp_p.n676 vp_p.n319 0.001
R27929 vp_p.n2102 vp_p.n1803 0.001
R27930 vp_p.n3527 vp_p.n3228 0.001
R27931 vp_p.n4951 vp_p.n4652 0.001
R27932 vp_p.n6374 vp_p.n6075 0.001
R27933 vp_p.n7796 vp_p.n7497 0.001
R27934 vp_p.n15100 vp_p.n14801 0.001
R27935 vp_p.n16528 vp_p.n16229 0.001
R27936 vp_p.n17955 vp_p.n17656 0.001
R27937 vp_p.n19381 vp_p.n19082 0.001
R27938 vp_p.n20806 vp_p.n20507 0.001
R27939 vp_p.n22230 vp_p.n21931 0.001
R27940 vp_p.n23653 vp_p.n23354 0.001
R27941 vp_p.n25075 vp_p.n24776 0.001
R27942 vp_p.n26500 vp_p.n26202 0.001
R27943 vp_p.n13971 vp_p.n13687 0.001
R27944 vp_p.n13975 vp_p.n13682 0.001
R27945 vp_p.n12311 vp_p.n11993 0.001
R27946 vp_p.n10873 vp_p.n10555 0.001
R27947 vp_p.n9436 vp_p.n9053 0.001
R27948 vp_p.n690 vp_p.n314 0.001
R27949 vp_p.n2116 vp_p.n1798 0.001
R27950 vp_p.n3541 vp_p.n3223 0.001
R27951 vp_p.n4965 vp_p.n4647 0.001
R27952 vp_p.n6388 vp_p.n6070 0.001
R27953 vp_p.n7810 vp_p.n7492 0.001
R27954 vp_p.n15114 vp_p.n14796 0.001
R27955 vp_p.n16542 vp_p.n16224 0.001
R27956 vp_p.n17969 vp_p.n17651 0.001
R27957 vp_p.n19395 vp_p.n19077 0.001
R27958 vp_p.n20820 vp_p.n20502 0.001
R27959 vp_p.n22244 vp_p.n21926 0.001
R27960 vp_p.n23667 vp_p.n23349 0.001
R27961 vp_p.n25089 vp_p.n24771 0.001
R27962 vp_p.n26514 vp_p.n26197 0.001
R27963 vp_p.n13979 vp_p.n13677 0.001
R27964 vp_p.n13983 vp_p.n13672 0.001
R27965 vp_p.n12325 vp_p.n11988 0.001
R27966 vp_p.n10887 vp_p.n10550 0.001
R27967 vp_p.n9450 vp_p.n9048 0.001
R27968 vp_p.n704 vp_p.n309 0.001
R27969 vp_p.n2130 vp_p.n1793 0.001
R27970 vp_p.n3555 vp_p.n3218 0.001
R27971 vp_p.n4979 vp_p.n4642 0.001
R27972 vp_p.n6402 vp_p.n6065 0.001
R27973 vp_p.n7824 vp_p.n7487 0.001
R27974 vp_p.n15128 vp_p.n14791 0.001
R27975 vp_p.n16556 vp_p.n16219 0.001
R27976 vp_p.n17983 vp_p.n17646 0.001
R27977 vp_p.n19409 vp_p.n19072 0.001
R27978 vp_p.n20834 vp_p.n20497 0.001
R27979 vp_p.n22258 vp_p.n21921 0.001
R27980 vp_p.n23681 vp_p.n23344 0.001
R27981 vp_p.n25103 vp_p.n24766 0.001
R27982 vp_p.n26528 vp_p.n26192 0.001
R27983 vp_p.n13987 vp_p.n13667 0.001
R27984 vp_p.n13991 vp_p.n13662 0.001
R27985 vp_p.n12339 vp_p.n11983 0.001
R27986 vp_p.n10901 vp_p.n10545 0.001
R27987 vp_p.n9464 vp_p.n9043 0.001
R27988 vp_p.n718 vp_p.n304 0.001
R27989 vp_p.n2144 vp_p.n1788 0.001
R27990 vp_p.n3569 vp_p.n3213 0.001
R27991 vp_p.n4993 vp_p.n4637 0.001
R27992 vp_p.n6416 vp_p.n6060 0.001
R27993 vp_p.n7838 vp_p.n7482 0.001
R27994 vp_p.n15142 vp_p.n14786 0.001
R27995 vp_p.n16570 vp_p.n16214 0.001
R27996 vp_p.n17997 vp_p.n17641 0.001
R27997 vp_p.n19423 vp_p.n19067 0.001
R27998 vp_p.n20848 vp_p.n20492 0.001
R27999 vp_p.n22272 vp_p.n21916 0.001
R28000 vp_p.n23695 vp_p.n23339 0.001
R28001 vp_p.n25117 vp_p.n24761 0.001
R28002 vp_p.n26542 vp_p.n26187 0.001
R28003 vp_p.n13995 vp_p.n13657 0.001
R28004 vp_p.n13999 vp_p.n13652 0.001
R28005 vp_p.n12353 vp_p.n11978 0.001
R28006 vp_p.n10915 vp_p.n10540 0.001
R28007 vp_p.n9478 vp_p.n9038 0.001
R28008 vp_p.n732 vp_p.n299 0.001
R28009 vp_p.n2158 vp_p.n1783 0.001
R28010 vp_p.n3583 vp_p.n3208 0.001
R28011 vp_p.n5007 vp_p.n4632 0.001
R28012 vp_p.n6430 vp_p.n6055 0.001
R28013 vp_p.n7852 vp_p.n7477 0.001
R28014 vp_p.n15156 vp_p.n14781 0.001
R28015 vp_p.n16584 vp_p.n16209 0.001
R28016 vp_p.n18011 vp_p.n17636 0.001
R28017 vp_p.n19437 vp_p.n19062 0.001
R28018 vp_p.n20862 vp_p.n20487 0.001
R28019 vp_p.n22286 vp_p.n21911 0.001
R28020 vp_p.n23709 vp_p.n23334 0.001
R28021 vp_p.n25131 vp_p.n24756 0.001
R28022 vp_p.n26556 vp_p.n26182 0.001
R28023 vp_p.n14003 vp_p.n13647 0.001
R28024 vp_p.n14007 vp_p.n13642 0.001
R28025 vp_p.n12367 vp_p.n11973 0.001
R28026 vp_p.n10929 vp_p.n10535 0.001
R28027 vp_p.n9492 vp_p.n9033 0.001
R28028 vp_p.n746 vp_p.n294 0.001
R28029 vp_p.n2172 vp_p.n1778 0.001
R28030 vp_p.n3597 vp_p.n3203 0.001
R28031 vp_p.n5021 vp_p.n4627 0.001
R28032 vp_p.n6444 vp_p.n6050 0.001
R28033 vp_p.n7866 vp_p.n7472 0.001
R28034 vp_p.n15170 vp_p.n14776 0.001
R28035 vp_p.n16598 vp_p.n16204 0.001
R28036 vp_p.n18025 vp_p.n17631 0.001
R28037 vp_p.n19451 vp_p.n19057 0.001
R28038 vp_p.n20876 vp_p.n20482 0.001
R28039 vp_p.n22300 vp_p.n21906 0.001
R28040 vp_p.n23723 vp_p.n23329 0.001
R28041 vp_p.n25145 vp_p.n24751 0.001
R28042 vp_p.n26570 vp_p.n26177 0.001
R28043 vp_p.n14011 vp_p.n13637 0.001
R28044 vp_p.n14015 vp_p.n13632 0.001
R28045 vp_p.n12381 vp_p.n11968 0.001
R28046 vp_p.n10943 vp_p.n10530 0.001
R28047 vp_p.n9506 vp_p.n9028 0.001
R28048 vp_p.n760 vp_p.n289 0.001
R28049 vp_p.n2186 vp_p.n1773 0.001
R28050 vp_p.n3611 vp_p.n3198 0.001
R28051 vp_p.n5035 vp_p.n4622 0.001
R28052 vp_p.n6458 vp_p.n6045 0.001
R28053 vp_p.n7880 vp_p.n7467 0.001
R28054 vp_p.n15184 vp_p.n14771 0.001
R28055 vp_p.n16612 vp_p.n16199 0.001
R28056 vp_p.n18039 vp_p.n17626 0.001
R28057 vp_p.n19465 vp_p.n19052 0.001
R28058 vp_p.n20890 vp_p.n20477 0.001
R28059 vp_p.n22314 vp_p.n21901 0.001
R28060 vp_p.n23737 vp_p.n23324 0.001
R28061 vp_p.n25159 vp_p.n24746 0.001
R28062 vp_p.n26584 vp_p.n26172 0.001
R28063 vp_p.n14019 vp_p.n13627 0.001
R28064 vp_p.n14023 vp_p.n13622 0.001
R28065 vp_p.n12395 vp_p.n11963 0.001
R28066 vp_p.n10957 vp_p.n10525 0.001
R28067 vp_p.n9520 vp_p.n9023 0.001
R28068 vp_p.n774 vp_p.n284 0.001
R28069 vp_p.n2200 vp_p.n1768 0.001
R28070 vp_p.n3625 vp_p.n3193 0.001
R28071 vp_p.n5049 vp_p.n4617 0.001
R28072 vp_p.n6472 vp_p.n6040 0.001
R28073 vp_p.n7894 vp_p.n7462 0.001
R28074 vp_p.n15198 vp_p.n14766 0.001
R28075 vp_p.n16626 vp_p.n16194 0.001
R28076 vp_p.n18053 vp_p.n17621 0.001
R28077 vp_p.n19479 vp_p.n19047 0.001
R28078 vp_p.n20904 vp_p.n20472 0.001
R28079 vp_p.n22328 vp_p.n21896 0.001
R28080 vp_p.n23751 vp_p.n23319 0.001
R28081 vp_p.n25173 vp_p.n24741 0.001
R28082 vp_p.n26598 vp_p.n26167 0.001
R28083 vp_p.n14027 vp_p.n13617 0.001
R28084 vp_p.n14031 vp_p.n13612 0.001
R28085 vp_p.n12409 vp_p.n11958 0.001
R28086 vp_p.n10971 vp_p.n10520 0.001
R28087 vp_p.n9534 vp_p.n9018 0.001
R28088 vp_p.n788 vp_p.n279 0.001
R28089 vp_p.n2214 vp_p.n1763 0.001
R28090 vp_p.n3639 vp_p.n3188 0.001
R28091 vp_p.n5063 vp_p.n4612 0.001
R28092 vp_p.n6486 vp_p.n6035 0.001
R28093 vp_p.n7908 vp_p.n7457 0.001
R28094 vp_p.n15212 vp_p.n14761 0.001
R28095 vp_p.n16640 vp_p.n16189 0.001
R28096 vp_p.n18067 vp_p.n17616 0.001
R28097 vp_p.n19493 vp_p.n19042 0.001
R28098 vp_p.n20918 vp_p.n20467 0.001
R28099 vp_p.n22342 vp_p.n21891 0.001
R28100 vp_p.n23765 vp_p.n23314 0.001
R28101 vp_p.n25187 vp_p.n24736 0.001
R28102 vp_p.n26612 vp_p.n26162 0.001
R28103 vp_p.n14035 vp_p.n13607 0.001
R28104 vp_p.n14039 vp_p.n13602 0.001
R28105 vp_p.n12423 vp_p.n11953 0.001
R28106 vp_p.n10985 vp_p.n10515 0.001
R28107 vp_p.n9548 vp_p.n9013 0.001
R28108 vp_p.n802 vp_p.n274 0.001
R28109 vp_p.n2228 vp_p.n1758 0.001
R28110 vp_p.n3653 vp_p.n3183 0.001
R28111 vp_p.n5077 vp_p.n4607 0.001
R28112 vp_p.n6500 vp_p.n6030 0.001
R28113 vp_p.n7922 vp_p.n7452 0.001
R28114 vp_p.n15226 vp_p.n14756 0.001
R28115 vp_p.n16654 vp_p.n16184 0.001
R28116 vp_p.n18081 vp_p.n17611 0.001
R28117 vp_p.n19507 vp_p.n19037 0.001
R28118 vp_p.n20932 vp_p.n20462 0.001
R28119 vp_p.n22356 vp_p.n21886 0.001
R28120 vp_p.n23779 vp_p.n23309 0.001
R28121 vp_p.n25201 vp_p.n24731 0.001
R28122 vp_p.n26626 vp_p.n26157 0.001
R28123 vp_p.n14043 vp_p.n13597 0.001
R28124 vp_p.n14047 vp_p.n13592 0.001
R28125 vp_p.n12437 vp_p.n11948 0.001
R28126 vp_p.n10999 vp_p.n10510 0.001
R28127 vp_p.n9562 vp_p.n9008 0.001
R28128 vp_p.n816 vp_p.n269 0.001
R28129 vp_p.n2242 vp_p.n1753 0.001
R28130 vp_p.n3667 vp_p.n3178 0.001
R28131 vp_p.n5091 vp_p.n4602 0.001
R28132 vp_p.n6514 vp_p.n6025 0.001
R28133 vp_p.n7936 vp_p.n7447 0.001
R28134 vp_p.n15240 vp_p.n14751 0.001
R28135 vp_p.n16668 vp_p.n16179 0.001
R28136 vp_p.n18095 vp_p.n17606 0.001
R28137 vp_p.n19521 vp_p.n19032 0.001
R28138 vp_p.n20946 vp_p.n20457 0.001
R28139 vp_p.n22370 vp_p.n21881 0.001
R28140 vp_p.n23793 vp_p.n23304 0.001
R28141 vp_p.n25215 vp_p.n24726 0.001
R28142 vp_p.n26640 vp_p.n26152 0.001
R28143 vp_p.n14051 vp_p.n13587 0.001
R28144 vp_p.n14055 vp_p.n13582 0.001
R28145 vp_p.n12451 vp_p.n11943 0.001
R28146 vp_p.n11013 vp_p.n10505 0.001
R28147 vp_p.n9576 vp_p.n9003 0.001
R28148 vp_p.n830 vp_p.n264 0.001
R28149 vp_p.n2256 vp_p.n1748 0.001
R28150 vp_p.n3681 vp_p.n3173 0.001
R28151 vp_p.n5105 vp_p.n4597 0.001
R28152 vp_p.n6528 vp_p.n6020 0.001
R28153 vp_p.n7950 vp_p.n7442 0.001
R28154 vp_p.n15254 vp_p.n14746 0.001
R28155 vp_p.n16682 vp_p.n16174 0.001
R28156 vp_p.n18109 vp_p.n17601 0.001
R28157 vp_p.n19535 vp_p.n19027 0.001
R28158 vp_p.n20960 vp_p.n20452 0.001
R28159 vp_p.n22384 vp_p.n21876 0.001
R28160 vp_p.n23807 vp_p.n23299 0.001
R28161 vp_p.n25229 vp_p.n24721 0.001
R28162 vp_p.n26654 vp_p.n26147 0.001
R28163 vp_p.n14059 vp_p.n13577 0.001
R28164 vp_p.n14063 vp_p.n13572 0.001
R28165 vp_p.n12465 vp_p.n11938 0.001
R28166 vp_p.n11027 vp_p.n10500 0.001
R28167 vp_p.n9590 vp_p.n8998 0.001
R28168 vp_p.n844 vp_p.n259 0.001
R28169 vp_p.n2270 vp_p.n1743 0.001
R28170 vp_p.n3695 vp_p.n3168 0.001
R28171 vp_p.n5119 vp_p.n4592 0.001
R28172 vp_p.n6542 vp_p.n6015 0.001
R28173 vp_p.n7964 vp_p.n7437 0.001
R28174 vp_p.n15268 vp_p.n14741 0.001
R28175 vp_p.n16696 vp_p.n16169 0.001
R28176 vp_p.n18123 vp_p.n17596 0.001
R28177 vp_p.n19549 vp_p.n19022 0.001
R28178 vp_p.n20974 vp_p.n20447 0.001
R28179 vp_p.n22398 vp_p.n21871 0.001
R28180 vp_p.n23821 vp_p.n23294 0.001
R28181 vp_p.n25243 vp_p.n24716 0.001
R28182 vp_p.n26668 vp_p.n26142 0.001
R28183 vp_p.n14067 vp_p.n13567 0.001
R28184 vp_p.n14071 vp_p.n13562 0.001
R28185 vp_p.n12479 vp_p.n11933 0.001
R28186 vp_p.n11041 vp_p.n10495 0.001
R28187 vp_p.n9604 vp_p.n8993 0.001
R28188 vp_p.n858 vp_p.n254 0.001
R28189 vp_p.n2284 vp_p.n1738 0.001
R28190 vp_p.n3709 vp_p.n3163 0.001
R28191 vp_p.n5133 vp_p.n4587 0.001
R28192 vp_p.n6556 vp_p.n6010 0.001
R28193 vp_p.n7978 vp_p.n7432 0.001
R28194 vp_p.n15282 vp_p.n14736 0.001
R28195 vp_p.n16710 vp_p.n16164 0.001
R28196 vp_p.n18137 vp_p.n17591 0.001
R28197 vp_p.n19563 vp_p.n19017 0.001
R28198 vp_p.n20988 vp_p.n20442 0.001
R28199 vp_p.n22412 vp_p.n21866 0.001
R28200 vp_p.n23835 vp_p.n23289 0.001
R28201 vp_p.n25257 vp_p.n24711 0.001
R28202 vp_p.n26682 vp_p.n26137 0.001
R28203 vp_p.n14075 vp_p.n13557 0.001
R28204 vp_p.n14079 vp_p.n13552 0.001
R28205 vp_p.n12493 vp_p.n11928 0.001
R28206 vp_p.n11055 vp_p.n10490 0.001
R28207 vp_p.n9618 vp_p.n8988 0.001
R28208 vp_p.n872 vp_p.n249 0.001
R28209 vp_p.n2298 vp_p.n1733 0.001
R28210 vp_p.n3723 vp_p.n3158 0.001
R28211 vp_p.n5147 vp_p.n4582 0.001
R28212 vp_p.n6570 vp_p.n6005 0.001
R28213 vp_p.n7992 vp_p.n7427 0.001
R28214 vp_p.n15296 vp_p.n14731 0.001
R28215 vp_p.n16724 vp_p.n16159 0.001
R28216 vp_p.n18151 vp_p.n17586 0.001
R28217 vp_p.n19577 vp_p.n19012 0.001
R28218 vp_p.n21002 vp_p.n20437 0.001
R28219 vp_p.n22426 vp_p.n21861 0.001
R28220 vp_p.n23849 vp_p.n23284 0.001
R28221 vp_p.n25271 vp_p.n24706 0.001
R28222 vp_p.n26696 vp_p.n26132 0.001
R28223 vp_p.n14083 vp_p.n13547 0.001
R28224 vp_p.n14087 vp_p.n13542 0.001
R28225 vp_p.n12507 vp_p.n11923 0.001
R28226 vp_p.n11069 vp_p.n10485 0.001
R28227 vp_p.n9632 vp_p.n8983 0.001
R28228 vp_p.n886 vp_p.n244 0.001
R28229 vp_p.n2312 vp_p.n1728 0.001
R28230 vp_p.n3737 vp_p.n3153 0.001
R28231 vp_p.n5161 vp_p.n4577 0.001
R28232 vp_p.n6584 vp_p.n6000 0.001
R28233 vp_p.n8006 vp_p.n7422 0.001
R28234 vp_p.n15310 vp_p.n14726 0.001
R28235 vp_p.n16738 vp_p.n16154 0.001
R28236 vp_p.n18165 vp_p.n17581 0.001
R28237 vp_p.n19591 vp_p.n19007 0.001
R28238 vp_p.n21016 vp_p.n20432 0.001
R28239 vp_p.n22440 vp_p.n21856 0.001
R28240 vp_p.n23863 vp_p.n23279 0.001
R28241 vp_p.n25285 vp_p.n24701 0.001
R28242 vp_p.n26710 vp_p.n26127 0.001
R28243 vp_p.n14091 vp_p.n13537 0.001
R28244 vp_p.n14095 vp_p.n13532 0.001
R28245 vp_p.n12521 vp_p.n11918 0.001
R28246 vp_p.n11083 vp_p.n10480 0.001
R28247 vp_p.n9646 vp_p.n8978 0.001
R28248 vp_p.n900 vp_p.n239 0.001
R28249 vp_p.n2326 vp_p.n1723 0.001
R28250 vp_p.n3751 vp_p.n3148 0.001
R28251 vp_p.n5175 vp_p.n4572 0.001
R28252 vp_p.n6598 vp_p.n5995 0.001
R28253 vp_p.n8020 vp_p.n7417 0.001
R28254 vp_p.n15324 vp_p.n14721 0.001
R28255 vp_p.n16752 vp_p.n16149 0.001
R28256 vp_p.n18179 vp_p.n17576 0.001
R28257 vp_p.n19605 vp_p.n19002 0.001
R28258 vp_p.n21030 vp_p.n20427 0.001
R28259 vp_p.n22454 vp_p.n21851 0.001
R28260 vp_p.n23877 vp_p.n23274 0.001
R28261 vp_p.n25299 vp_p.n24696 0.001
R28262 vp_p.n26724 vp_p.n26122 0.001
R28263 vp_p.n14099 vp_p.n13527 0.001
R28264 vp_p.n14103 vp_p.n13522 0.001
R28265 vp_p.n12535 vp_p.n11913 0.001
R28266 vp_p.n11097 vp_p.n10475 0.001
R28267 vp_p.n9660 vp_p.n8973 0.001
R28268 vp_p.n914 vp_p.n234 0.001
R28269 vp_p.n2340 vp_p.n1718 0.001
R28270 vp_p.n3765 vp_p.n3143 0.001
R28271 vp_p.n5189 vp_p.n4567 0.001
R28272 vp_p.n6612 vp_p.n5990 0.001
R28273 vp_p.n8034 vp_p.n7412 0.001
R28274 vp_p.n15338 vp_p.n14716 0.001
R28275 vp_p.n16766 vp_p.n16144 0.001
R28276 vp_p.n18193 vp_p.n17571 0.001
R28277 vp_p.n19619 vp_p.n18997 0.001
R28278 vp_p.n21044 vp_p.n20422 0.001
R28279 vp_p.n22468 vp_p.n21846 0.001
R28280 vp_p.n23891 vp_p.n23269 0.001
R28281 vp_p.n25313 vp_p.n24691 0.001
R28282 vp_p.n26738 vp_p.n26117 0.001
R28283 vp_p.n14107 vp_p.n13517 0.001
R28284 vp_p.n14111 vp_p.n13512 0.001
R28285 vp_p.n12549 vp_p.n11908 0.001
R28286 vp_p.n11111 vp_p.n10470 0.001
R28287 vp_p.n9674 vp_p.n8968 0.001
R28288 vp_p.n928 vp_p.n229 0.001
R28289 vp_p.n2354 vp_p.n1713 0.001
R28290 vp_p.n3779 vp_p.n3138 0.001
R28291 vp_p.n5203 vp_p.n4562 0.001
R28292 vp_p.n6626 vp_p.n5985 0.001
R28293 vp_p.n8048 vp_p.n7407 0.001
R28294 vp_p.n15352 vp_p.n14711 0.001
R28295 vp_p.n16780 vp_p.n16139 0.001
R28296 vp_p.n18207 vp_p.n17566 0.001
R28297 vp_p.n19633 vp_p.n18992 0.001
R28298 vp_p.n21058 vp_p.n20417 0.001
R28299 vp_p.n22482 vp_p.n21841 0.001
R28300 vp_p.n23905 vp_p.n23264 0.001
R28301 vp_p.n25327 vp_p.n24686 0.001
R28302 vp_p.n26752 vp_p.n26112 0.001
R28303 vp_p.n14115 vp_p.n13507 0.001
R28304 vp_p.n14119 vp_p.n13502 0.001
R28305 vp_p.n12563 vp_p.n11903 0.001
R28306 vp_p.n11125 vp_p.n10465 0.001
R28307 vp_p.n9688 vp_p.n8963 0.001
R28308 vp_p.n942 vp_p.n224 0.001
R28309 vp_p.n2368 vp_p.n1708 0.001
R28310 vp_p.n3793 vp_p.n3133 0.001
R28311 vp_p.n5217 vp_p.n4557 0.001
R28312 vp_p.n6640 vp_p.n5980 0.001
R28313 vp_p.n8062 vp_p.n7402 0.001
R28314 vp_p.n15366 vp_p.n14706 0.001
R28315 vp_p.n16794 vp_p.n16134 0.001
R28316 vp_p.n18221 vp_p.n17561 0.001
R28317 vp_p.n19647 vp_p.n18987 0.001
R28318 vp_p.n21072 vp_p.n20412 0.001
R28319 vp_p.n22496 vp_p.n21836 0.001
R28320 vp_p.n23919 vp_p.n23259 0.001
R28321 vp_p.n25341 vp_p.n24681 0.001
R28322 vp_p.n26766 vp_p.n26107 0.001
R28323 vp_p.n14123 vp_p.n13497 0.001
R28324 vp_p.n14127 vp_p.n13492 0.001
R28325 vp_p.n12577 vp_p.n11898 0.001
R28326 vp_p.n11139 vp_p.n10460 0.001
R28327 vp_p.n9702 vp_p.n8958 0.001
R28328 vp_p.n956 vp_p.n219 0.001
R28329 vp_p.n2382 vp_p.n1703 0.001
R28330 vp_p.n3807 vp_p.n3128 0.001
R28331 vp_p.n5231 vp_p.n4552 0.001
R28332 vp_p.n6654 vp_p.n5975 0.001
R28333 vp_p.n8076 vp_p.n7397 0.001
R28334 vp_p.n15380 vp_p.n14701 0.001
R28335 vp_p.n16808 vp_p.n16129 0.001
R28336 vp_p.n18235 vp_p.n17556 0.001
R28337 vp_p.n19661 vp_p.n18982 0.001
R28338 vp_p.n21086 vp_p.n20407 0.001
R28339 vp_p.n22510 vp_p.n21831 0.001
R28340 vp_p.n23933 vp_p.n23254 0.001
R28341 vp_p.n25355 vp_p.n24676 0.001
R28342 vp_p.n26780 vp_p.n26102 0.001
R28343 vp_p.n14131 vp_p.n13487 0.001
R28344 vp_p.n14135 vp_p.n13482 0.001
R28345 vp_p.n12591 vp_p.n11893 0.001
R28346 vp_p.n11153 vp_p.n10455 0.001
R28347 vp_p.n9716 vp_p.n8953 0.001
R28348 vp_p.n970 vp_p.n214 0.001
R28349 vp_p.n2396 vp_p.n1698 0.001
R28350 vp_p.n3821 vp_p.n3123 0.001
R28351 vp_p.n5245 vp_p.n4547 0.001
R28352 vp_p.n6668 vp_p.n5970 0.001
R28353 vp_p.n8090 vp_p.n7392 0.001
R28354 vp_p.n15394 vp_p.n14696 0.001
R28355 vp_p.n16822 vp_p.n16124 0.001
R28356 vp_p.n18249 vp_p.n17551 0.001
R28357 vp_p.n19675 vp_p.n18977 0.001
R28358 vp_p.n21100 vp_p.n20402 0.001
R28359 vp_p.n22524 vp_p.n21826 0.001
R28360 vp_p.n23947 vp_p.n23249 0.001
R28361 vp_p.n25369 vp_p.n24671 0.001
R28362 vp_p.n26794 vp_p.n26097 0.001
R28363 vp_p.n14139 vp_p.n13477 0.001
R28364 vp_p.n14143 vp_p.n13472 0.001
R28365 vp_p.n12605 vp_p.n11888 0.001
R28366 vp_p.n11167 vp_p.n10450 0.001
R28367 vp_p.n9730 vp_p.n8948 0.001
R28368 vp_p.n984 vp_p.n209 0.001
R28369 vp_p.n2410 vp_p.n1693 0.001
R28370 vp_p.n3835 vp_p.n3118 0.001
R28371 vp_p.n5259 vp_p.n4542 0.001
R28372 vp_p.n6682 vp_p.n5965 0.001
R28373 vp_p.n8104 vp_p.n7387 0.001
R28374 vp_p.n15408 vp_p.n14691 0.001
R28375 vp_p.n16836 vp_p.n16119 0.001
R28376 vp_p.n18263 vp_p.n17546 0.001
R28377 vp_p.n19689 vp_p.n18972 0.001
R28378 vp_p.n21114 vp_p.n20397 0.001
R28379 vp_p.n22538 vp_p.n21821 0.001
R28380 vp_p.n23961 vp_p.n23244 0.001
R28381 vp_p.n25383 vp_p.n24666 0.001
R28382 vp_p.n26808 vp_p.n26092 0.001
R28383 vp_p.n14147 vp_p.n13467 0.001
R28384 vp_p.n14151 vp_p.n13462 0.001
R28385 vp_p.n12619 vp_p.n11883 0.001
R28386 vp_p.n11181 vp_p.n10445 0.001
R28387 vp_p.n9744 vp_p.n8943 0.001
R28388 vp_p.n998 vp_p.n204 0.001
R28389 vp_p.n2424 vp_p.n1688 0.001
R28390 vp_p.n3849 vp_p.n3113 0.001
R28391 vp_p.n5273 vp_p.n4537 0.001
R28392 vp_p.n6696 vp_p.n5960 0.001
R28393 vp_p.n8118 vp_p.n7382 0.001
R28394 vp_p.n15422 vp_p.n14686 0.001
R28395 vp_p.n16850 vp_p.n16114 0.001
R28396 vp_p.n18277 vp_p.n17541 0.001
R28397 vp_p.n19703 vp_p.n18967 0.001
R28398 vp_p.n21128 vp_p.n20392 0.001
R28399 vp_p.n22552 vp_p.n21816 0.001
R28400 vp_p.n23975 vp_p.n23239 0.001
R28401 vp_p.n25397 vp_p.n24661 0.001
R28402 vp_p.n26822 vp_p.n26087 0.001
R28403 vp_p.n14155 vp_p.n13457 0.001
R28404 vp_p.n14159 vp_p.n13452 0.001
R28405 vp_p.n12633 vp_p.n11878 0.001
R28406 vp_p.n11195 vp_p.n10440 0.001
R28407 vp_p.n9758 vp_p.n8938 0.001
R28408 vp_p.n1012 vp_p.n199 0.001
R28409 vp_p.n2438 vp_p.n1683 0.001
R28410 vp_p.n3863 vp_p.n3108 0.001
R28411 vp_p.n5287 vp_p.n4532 0.001
R28412 vp_p.n6710 vp_p.n5955 0.001
R28413 vp_p.n8132 vp_p.n7377 0.001
R28414 vp_p.n15436 vp_p.n14681 0.001
R28415 vp_p.n16864 vp_p.n16109 0.001
R28416 vp_p.n18291 vp_p.n17536 0.001
R28417 vp_p.n19717 vp_p.n18962 0.001
R28418 vp_p.n21142 vp_p.n20387 0.001
R28419 vp_p.n22566 vp_p.n21811 0.001
R28420 vp_p.n23989 vp_p.n23234 0.001
R28421 vp_p.n25411 vp_p.n24656 0.001
R28422 vp_p.n26836 vp_p.n26082 0.001
R28423 vp_p.n14163 vp_p.n13447 0.001
R28424 vp_p.n14167 vp_p.n13442 0.001
R28425 vp_p.n12647 vp_p.n11873 0.001
R28426 vp_p.n11209 vp_p.n10435 0.001
R28427 vp_p.n9772 vp_p.n8933 0.001
R28428 vp_p.n1026 vp_p.n194 0.001
R28429 vp_p.n2452 vp_p.n1678 0.001
R28430 vp_p.n3877 vp_p.n3103 0.001
R28431 vp_p.n5301 vp_p.n4527 0.001
R28432 vp_p.n6724 vp_p.n5950 0.001
R28433 vp_p.n8146 vp_p.n7372 0.001
R28434 vp_p.n15450 vp_p.n14676 0.001
R28435 vp_p.n16878 vp_p.n16104 0.001
R28436 vp_p.n18305 vp_p.n17531 0.001
R28437 vp_p.n19731 vp_p.n18957 0.001
R28438 vp_p.n21156 vp_p.n20382 0.001
R28439 vp_p.n22580 vp_p.n21806 0.001
R28440 vp_p.n24003 vp_p.n23229 0.001
R28441 vp_p.n25425 vp_p.n24651 0.001
R28442 vp_p.n26850 vp_p.n26077 0.001
R28443 vp_p.n14171 vp_p.n13437 0.001
R28444 vp_p.n14175 vp_p.n13432 0.001
R28445 vp_p.n12661 vp_p.n11868 0.001
R28446 vp_p.n11223 vp_p.n10430 0.001
R28447 vp_p.n9786 vp_p.n8928 0.001
R28448 vp_p.n1040 vp_p.n189 0.001
R28449 vp_p.n2466 vp_p.n1673 0.001
R28450 vp_p.n3891 vp_p.n3098 0.001
R28451 vp_p.n5315 vp_p.n4522 0.001
R28452 vp_p.n6738 vp_p.n5945 0.001
R28453 vp_p.n8160 vp_p.n7367 0.001
R28454 vp_p.n15464 vp_p.n14671 0.001
R28455 vp_p.n16892 vp_p.n16099 0.001
R28456 vp_p.n18319 vp_p.n17526 0.001
R28457 vp_p.n19745 vp_p.n18952 0.001
R28458 vp_p.n21170 vp_p.n20377 0.001
R28459 vp_p.n22594 vp_p.n21801 0.001
R28460 vp_p.n24017 vp_p.n23224 0.001
R28461 vp_p.n25439 vp_p.n24646 0.001
R28462 vp_p.n26864 vp_p.n26072 0.001
R28463 vp_p.n14179 vp_p.n13427 0.001
R28464 vp_p.n14183 vp_p.n13422 0.001
R28465 vp_p.n12675 vp_p.n11863 0.001
R28466 vp_p.n11237 vp_p.n10425 0.001
R28467 vp_p.n9800 vp_p.n8923 0.001
R28468 vp_p.n1054 vp_p.n184 0.001
R28469 vp_p.n2480 vp_p.n1668 0.001
R28470 vp_p.n3905 vp_p.n3093 0.001
R28471 vp_p.n5329 vp_p.n4517 0.001
R28472 vp_p.n6752 vp_p.n5940 0.001
R28473 vp_p.n8174 vp_p.n7362 0.001
R28474 vp_p.n15478 vp_p.n14666 0.001
R28475 vp_p.n16906 vp_p.n16094 0.001
R28476 vp_p.n18333 vp_p.n17521 0.001
R28477 vp_p.n19759 vp_p.n18947 0.001
R28478 vp_p.n21184 vp_p.n20372 0.001
R28479 vp_p.n22608 vp_p.n21796 0.001
R28480 vp_p.n24031 vp_p.n23219 0.001
R28481 vp_p.n25453 vp_p.n24641 0.001
R28482 vp_p.n26878 vp_p.n26067 0.001
R28483 vp_p.n14187 vp_p.n13417 0.001
R28484 vp_p.n14191 vp_p.n13412 0.001
R28485 vp_p.n12689 vp_p.n11858 0.001
R28486 vp_p.n11251 vp_p.n10420 0.001
R28487 vp_p.n9814 vp_p.n8918 0.001
R28488 vp_p.n1068 vp_p.n179 0.001
R28489 vp_p.n2494 vp_p.n1663 0.001
R28490 vp_p.n3919 vp_p.n3088 0.001
R28491 vp_p.n5343 vp_p.n4512 0.001
R28492 vp_p.n6766 vp_p.n5935 0.001
R28493 vp_p.n8188 vp_p.n7357 0.001
R28494 vp_p.n15492 vp_p.n14661 0.001
R28495 vp_p.n16920 vp_p.n16089 0.001
R28496 vp_p.n18347 vp_p.n17516 0.001
R28497 vp_p.n19773 vp_p.n18942 0.001
R28498 vp_p.n21198 vp_p.n20367 0.001
R28499 vp_p.n22622 vp_p.n21791 0.001
R28500 vp_p.n24045 vp_p.n23214 0.001
R28501 vp_p.n25467 vp_p.n24636 0.001
R28502 vp_p.n26892 vp_p.n26062 0.001
R28503 vp_p.n14195 vp_p.n13407 0.001
R28504 vp_p.n14199 vp_p.n13402 0.001
R28505 vp_p.n12703 vp_p.n11853 0.001
R28506 vp_p.n11265 vp_p.n10415 0.001
R28507 vp_p.n9828 vp_p.n8913 0.001
R28508 vp_p.n1082 vp_p.n174 0.001
R28509 vp_p.n2508 vp_p.n1658 0.001
R28510 vp_p.n3933 vp_p.n3083 0.001
R28511 vp_p.n5357 vp_p.n4507 0.001
R28512 vp_p.n6780 vp_p.n5930 0.001
R28513 vp_p.n8202 vp_p.n7352 0.001
R28514 vp_p.n15506 vp_p.n14656 0.001
R28515 vp_p.n16934 vp_p.n16084 0.001
R28516 vp_p.n18361 vp_p.n17511 0.001
R28517 vp_p.n19787 vp_p.n18937 0.001
R28518 vp_p.n21212 vp_p.n20362 0.001
R28519 vp_p.n22636 vp_p.n21786 0.001
R28520 vp_p.n24059 vp_p.n23209 0.001
R28521 vp_p.n25481 vp_p.n24631 0.001
R28522 vp_p.n26906 vp_p.n26057 0.001
R28523 vp_p.n14203 vp_p.n13397 0.001
R28524 vp_p.n14207 vp_p.n13392 0.001
R28525 vp_p.n12717 vp_p.n11848 0.001
R28526 vp_p.n11279 vp_p.n10410 0.001
R28527 vp_p.n9842 vp_p.n8908 0.001
R28528 vp_p.n1096 vp_p.n169 0.001
R28529 vp_p.n2522 vp_p.n1653 0.001
R28530 vp_p.n3947 vp_p.n3078 0.001
R28531 vp_p.n5371 vp_p.n4502 0.001
R28532 vp_p.n6794 vp_p.n5925 0.001
R28533 vp_p.n8216 vp_p.n7347 0.001
R28534 vp_p.n15520 vp_p.n14651 0.001
R28535 vp_p.n16948 vp_p.n16079 0.001
R28536 vp_p.n18375 vp_p.n17506 0.001
R28537 vp_p.n19801 vp_p.n18932 0.001
R28538 vp_p.n21226 vp_p.n20357 0.001
R28539 vp_p.n22650 vp_p.n21781 0.001
R28540 vp_p.n24073 vp_p.n23204 0.001
R28541 vp_p.n25495 vp_p.n24626 0.001
R28542 vp_p.n26920 vp_p.n26052 0.001
R28543 vp_p.n14211 vp_p.n13387 0.001
R28544 vp_p.n14215 vp_p.n13382 0.001
R28545 vp_p.n12731 vp_p.n11843 0.001
R28546 vp_p.n11293 vp_p.n10405 0.001
R28547 vp_p.n9856 vp_p.n8903 0.001
R28548 vp_p.n1110 vp_p.n164 0.001
R28549 vp_p.n2536 vp_p.n1648 0.001
R28550 vp_p.n3961 vp_p.n3073 0.001
R28551 vp_p.n5385 vp_p.n4497 0.001
R28552 vp_p.n6808 vp_p.n5920 0.001
R28553 vp_p.n8230 vp_p.n7342 0.001
R28554 vp_p.n15534 vp_p.n14646 0.001
R28555 vp_p.n16962 vp_p.n16074 0.001
R28556 vp_p.n18389 vp_p.n17501 0.001
R28557 vp_p.n19815 vp_p.n18927 0.001
R28558 vp_p.n21240 vp_p.n20352 0.001
R28559 vp_p.n22664 vp_p.n21776 0.001
R28560 vp_p.n24087 vp_p.n23199 0.001
R28561 vp_p.n25509 vp_p.n24621 0.001
R28562 vp_p.n26934 vp_p.n26047 0.001
R28563 vp_p.n14219 vp_p.n13377 0.001
R28564 vp_p.n14223 vp_p.n13372 0.001
R28565 vp_p.n12745 vp_p.n11838 0.001
R28566 vp_p.n11307 vp_p.n10400 0.001
R28567 vp_p.n9870 vp_p.n8898 0.001
R28568 vp_p.n1124 vp_p.n159 0.001
R28569 vp_p.n2550 vp_p.n1643 0.001
R28570 vp_p.n3975 vp_p.n3068 0.001
R28571 vp_p.n5399 vp_p.n4492 0.001
R28572 vp_p.n6822 vp_p.n5915 0.001
R28573 vp_p.n8244 vp_p.n7337 0.001
R28574 vp_p.n15548 vp_p.n14641 0.001
R28575 vp_p.n16976 vp_p.n16069 0.001
R28576 vp_p.n18403 vp_p.n17496 0.001
R28577 vp_p.n19829 vp_p.n18922 0.001
R28578 vp_p.n21254 vp_p.n20347 0.001
R28579 vp_p.n22678 vp_p.n21771 0.001
R28580 vp_p.n24101 vp_p.n23194 0.001
R28581 vp_p.n25523 vp_p.n24616 0.001
R28582 vp_p.n26948 vp_p.n26042 0.001
R28583 vp_p.n14227 vp_p.n13367 0.001
R28584 vp_p.n14231 vp_p.n13362 0.001
R28585 vp_p.n12759 vp_p.n11833 0.001
R28586 vp_p.n11321 vp_p.n10395 0.001
R28587 vp_p.n9884 vp_p.n8893 0.001
R28588 vp_p.n1138 vp_p.n154 0.001
R28589 vp_p.n2564 vp_p.n1638 0.001
R28590 vp_p.n3989 vp_p.n3063 0.001
R28591 vp_p.n5413 vp_p.n4487 0.001
R28592 vp_p.n6836 vp_p.n5910 0.001
R28593 vp_p.n8258 vp_p.n7332 0.001
R28594 vp_p.n15562 vp_p.n14636 0.001
R28595 vp_p.n16990 vp_p.n16064 0.001
R28596 vp_p.n18417 vp_p.n17491 0.001
R28597 vp_p.n19843 vp_p.n18917 0.001
R28598 vp_p.n21268 vp_p.n20342 0.001
R28599 vp_p.n22692 vp_p.n21766 0.001
R28600 vp_p.n24115 vp_p.n23189 0.001
R28601 vp_p.n25537 vp_p.n24611 0.001
R28602 vp_p.n26962 vp_p.n26037 0.001
R28603 vp_p.n14235 vp_p.n13357 0.001
R28604 vp_p.n14239 vp_p.n13352 0.001
R28605 vp_p.n12773 vp_p.n11828 0.001
R28606 vp_p.n11335 vp_p.n10390 0.001
R28607 vp_p.n9898 vp_p.n8888 0.001
R28608 vp_p.n1152 vp_p.n149 0.001
R28609 vp_p.n2578 vp_p.n1633 0.001
R28610 vp_p.n4003 vp_p.n3058 0.001
R28611 vp_p.n5427 vp_p.n4482 0.001
R28612 vp_p.n6850 vp_p.n5905 0.001
R28613 vp_p.n8272 vp_p.n7327 0.001
R28614 vp_p.n15576 vp_p.n14631 0.001
R28615 vp_p.n17004 vp_p.n16059 0.001
R28616 vp_p.n18431 vp_p.n17486 0.001
R28617 vp_p.n19857 vp_p.n18912 0.001
R28618 vp_p.n21282 vp_p.n20337 0.001
R28619 vp_p.n22706 vp_p.n21761 0.001
R28620 vp_p.n24129 vp_p.n23184 0.001
R28621 vp_p.n25551 vp_p.n24606 0.001
R28622 vp_p.n26976 vp_p.n26032 0.001
R28623 vp_p.n14243 vp_p.n13347 0.001
R28624 vp_p.n14247 vp_p.n13342 0.001
R28625 vp_p.n12787 vp_p.n11823 0.001
R28626 vp_p.n11349 vp_p.n10385 0.001
R28627 vp_p.n9912 vp_p.n8883 0.001
R28628 vp_p.n1166 vp_p.n144 0.001
R28629 vp_p.n2592 vp_p.n1628 0.001
R28630 vp_p.n4017 vp_p.n3053 0.001
R28631 vp_p.n5441 vp_p.n4477 0.001
R28632 vp_p.n6864 vp_p.n5900 0.001
R28633 vp_p.n8286 vp_p.n7322 0.001
R28634 vp_p.n15590 vp_p.n14626 0.001
R28635 vp_p.n17018 vp_p.n16054 0.001
R28636 vp_p.n18445 vp_p.n17481 0.001
R28637 vp_p.n19871 vp_p.n18907 0.001
R28638 vp_p.n21296 vp_p.n20332 0.001
R28639 vp_p.n22720 vp_p.n21756 0.001
R28640 vp_p.n24143 vp_p.n23179 0.001
R28641 vp_p.n25565 vp_p.n24601 0.001
R28642 vp_p.n26990 vp_p.n26027 0.001
R28643 vp_p.n14251 vp_p.n13337 0.001
R28644 vp_p.n14255 vp_p.n13332 0.001
R28645 vp_p.n12801 vp_p.n11818 0.001
R28646 vp_p.n11363 vp_p.n10380 0.001
R28647 vp_p.n9926 vp_p.n8878 0.001
R28648 vp_p.n1180 vp_p.n139 0.001
R28649 vp_p.n2606 vp_p.n1623 0.001
R28650 vp_p.n4031 vp_p.n3048 0.001
R28651 vp_p.n5455 vp_p.n4472 0.001
R28652 vp_p.n6878 vp_p.n5895 0.001
R28653 vp_p.n8300 vp_p.n7317 0.001
R28654 vp_p.n15604 vp_p.n14621 0.001
R28655 vp_p.n17032 vp_p.n16049 0.001
R28656 vp_p.n18459 vp_p.n17476 0.001
R28657 vp_p.n19885 vp_p.n18902 0.001
R28658 vp_p.n21310 vp_p.n20327 0.001
R28659 vp_p.n22734 vp_p.n21751 0.001
R28660 vp_p.n24157 vp_p.n23174 0.001
R28661 vp_p.n25579 vp_p.n24596 0.001
R28662 vp_p.n27004 vp_p.n26022 0.001
R28663 vp_p.n14259 vp_p.n13327 0.001
R28664 vp_p.n14263 vp_p.n13322 0.001
R28665 vp_p.n12815 vp_p.n11813 0.001
R28666 vp_p.n11377 vp_p.n10375 0.001
R28667 vp_p.n9940 vp_p.n8873 0.001
R28668 vp_p.n1194 vp_p.n134 0.001
R28669 vp_p.n2620 vp_p.n1618 0.001
R28670 vp_p.n4045 vp_p.n3043 0.001
R28671 vp_p.n5469 vp_p.n4467 0.001
R28672 vp_p.n6892 vp_p.n5890 0.001
R28673 vp_p.n8314 vp_p.n7312 0.001
R28674 vp_p.n15618 vp_p.n14616 0.001
R28675 vp_p.n17046 vp_p.n16044 0.001
R28676 vp_p.n18473 vp_p.n17471 0.001
R28677 vp_p.n19899 vp_p.n18897 0.001
R28678 vp_p.n21324 vp_p.n20322 0.001
R28679 vp_p.n22748 vp_p.n21746 0.001
R28680 vp_p.n24171 vp_p.n23169 0.001
R28681 vp_p.n25593 vp_p.n24591 0.001
R28682 vp_p.n27018 vp_p.n26017 0.001
R28683 vp_p.n14267 vp_p.n13317 0.001
R28684 vp_p.n14271 vp_p.n13312 0.001
R28685 vp_p.n12829 vp_p.n11808 0.001
R28686 vp_p.n11391 vp_p.n10370 0.001
R28687 vp_p.n9954 vp_p.n8868 0.001
R28688 vp_p.n1208 vp_p.n129 0.001
R28689 vp_p.n2634 vp_p.n1613 0.001
R28690 vp_p.n4059 vp_p.n3038 0.001
R28691 vp_p.n5483 vp_p.n4462 0.001
R28692 vp_p.n6906 vp_p.n5885 0.001
R28693 vp_p.n8328 vp_p.n7307 0.001
R28694 vp_p.n15632 vp_p.n14611 0.001
R28695 vp_p.n17060 vp_p.n16039 0.001
R28696 vp_p.n18487 vp_p.n17466 0.001
R28697 vp_p.n19913 vp_p.n18892 0.001
R28698 vp_p.n21338 vp_p.n20317 0.001
R28699 vp_p.n22762 vp_p.n21741 0.001
R28700 vp_p.n24185 vp_p.n23164 0.001
R28701 vp_p.n25607 vp_p.n24586 0.001
R28702 vp_p.n27032 vp_p.n26012 0.001
R28703 vp_p.n14275 vp_p.n13307 0.001
R28704 vp_p.n14279 vp_p.n13302 0.001
R28705 vp_p.n12843 vp_p.n11803 0.001
R28706 vp_p.n11405 vp_p.n10365 0.001
R28707 vp_p.n9968 vp_p.n8863 0.001
R28708 vp_p.n1222 vp_p.n124 0.001
R28709 vp_p.n2648 vp_p.n1608 0.001
R28710 vp_p.n4073 vp_p.n3033 0.001
R28711 vp_p.n5497 vp_p.n4457 0.001
R28712 vp_p.n6920 vp_p.n5880 0.001
R28713 vp_p.n8342 vp_p.n7302 0.001
R28714 vp_p.n15646 vp_p.n14606 0.001
R28715 vp_p.n17074 vp_p.n16034 0.001
R28716 vp_p.n18501 vp_p.n17461 0.001
R28717 vp_p.n19927 vp_p.n18887 0.001
R28718 vp_p.n21352 vp_p.n20312 0.001
R28719 vp_p.n22776 vp_p.n21736 0.001
R28720 vp_p.n24199 vp_p.n23159 0.001
R28721 vp_p.n25621 vp_p.n24581 0.001
R28722 vp_p.n27046 vp_p.n26007 0.001
R28723 vp_p.n14283 vp_p.n13297 0.001
R28724 vp_p.n14287 vp_p.n13292 0.001
R28725 vp_p.n12857 vp_p.n11798 0.001
R28726 vp_p.n11419 vp_p.n10360 0.001
R28727 vp_p.n9982 vp_p.n8858 0.001
R28728 vp_p.n1236 vp_p.n119 0.001
R28729 vp_p.n2662 vp_p.n1603 0.001
R28730 vp_p.n4087 vp_p.n3028 0.001
R28731 vp_p.n5511 vp_p.n4452 0.001
R28732 vp_p.n6934 vp_p.n5875 0.001
R28733 vp_p.n8356 vp_p.n7297 0.001
R28734 vp_p.n15660 vp_p.n14601 0.001
R28735 vp_p.n17088 vp_p.n16029 0.001
R28736 vp_p.n18515 vp_p.n17456 0.001
R28737 vp_p.n19941 vp_p.n18882 0.001
R28738 vp_p.n21366 vp_p.n20307 0.001
R28739 vp_p.n22790 vp_p.n21731 0.001
R28740 vp_p.n24213 vp_p.n23154 0.001
R28741 vp_p.n25635 vp_p.n24576 0.001
R28742 vp_p.n27060 vp_p.n26002 0.001
R28743 vp_p.n14291 vp_p.n13287 0.001
R28744 vp_p.n14295 vp_p.n13282 0.001
R28745 vp_p.n12871 vp_p.n11793 0.001
R28746 vp_p.n11433 vp_p.n10355 0.001
R28747 vp_p.n9996 vp_p.n8853 0.001
R28748 vp_p.n1250 vp_p.n114 0.001
R28749 vp_p.n2676 vp_p.n1598 0.001
R28750 vp_p.n4101 vp_p.n3023 0.001
R28751 vp_p.n5525 vp_p.n4447 0.001
R28752 vp_p.n6948 vp_p.n5870 0.001
R28753 vp_p.n8370 vp_p.n7292 0.001
R28754 vp_p.n15674 vp_p.n14596 0.001
R28755 vp_p.n17102 vp_p.n16024 0.001
R28756 vp_p.n18529 vp_p.n17451 0.001
R28757 vp_p.n19955 vp_p.n18877 0.001
R28758 vp_p.n21380 vp_p.n20302 0.001
R28759 vp_p.n22804 vp_p.n21726 0.001
R28760 vp_p.n24227 vp_p.n23149 0.001
R28761 vp_p.n25649 vp_p.n24571 0.001
R28762 vp_p.n27074 vp_p.n25997 0.001
R28763 vp_p.n14299 vp_p.n13277 0.001
R28764 vp_p.n14303 vp_p.n13272 0.001
R28765 vp_p.n12885 vp_p.n11788 0.001
R28766 vp_p.n11447 vp_p.n10350 0.001
R28767 vp_p.n10010 vp_p.n8848 0.001
R28768 vp_p.n1264 vp_p.n109 0.001
R28769 vp_p.n2690 vp_p.n1593 0.001
R28770 vp_p.n4115 vp_p.n3018 0.001
R28771 vp_p.n5539 vp_p.n4442 0.001
R28772 vp_p.n6962 vp_p.n5865 0.001
R28773 vp_p.n8384 vp_p.n7287 0.001
R28774 vp_p.n15688 vp_p.n14591 0.001
R28775 vp_p.n17116 vp_p.n16019 0.001
R28776 vp_p.n18543 vp_p.n17446 0.001
R28777 vp_p.n19969 vp_p.n18872 0.001
R28778 vp_p.n21394 vp_p.n20297 0.001
R28779 vp_p.n22818 vp_p.n21721 0.001
R28780 vp_p.n24241 vp_p.n23144 0.001
R28781 vp_p.n25663 vp_p.n24566 0.001
R28782 vp_p.n27088 vp_p.n25992 0.001
R28783 vp_p.n14307 vp_p.n13267 0.001
R28784 vp_p.n14311 vp_p.n13262 0.001
R28785 vp_p.n12899 vp_p.n11783 0.001
R28786 vp_p.n11461 vp_p.n10345 0.001
R28787 vp_p.n10024 vp_p.n8843 0.001
R28788 vp_p.n1278 vp_p.n104 0.001
R28789 vp_p.n2704 vp_p.n1588 0.001
R28790 vp_p.n4129 vp_p.n3013 0.001
R28791 vp_p.n5553 vp_p.n4437 0.001
R28792 vp_p.n6976 vp_p.n5860 0.001
R28793 vp_p.n8398 vp_p.n7282 0.001
R28794 vp_p.n15702 vp_p.n14586 0.001
R28795 vp_p.n17130 vp_p.n16014 0.001
R28796 vp_p.n18557 vp_p.n17441 0.001
R28797 vp_p.n19983 vp_p.n18867 0.001
R28798 vp_p.n21408 vp_p.n20292 0.001
R28799 vp_p.n22832 vp_p.n21716 0.001
R28800 vp_p.n24255 vp_p.n23139 0.001
R28801 vp_p.n25677 vp_p.n24561 0.001
R28802 vp_p.n27102 vp_p.n25987 0.001
R28803 vp_p.n14315 vp_p.n13257 0.001
R28804 vp_p.n14319 vp_p.n13252 0.001
R28805 vp_p.n12913 vp_p.n11778 0.001
R28806 vp_p.n11475 vp_p.n10340 0.001
R28807 vp_p.n10038 vp_p.n8838 0.001
R28808 vp_p.n1292 vp_p.n99 0.001
R28809 vp_p.n2718 vp_p.n1583 0.001
R28810 vp_p.n4143 vp_p.n3008 0.001
R28811 vp_p.n5567 vp_p.n4432 0.001
R28812 vp_p.n6990 vp_p.n5855 0.001
R28813 vp_p.n8412 vp_p.n7277 0.001
R28814 vp_p.n15716 vp_p.n14581 0.001
R28815 vp_p.n17144 vp_p.n16009 0.001
R28816 vp_p.n18571 vp_p.n17436 0.001
R28817 vp_p.n19997 vp_p.n18862 0.001
R28818 vp_p.n21422 vp_p.n20287 0.001
R28819 vp_p.n22846 vp_p.n21711 0.001
R28820 vp_p.n24269 vp_p.n23134 0.001
R28821 vp_p.n25691 vp_p.n24556 0.001
R28822 vp_p.n27116 vp_p.n25982 0.001
R28823 vp_p.n14323 vp_p.n13247 0.001
R28824 vp_p.n14327 vp_p.n13242 0.001
R28825 vp_p.n12927 vp_p.n11773 0.001
R28826 vp_p.n11489 vp_p.n10335 0.001
R28827 vp_p.n10052 vp_p.n8833 0.001
R28828 vp_p.n1306 vp_p.n94 0.001
R28829 vp_p.n2732 vp_p.n1578 0.001
R28830 vp_p.n4157 vp_p.n3003 0.001
R28831 vp_p.n5581 vp_p.n4427 0.001
R28832 vp_p.n7004 vp_p.n5850 0.001
R28833 vp_p.n8426 vp_p.n7272 0.001
R28834 vp_p.n15730 vp_p.n14576 0.001
R28835 vp_p.n17158 vp_p.n16004 0.001
R28836 vp_p.n18585 vp_p.n17431 0.001
R28837 vp_p.n20011 vp_p.n18857 0.001
R28838 vp_p.n21436 vp_p.n20282 0.001
R28839 vp_p.n22860 vp_p.n21706 0.001
R28840 vp_p.n24283 vp_p.n23129 0.001
R28841 vp_p.n25705 vp_p.n24551 0.001
R28842 vp_p.n27130 vp_p.n25977 0.001
R28843 vp_p.n14331 vp_p.n13237 0.001
R28844 vp_p.n14335 vp_p.n13232 0.001
R28845 vp_p.n12941 vp_p.n11768 0.001
R28846 vp_p.n11503 vp_p.n10330 0.001
R28847 vp_p.n10066 vp_p.n8828 0.001
R28848 vp_p.n1320 vp_p.n89 0.001
R28849 vp_p.n2746 vp_p.n1573 0.001
R28850 vp_p.n4171 vp_p.n2998 0.001
R28851 vp_p.n5595 vp_p.n4422 0.001
R28852 vp_p.n7018 vp_p.n5845 0.001
R28853 vp_p.n8440 vp_p.n7267 0.001
R28854 vp_p.n15744 vp_p.n14571 0.001
R28855 vp_p.n17172 vp_p.n15999 0.001
R28856 vp_p.n18599 vp_p.n17426 0.001
R28857 vp_p.n20025 vp_p.n18852 0.001
R28858 vp_p.n21450 vp_p.n20277 0.001
R28859 vp_p.n22874 vp_p.n21701 0.001
R28860 vp_p.n24297 vp_p.n23124 0.001
R28861 vp_p.n25719 vp_p.n24546 0.001
R28862 vp_p.n27144 vp_p.n25972 0.001
R28863 vp_p.n14339 vp_p.n13227 0.001
R28864 vp_p.n14343 vp_p.n13222 0.001
R28865 vp_p.n12955 vp_p.n11763 0.001
R28866 vp_p.n11517 vp_p.n10325 0.001
R28867 vp_p.n10080 vp_p.n8823 0.001
R28868 vp_p.n1334 vp_p.n84 0.001
R28869 vp_p.n2760 vp_p.n1568 0.001
R28870 vp_p.n4185 vp_p.n2993 0.001
R28871 vp_p.n5609 vp_p.n4417 0.001
R28872 vp_p.n7032 vp_p.n5840 0.001
R28873 vp_p.n8454 vp_p.n7262 0.001
R28874 vp_p.n15758 vp_p.n14566 0.001
R28875 vp_p.n17186 vp_p.n15994 0.001
R28876 vp_p.n18613 vp_p.n17421 0.001
R28877 vp_p.n20039 vp_p.n18847 0.001
R28878 vp_p.n21464 vp_p.n20272 0.001
R28879 vp_p.n22888 vp_p.n21696 0.001
R28880 vp_p.n24311 vp_p.n23119 0.001
R28881 vp_p.n25733 vp_p.n24541 0.001
R28882 vp_p.n27158 vp_p.n25967 0.001
R28883 vp_p.n14347 vp_p.n13217 0.001
R28884 vp_p.n14351 vp_p.n13212 0.001
R28885 vp_p.n12969 vp_p.n11758 0.001
R28886 vp_p.n11531 vp_p.n10320 0.001
R28887 vp_p.n10094 vp_p.n8818 0.001
R28888 vp_p.n1348 vp_p.n79 0.001
R28889 vp_p.n2774 vp_p.n1563 0.001
R28890 vp_p.n4199 vp_p.n2988 0.001
R28891 vp_p.n5623 vp_p.n4412 0.001
R28892 vp_p.n7046 vp_p.n5835 0.001
R28893 vp_p.n8468 vp_p.n7257 0.001
R28894 vp_p.n15772 vp_p.n14561 0.001
R28895 vp_p.n17200 vp_p.n15989 0.001
R28896 vp_p.n18627 vp_p.n17416 0.001
R28897 vp_p.n20053 vp_p.n18842 0.001
R28898 vp_p.n21478 vp_p.n20267 0.001
R28899 vp_p.n22902 vp_p.n21691 0.001
R28900 vp_p.n24325 vp_p.n23114 0.001
R28901 vp_p.n25747 vp_p.n24536 0.001
R28902 vp_p.n27172 vp_p.n25962 0.001
R28903 vp_p.n14355 vp_p.n13207 0.001
R28904 vp_p.n14359 vp_p.n13202 0.001
R28905 vp_p.n12983 vp_p.n11753 0.001
R28906 vp_p.n11545 vp_p.n10315 0.001
R28907 vp_p.n10108 vp_p.n8813 0.001
R28908 vp_p.n1362 vp_p.n74 0.001
R28909 vp_p.n2788 vp_p.n1558 0.001
R28910 vp_p.n4213 vp_p.n2983 0.001
R28911 vp_p.n5637 vp_p.n4407 0.001
R28912 vp_p.n7060 vp_p.n5830 0.001
R28913 vp_p.n8482 vp_p.n7252 0.001
R28914 vp_p.n15786 vp_p.n14556 0.001
R28915 vp_p.n17214 vp_p.n15984 0.001
R28916 vp_p.n18641 vp_p.n17411 0.001
R28917 vp_p.n20067 vp_p.n18837 0.001
R28918 vp_p.n21492 vp_p.n20262 0.001
R28919 vp_p.n22916 vp_p.n21686 0.001
R28920 vp_p.n24339 vp_p.n23109 0.001
R28921 vp_p.n25761 vp_p.n24531 0.001
R28922 vp_p.n27186 vp_p.n25957 0.001
R28923 vp_p.n14363 vp_p.n13197 0.001
R28924 vp_p.n14367 vp_p.n13192 0.001
R28925 vp_p.n12997 vp_p.n11748 0.001
R28926 vp_p.n11559 vp_p.n10310 0.001
R28927 vp_p.n10122 vp_p.n8808 0.001
R28928 vp_p.n1376 vp_p.n69 0.001
R28929 vp_p.n2802 vp_p.n1553 0.001
R28930 vp_p.n4227 vp_p.n2978 0.001
R28931 vp_p.n5651 vp_p.n4402 0.001
R28932 vp_p.n7074 vp_p.n5825 0.001
R28933 vp_p.n8496 vp_p.n7247 0.001
R28934 vp_p.n15800 vp_p.n14551 0.001
R28935 vp_p.n17228 vp_p.n15979 0.001
R28936 vp_p.n18655 vp_p.n17406 0.001
R28937 vp_p.n20081 vp_p.n18832 0.001
R28938 vp_p.n21506 vp_p.n20257 0.001
R28939 vp_p.n22930 vp_p.n21681 0.001
R28940 vp_p.n24353 vp_p.n23104 0.001
R28941 vp_p.n25775 vp_p.n24526 0.001
R28942 vp_p.n27200 vp_p.n25952 0.001
R28943 vp_p.n14371 vp_p.n13187 0.001
R28944 vp_p.n14375 vp_p.n13182 0.001
R28945 vp_p.n15814 vp_p.n14546 0.001
R28946 vp_p.n17242 vp_p.n15974 0.001
R28947 vp_p.n18669 vp_p.n17401 0.001
R28948 vp_p.n20095 vp_p.n18827 0.001
R28949 vp_p.n21520 vp_p.n20252 0.001
R28950 vp_p.n22944 vp_p.n21676 0.001
R28951 vp_p.n24367 vp_p.n23099 0.001
R28952 vp_p.n25789 vp_p.n24521 0.001
R28953 vp_p.n27214 vp_p.n25947 0.001
R28954 vp_p.n13011 vp_p.n11743 0.001
R28955 vp_p.n15818 vp_p.n14541 0.001
R28956 vp_p.n17256 vp_p.n15969 0.001
R28957 vp_p.n18683 vp_p.n17396 0.001
R28958 vp_p.n20109 vp_p.n18822 0.001
R28959 vp_p.n21534 vp_p.n20247 0.001
R28960 vp_p.n22958 vp_p.n21671 0.001
R28961 vp_p.n24381 vp_p.n23094 0.001
R28962 vp_p.n25803 vp_p.n24516 0.001
R28963 vp_p.n27228 vp_p.n25942 0.001
R28964 vp_p.n11587 vp_p.n10300 0.001
R28965 vp_p.n17260 vp_p.n15964 0.001
R28966 vp_p.n18697 vp_p.n17391 0.001
R28967 vp_p.n20123 vp_p.n18817 0.001
R28968 vp_p.n21548 vp_p.n20242 0.001
R28969 vp_p.n22972 vp_p.n21666 0.001
R28970 vp_p.n24395 vp_p.n23089 0.001
R28971 vp_p.n25817 vp_p.n24511 0.001
R28972 vp_p.n27242 vp_p.n25937 0.001
R28973 vp_p.n10164 vp_p.n8793 0.001
R28974 vp_p.n18701 vp_p.n17386 0.001
R28975 vp_p.n20137 vp_p.n18812 0.001
R28976 vp_p.n21562 vp_p.n20237 0.001
R28977 vp_p.n22986 vp_p.n21661 0.001
R28978 vp_p.n24409 vp_p.n23084 0.001
R28979 vp_p.n25831 vp_p.n24506 0.001
R28980 vp_p.n27256 vp_p.n25932 0.001
R28981 vp_p.n1432 vp_p.n49 0.001
R28982 vp_p.n20141 vp_p.n18807 0.001
R28983 vp_p.n21576 vp_p.n20232 0.001
R28984 vp_p.n23000 vp_p.n21656 0.001
R28985 vp_p.n24423 vp_p.n23079 0.001
R28986 vp_p.n25845 vp_p.n24501 0.001
R28987 vp_p.n27270 vp_p.n25927 0.001
R28988 vp_p.n2872 vp_p.n1528 0.001
R28989 vp_p.n21580 vp_p.n20227 0.001
R28990 vp_p.n23014 vp_p.n21651 0.001
R28991 vp_p.n24437 vp_p.n23074 0.001
R28992 vp_p.n25859 vp_p.n24496 0.001
R28993 vp_p.n27284 vp_p.n25922 0.001
R28994 vp_p.n4311 vp_p.n2948 0.001
R28995 vp_p.n23018 vp_p.n21646 0.001
R28996 vp_p.n24451 vp_p.n23069 0.001
R28997 vp_p.n25873 vp_p.n24491 0.001
R28998 vp_p.n27298 vp_p.n25917 0.001
R28999 vp_p.n5749 vp_p.n4367 0.001
R29000 vp_p.n24455 vp_p.n23064 0.001
R29001 vp_p.n25887 vp_p.n24486 0.001
R29002 vp_p.n27312 vp_p.n25912 0.001
R29003 vp_p.n7186 vp_p.n5785 0.001
R29004 vp_p.n25891 vp_p.n24481 0.001
R29005 vp_p.n27326 vp_p.n25907 0.001
R29006 vp_p.n26290 vp_p.n26277 0.001
R29007 vp_p.n12096 vp_p.n12095 0.001
R29008 vp_p.n10658 vp_p.n10657 0.001
R29009 vp_p.n9221 vp_p.n9220 0.001
R29010 vp_p.n475 vp_p.n474 0.001
R29011 vp_p.n1901 vp_p.n1900 0.001
R29012 vp_p.n3326 vp_p.n3325 0.001
R29013 vp_p.n4750 vp_p.n4749 0.001
R29014 vp_p.n6173 vp_p.n6172 0.001
R29015 vp_p.n7595 vp_p.n7594 0.001
R29016 vp_p.n14899 vp_p.n14898 0.001
R29017 vp_p.n16327 vp_p.n16326 0.001
R29018 vp_p.n17754 vp_p.n17753 0.001
R29019 vp_p.n19180 vp_p.n19179 0.001
R29020 vp_p.n20605 vp_p.n20604 0.001
R29021 vp_p.n22029 vp_p.n22028 0.001
R29022 vp_p.n23452 vp_p.n23451 0.001
R29023 vp_p.n24874 vp_p.n24873 0.001
R29024 vp_p.n26299 vp_p.n26298 0.001
R29025 vp_p.n12110 vp_p.n12109 0.001
R29026 vp_p.n10672 vp_p.n10671 0.001
R29027 vp_p.n9235 vp_p.n9234 0.001
R29028 vp_p.n489 vp_p.n488 0.001
R29029 vp_p.n1915 vp_p.n1914 0.001
R29030 vp_p.n3340 vp_p.n3339 0.001
R29031 vp_p.n4764 vp_p.n4763 0.001
R29032 vp_p.n6187 vp_p.n6186 0.001
R29033 vp_p.n7609 vp_p.n7608 0.001
R29034 vp_p.n14913 vp_p.n14912 0.001
R29035 vp_p.n16341 vp_p.n16340 0.001
R29036 vp_p.n17768 vp_p.n17767 0.001
R29037 vp_p.n19194 vp_p.n19193 0.001
R29038 vp_p.n20619 vp_p.n20618 0.001
R29039 vp_p.n22043 vp_p.n22042 0.001
R29040 vp_p.n23466 vp_p.n23465 0.001
R29041 vp_p.n24888 vp_p.n24887 0.001
R29042 vp_p.n26313 vp_p.n26312 0.001
R29043 vp_p.n12124 vp_p.n12123 0.001
R29044 vp_p.n10686 vp_p.n10685 0.001
R29045 vp_p.n9249 vp_p.n9248 0.001
R29046 vp_p.n503 vp_p.n502 0.001
R29047 vp_p.n1929 vp_p.n1928 0.001
R29048 vp_p.n3354 vp_p.n3353 0.001
R29049 vp_p.n4778 vp_p.n4777 0.001
R29050 vp_p.n6201 vp_p.n6200 0.001
R29051 vp_p.n7623 vp_p.n7622 0.001
R29052 vp_p.n14927 vp_p.n14926 0.001
R29053 vp_p.n16355 vp_p.n16354 0.001
R29054 vp_p.n17782 vp_p.n17781 0.001
R29055 vp_p.n19208 vp_p.n19207 0.001
R29056 vp_p.n20633 vp_p.n20632 0.001
R29057 vp_p.n22057 vp_p.n22056 0.001
R29058 vp_p.n23480 vp_p.n23479 0.001
R29059 vp_p.n24902 vp_p.n24901 0.001
R29060 vp_p.n26327 vp_p.n26326 0.001
R29061 vp_p.n12138 vp_p.n12137 0.001
R29062 vp_p.n10700 vp_p.n10699 0.001
R29063 vp_p.n9263 vp_p.n9262 0.001
R29064 vp_p.n517 vp_p.n516 0.001
R29065 vp_p.n1943 vp_p.n1942 0.001
R29066 vp_p.n3368 vp_p.n3367 0.001
R29067 vp_p.n4792 vp_p.n4791 0.001
R29068 vp_p.n6215 vp_p.n6214 0.001
R29069 vp_p.n7637 vp_p.n7636 0.001
R29070 vp_p.n14941 vp_p.n14940 0.001
R29071 vp_p.n16369 vp_p.n16368 0.001
R29072 vp_p.n17796 vp_p.n17795 0.001
R29073 vp_p.n19222 vp_p.n19221 0.001
R29074 vp_p.n20647 vp_p.n20646 0.001
R29075 vp_p.n22071 vp_p.n22070 0.001
R29076 vp_p.n23494 vp_p.n23493 0.001
R29077 vp_p.n24916 vp_p.n24915 0.001
R29078 vp_p.n26341 vp_p.n26340 0.001
R29079 vp_p.n12152 vp_p.n12151 0.001
R29080 vp_p.n10714 vp_p.n10713 0.001
R29081 vp_p.n9277 vp_p.n9276 0.001
R29082 vp_p.n531 vp_p.n530 0.001
R29083 vp_p.n1957 vp_p.n1956 0.001
R29084 vp_p.n3382 vp_p.n3381 0.001
R29085 vp_p.n4806 vp_p.n4805 0.001
R29086 vp_p.n6229 vp_p.n6228 0.001
R29087 vp_p.n7651 vp_p.n7650 0.001
R29088 vp_p.n14955 vp_p.n14954 0.001
R29089 vp_p.n16383 vp_p.n16382 0.001
R29090 vp_p.n17810 vp_p.n17809 0.001
R29091 vp_p.n19236 vp_p.n19235 0.001
R29092 vp_p.n20661 vp_p.n20660 0.001
R29093 vp_p.n22085 vp_p.n22084 0.001
R29094 vp_p.n23508 vp_p.n23507 0.001
R29095 vp_p.n24930 vp_p.n24929 0.001
R29096 vp_p.n26355 vp_p.n26354 0.001
R29097 vp_p.n12166 vp_p.n12165 0.001
R29098 vp_p.n10728 vp_p.n10727 0.001
R29099 vp_p.n9291 vp_p.n9290 0.001
R29100 vp_p.n545 vp_p.n544 0.001
R29101 vp_p.n1971 vp_p.n1970 0.001
R29102 vp_p.n3396 vp_p.n3395 0.001
R29103 vp_p.n4820 vp_p.n4819 0.001
R29104 vp_p.n6243 vp_p.n6242 0.001
R29105 vp_p.n7665 vp_p.n7664 0.001
R29106 vp_p.n14969 vp_p.n14968 0.001
R29107 vp_p.n16397 vp_p.n16396 0.001
R29108 vp_p.n17824 vp_p.n17823 0.001
R29109 vp_p.n19250 vp_p.n19249 0.001
R29110 vp_p.n20675 vp_p.n20674 0.001
R29111 vp_p.n22099 vp_p.n22098 0.001
R29112 vp_p.n23522 vp_p.n23521 0.001
R29113 vp_p.n24944 vp_p.n24943 0.001
R29114 vp_p.n26369 vp_p.n26368 0.001
R29115 vp_p.n12180 vp_p.n12179 0.001
R29116 vp_p.n10742 vp_p.n10741 0.001
R29117 vp_p.n9305 vp_p.n9304 0.001
R29118 vp_p.n559 vp_p.n558 0.001
R29119 vp_p.n1985 vp_p.n1984 0.001
R29120 vp_p.n3410 vp_p.n3409 0.001
R29121 vp_p.n4834 vp_p.n4833 0.001
R29122 vp_p.n6257 vp_p.n6256 0.001
R29123 vp_p.n7679 vp_p.n7678 0.001
R29124 vp_p.n14983 vp_p.n14982 0.001
R29125 vp_p.n16411 vp_p.n16410 0.001
R29126 vp_p.n17838 vp_p.n17837 0.001
R29127 vp_p.n19264 vp_p.n19263 0.001
R29128 vp_p.n20689 vp_p.n20688 0.001
R29129 vp_p.n22113 vp_p.n22112 0.001
R29130 vp_p.n23536 vp_p.n23535 0.001
R29131 vp_p.n24958 vp_p.n24957 0.001
R29132 vp_p.n26383 vp_p.n26382 0.001
R29133 vp_p.n12194 vp_p.n12193 0.001
R29134 vp_p.n10756 vp_p.n10755 0.001
R29135 vp_p.n9319 vp_p.n9318 0.001
R29136 vp_p.n573 vp_p.n572 0.001
R29137 vp_p.n1999 vp_p.n1998 0.001
R29138 vp_p.n3424 vp_p.n3423 0.001
R29139 vp_p.n4848 vp_p.n4847 0.001
R29140 vp_p.n6271 vp_p.n6270 0.001
R29141 vp_p.n7693 vp_p.n7692 0.001
R29142 vp_p.n14997 vp_p.n14996 0.001
R29143 vp_p.n16425 vp_p.n16424 0.001
R29144 vp_p.n17852 vp_p.n17851 0.001
R29145 vp_p.n19278 vp_p.n19277 0.001
R29146 vp_p.n20703 vp_p.n20702 0.001
R29147 vp_p.n22127 vp_p.n22126 0.001
R29148 vp_p.n23550 vp_p.n23549 0.001
R29149 vp_p.n24972 vp_p.n24971 0.001
R29150 vp_p.n26397 vp_p.n26396 0.001
R29151 vp_p.n12208 vp_p.n12207 0.001
R29152 vp_p.n10770 vp_p.n10769 0.001
R29153 vp_p.n9333 vp_p.n9332 0.001
R29154 vp_p.n587 vp_p.n586 0.001
R29155 vp_p.n2013 vp_p.n2012 0.001
R29156 vp_p.n3438 vp_p.n3437 0.001
R29157 vp_p.n4862 vp_p.n4861 0.001
R29158 vp_p.n6285 vp_p.n6284 0.001
R29159 vp_p.n7707 vp_p.n7706 0.001
R29160 vp_p.n15011 vp_p.n15010 0.001
R29161 vp_p.n16439 vp_p.n16438 0.001
R29162 vp_p.n17866 vp_p.n17865 0.001
R29163 vp_p.n19292 vp_p.n19291 0.001
R29164 vp_p.n20717 vp_p.n20716 0.001
R29165 vp_p.n22141 vp_p.n22140 0.001
R29166 vp_p.n23564 vp_p.n23563 0.001
R29167 vp_p.n24986 vp_p.n24985 0.001
R29168 vp_p.n26411 vp_p.n26410 0.001
R29169 vp_p.n12222 vp_p.n12221 0.001
R29170 vp_p.n10784 vp_p.n10783 0.001
R29171 vp_p.n9347 vp_p.n9346 0.001
R29172 vp_p.n601 vp_p.n600 0.001
R29173 vp_p.n2027 vp_p.n2026 0.001
R29174 vp_p.n3452 vp_p.n3451 0.001
R29175 vp_p.n4876 vp_p.n4875 0.001
R29176 vp_p.n6299 vp_p.n6298 0.001
R29177 vp_p.n7721 vp_p.n7720 0.001
R29178 vp_p.n15025 vp_p.n15024 0.001
R29179 vp_p.n16453 vp_p.n16452 0.001
R29180 vp_p.n17880 vp_p.n17879 0.001
R29181 vp_p.n19306 vp_p.n19305 0.001
R29182 vp_p.n20731 vp_p.n20730 0.001
R29183 vp_p.n22155 vp_p.n22154 0.001
R29184 vp_p.n23578 vp_p.n23577 0.001
R29185 vp_p.n25000 vp_p.n24999 0.001
R29186 vp_p.n26425 vp_p.n26424 0.001
R29187 vp_p.n12236 vp_p.n12235 0.001
R29188 vp_p.n10798 vp_p.n10797 0.001
R29189 vp_p.n9361 vp_p.n9360 0.001
R29190 vp_p.n615 vp_p.n614 0.001
R29191 vp_p.n2041 vp_p.n2040 0.001
R29192 vp_p.n3466 vp_p.n3465 0.001
R29193 vp_p.n4890 vp_p.n4889 0.001
R29194 vp_p.n6313 vp_p.n6312 0.001
R29195 vp_p.n7735 vp_p.n7734 0.001
R29196 vp_p.n15039 vp_p.n15038 0.001
R29197 vp_p.n16467 vp_p.n16466 0.001
R29198 vp_p.n17894 vp_p.n17893 0.001
R29199 vp_p.n19320 vp_p.n19319 0.001
R29200 vp_p.n20745 vp_p.n20744 0.001
R29201 vp_p.n22169 vp_p.n22168 0.001
R29202 vp_p.n23592 vp_p.n23591 0.001
R29203 vp_p.n25014 vp_p.n25013 0.001
R29204 vp_p.n26439 vp_p.n26438 0.001
R29205 vp_p.n12250 vp_p.n12249 0.001
R29206 vp_p.n10812 vp_p.n10811 0.001
R29207 vp_p.n9375 vp_p.n9374 0.001
R29208 vp_p.n629 vp_p.n628 0.001
R29209 vp_p.n2055 vp_p.n2054 0.001
R29210 vp_p.n3480 vp_p.n3479 0.001
R29211 vp_p.n4904 vp_p.n4903 0.001
R29212 vp_p.n6327 vp_p.n6326 0.001
R29213 vp_p.n7749 vp_p.n7748 0.001
R29214 vp_p.n15053 vp_p.n15052 0.001
R29215 vp_p.n16481 vp_p.n16480 0.001
R29216 vp_p.n17908 vp_p.n17907 0.001
R29217 vp_p.n19334 vp_p.n19333 0.001
R29218 vp_p.n20759 vp_p.n20758 0.001
R29219 vp_p.n22183 vp_p.n22182 0.001
R29220 vp_p.n23606 vp_p.n23605 0.001
R29221 vp_p.n25028 vp_p.n25027 0.001
R29222 vp_p.n26453 vp_p.n26452 0.001
R29223 vp_p.n12264 vp_p.n12263 0.001
R29224 vp_p.n10826 vp_p.n10825 0.001
R29225 vp_p.n9389 vp_p.n9388 0.001
R29226 vp_p.n643 vp_p.n642 0.001
R29227 vp_p.n2069 vp_p.n2068 0.001
R29228 vp_p.n3494 vp_p.n3493 0.001
R29229 vp_p.n4918 vp_p.n4917 0.001
R29230 vp_p.n6341 vp_p.n6340 0.001
R29231 vp_p.n7763 vp_p.n7762 0.001
R29232 vp_p.n15067 vp_p.n15066 0.001
R29233 vp_p.n16495 vp_p.n16494 0.001
R29234 vp_p.n17922 vp_p.n17921 0.001
R29235 vp_p.n19348 vp_p.n19347 0.001
R29236 vp_p.n20773 vp_p.n20772 0.001
R29237 vp_p.n22197 vp_p.n22196 0.001
R29238 vp_p.n23620 vp_p.n23619 0.001
R29239 vp_p.n25042 vp_p.n25041 0.001
R29240 vp_p.n26467 vp_p.n26466 0.001
R29241 vp_p.n12278 vp_p.n12277 0.001
R29242 vp_p.n10840 vp_p.n10839 0.001
R29243 vp_p.n9403 vp_p.n9402 0.001
R29244 vp_p.n657 vp_p.n656 0.001
R29245 vp_p.n2083 vp_p.n2082 0.001
R29246 vp_p.n3508 vp_p.n3507 0.001
R29247 vp_p.n4932 vp_p.n4931 0.001
R29248 vp_p.n6355 vp_p.n6354 0.001
R29249 vp_p.n7777 vp_p.n7776 0.001
R29250 vp_p.n15081 vp_p.n15080 0.001
R29251 vp_p.n16509 vp_p.n16508 0.001
R29252 vp_p.n17936 vp_p.n17935 0.001
R29253 vp_p.n19362 vp_p.n19361 0.001
R29254 vp_p.n20787 vp_p.n20786 0.001
R29255 vp_p.n22211 vp_p.n22210 0.001
R29256 vp_p.n23634 vp_p.n23633 0.001
R29257 vp_p.n25056 vp_p.n25055 0.001
R29258 vp_p.n26481 vp_p.n26480 0.001
R29259 vp_p.n12292 vp_p.n12291 0.001
R29260 vp_p.n10854 vp_p.n10853 0.001
R29261 vp_p.n9417 vp_p.n9416 0.001
R29262 vp_p.n671 vp_p.n670 0.001
R29263 vp_p.n2097 vp_p.n2096 0.001
R29264 vp_p.n3522 vp_p.n3521 0.001
R29265 vp_p.n4946 vp_p.n4945 0.001
R29266 vp_p.n6369 vp_p.n6368 0.001
R29267 vp_p.n7791 vp_p.n7790 0.001
R29268 vp_p.n15095 vp_p.n15094 0.001
R29269 vp_p.n16523 vp_p.n16522 0.001
R29270 vp_p.n17950 vp_p.n17949 0.001
R29271 vp_p.n19376 vp_p.n19375 0.001
R29272 vp_p.n20801 vp_p.n20800 0.001
R29273 vp_p.n22225 vp_p.n22224 0.001
R29274 vp_p.n23648 vp_p.n23647 0.001
R29275 vp_p.n25070 vp_p.n25069 0.001
R29276 vp_p.n26495 vp_p.n26494 0.001
R29277 vp_p.n12306 vp_p.n12305 0.001
R29278 vp_p.n10868 vp_p.n10867 0.001
R29279 vp_p.n9431 vp_p.n9430 0.001
R29280 vp_p.n685 vp_p.n684 0.001
R29281 vp_p.n2111 vp_p.n2110 0.001
R29282 vp_p.n3536 vp_p.n3535 0.001
R29283 vp_p.n4960 vp_p.n4959 0.001
R29284 vp_p.n6383 vp_p.n6382 0.001
R29285 vp_p.n7805 vp_p.n7804 0.001
R29286 vp_p.n15109 vp_p.n15108 0.001
R29287 vp_p.n16537 vp_p.n16536 0.001
R29288 vp_p.n17964 vp_p.n17963 0.001
R29289 vp_p.n19390 vp_p.n19389 0.001
R29290 vp_p.n20815 vp_p.n20814 0.001
R29291 vp_p.n22239 vp_p.n22238 0.001
R29292 vp_p.n23662 vp_p.n23661 0.001
R29293 vp_p.n25084 vp_p.n25083 0.001
R29294 vp_p.n26509 vp_p.n26508 0.001
R29295 vp_p.n12320 vp_p.n12319 0.001
R29296 vp_p.n10882 vp_p.n10881 0.001
R29297 vp_p.n9445 vp_p.n9444 0.001
R29298 vp_p.n699 vp_p.n698 0.001
R29299 vp_p.n2125 vp_p.n2124 0.001
R29300 vp_p.n3550 vp_p.n3549 0.001
R29301 vp_p.n4974 vp_p.n4973 0.001
R29302 vp_p.n6397 vp_p.n6396 0.001
R29303 vp_p.n7819 vp_p.n7818 0.001
R29304 vp_p.n15123 vp_p.n15122 0.001
R29305 vp_p.n16551 vp_p.n16550 0.001
R29306 vp_p.n17978 vp_p.n17977 0.001
R29307 vp_p.n19404 vp_p.n19403 0.001
R29308 vp_p.n20829 vp_p.n20828 0.001
R29309 vp_p.n22253 vp_p.n22252 0.001
R29310 vp_p.n23676 vp_p.n23675 0.001
R29311 vp_p.n25098 vp_p.n25097 0.001
R29312 vp_p.n26523 vp_p.n26522 0.001
R29313 vp_p.n12334 vp_p.n12333 0.001
R29314 vp_p.n10896 vp_p.n10895 0.001
R29315 vp_p.n9459 vp_p.n9458 0.001
R29316 vp_p.n713 vp_p.n712 0.001
R29317 vp_p.n2139 vp_p.n2138 0.001
R29318 vp_p.n3564 vp_p.n3563 0.001
R29319 vp_p.n4988 vp_p.n4987 0.001
R29320 vp_p.n6411 vp_p.n6410 0.001
R29321 vp_p.n7833 vp_p.n7832 0.001
R29322 vp_p.n15137 vp_p.n15136 0.001
R29323 vp_p.n16565 vp_p.n16564 0.001
R29324 vp_p.n17992 vp_p.n17991 0.001
R29325 vp_p.n19418 vp_p.n19417 0.001
R29326 vp_p.n20843 vp_p.n20842 0.001
R29327 vp_p.n22267 vp_p.n22266 0.001
R29328 vp_p.n23690 vp_p.n23689 0.001
R29329 vp_p.n25112 vp_p.n25111 0.001
R29330 vp_p.n26537 vp_p.n26536 0.001
R29331 vp_p.n12348 vp_p.n12347 0.001
R29332 vp_p.n10910 vp_p.n10909 0.001
R29333 vp_p.n9473 vp_p.n9472 0.001
R29334 vp_p.n727 vp_p.n726 0.001
R29335 vp_p.n2153 vp_p.n2152 0.001
R29336 vp_p.n3578 vp_p.n3577 0.001
R29337 vp_p.n5002 vp_p.n5001 0.001
R29338 vp_p.n6425 vp_p.n6424 0.001
R29339 vp_p.n7847 vp_p.n7846 0.001
R29340 vp_p.n15151 vp_p.n15150 0.001
R29341 vp_p.n16579 vp_p.n16578 0.001
R29342 vp_p.n18006 vp_p.n18005 0.001
R29343 vp_p.n19432 vp_p.n19431 0.001
R29344 vp_p.n20857 vp_p.n20856 0.001
R29345 vp_p.n22281 vp_p.n22280 0.001
R29346 vp_p.n23704 vp_p.n23703 0.001
R29347 vp_p.n25126 vp_p.n25125 0.001
R29348 vp_p.n26551 vp_p.n26550 0.001
R29349 vp_p.n12362 vp_p.n12361 0.001
R29350 vp_p.n10924 vp_p.n10923 0.001
R29351 vp_p.n9487 vp_p.n9486 0.001
R29352 vp_p.n741 vp_p.n740 0.001
R29353 vp_p.n2167 vp_p.n2166 0.001
R29354 vp_p.n3592 vp_p.n3591 0.001
R29355 vp_p.n5016 vp_p.n5015 0.001
R29356 vp_p.n6439 vp_p.n6438 0.001
R29357 vp_p.n7861 vp_p.n7860 0.001
R29358 vp_p.n15165 vp_p.n15164 0.001
R29359 vp_p.n16593 vp_p.n16592 0.001
R29360 vp_p.n18020 vp_p.n18019 0.001
R29361 vp_p.n19446 vp_p.n19445 0.001
R29362 vp_p.n20871 vp_p.n20870 0.001
R29363 vp_p.n22295 vp_p.n22294 0.001
R29364 vp_p.n23718 vp_p.n23717 0.001
R29365 vp_p.n25140 vp_p.n25139 0.001
R29366 vp_p.n26565 vp_p.n26564 0.001
R29367 vp_p.n12376 vp_p.n12375 0.001
R29368 vp_p.n10938 vp_p.n10937 0.001
R29369 vp_p.n9501 vp_p.n9500 0.001
R29370 vp_p.n755 vp_p.n754 0.001
R29371 vp_p.n2181 vp_p.n2180 0.001
R29372 vp_p.n3606 vp_p.n3605 0.001
R29373 vp_p.n5030 vp_p.n5029 0.001
R29374 vp_p.n6453 vp_p.n6452 0.001
R29375 vp_p.n7875 vp_p.n7874 0.001
R29376 vp_p.n15179 vp_p.n15178 0.001
R29377 vp_p.n16607 vp_p.n16606 0.001
R29378 vp_p.n18034 vp_p.n18033 0.001
R29379 vp_p.n19460 vp_p.n19459 0.001
R29380 vp_p.n20885 vp_p.n20884 0.001
R29381 vp_p.n22309 vp_p.n22308 0.001
R29382 vp_p.n23732 vp_p.n23731 0.001
R29383 vp_p.n25154 vp_p.n25153 0.001
R29384 vp_p.n26579 vp_p.n26578 0.001
R29385 vp_p.n12390 vp_p.n12389 0.001
R29386 vp_p.n10952 vp_p.n10951 0.001
R29387 vp_p.n9515 vp_p.n9514 0.001
R29388 vp_p.n769 vp_p.n768 0.001
R29389 vp_p.n2195 vp_p.n2194 0.001
R29390 vp_p.n3620 vp_p.n3619 0.001
R29391 vp_p.n5044 vp_p.n5043 0.001
R29392 vp_p.n6467 vp_p.n6466 0.001
R29393 vp_p.n7889 vp_p.n7888 0.001
R29394 vp_p.n15193 vp_p.n15192 0.001
R29395 vp_p.n16621 vp_p.n16620 0.001
R29396 vp_p.n18048 vp_p.n18047 0.001
R29397 vp_p.n19474 vp_p.n19473 0.001
R29398 vp_p.n20899 vp_p.n20898 0.001
R29399 vp_p.n22323 vp_p.n22322 0.001
R29400 vp_p.n23746 vp_p.n23745 0.001
R29401 vp_p.n25168 vp_p.n25167 0.001
R29402 vp_p.n26593 vp_p.n26592 0.001
R29403 vp_p.n12404 vp_p.n12403 0.001
R29404 vp_p.n10966 vp_p.n10965 0.001
R29405 vp_p.n9529 vp_p.n9528 0.001
R29406 vp_p.n783 vp_p.n782 0.001
R29407 vp_p.n2209 vp_p.n2208 0.001
R29408 vp_p.n3634 vp_p.n3633 0.001
R29409 vp_p.n5058 vp_p.n5057 0.001
R29410 vp_p.n6481 vp_p.n6480 0.001
R29411 vp_p.n7903 vp_p.n7902 0.001
R29412 vp_p.n15207 vp_p.n15206 0.001
R29413 vp_p.n16635 vp_p.n16634 0.001
R29414 vp_p.n18062 vp_p.n18061 0.001
R29415 vp_p.n19488 vp_p.n19487 0.001
R29416 vp_p.n20913 vp_p.n20912 0.001
R29417 vp_p.n22337 vp_p.n22336 0.001
R29418 vp_p.n23760 vp_p.n23759 0.001
R29419 vp_p.n25182 vp_p.n25181 0.001
R29420 vp_p.n26607 vp_p.n26606 0.001
R29421 vp_p.n12418 vp_p.n12417 0.001
R29422 vp_p.n10980 vp_p.n10979 0.001
R29423 vp_p.n9543 vp_p.n9542 0.001
R29424 vp_p.n797 vp_p.n796 0.001
R29425 vp_p.n2223 vp_p.n2222 0.001
R29426 vp_p.n3648 vp_p.n3647 0.001
R29427 vp_p.n5072 vp_p.n5071 0.001
R29428 vp_p.n6495 vp_p.n6494 0.001
R29429 vp_p.n7917 vp_p.n7916 0.001
R29430 vp_p.n15221 vp_p.n15220 0.001
R29431 vp_p.n16649 vp_p.n16648 0.001
R29432 vp_p.n18076 vp_p.n18075 0.001
R29433 vp_p.n19502 vp_p.n19501 0.001
R29434 vp_p.n20927 vp_p.n20926 0.001
R29435 vp_p.n22351 vp_p.n22350 0.001
R29436 vp_p.n23774 vp_p.n23773 0.001
R29437 vp_p.n25196 vp_p.n25195 0.001
R29438 vp_p.n26621 vp_p.n26620 0.001
R29439 vp_p.n12432 vp_p.n12431 0.001
R29440 vp_p.n10994 vp_p.n10993 0.001
R29441 vp_p.n9557 vp_p.n9556 0.001
R29442 vp_p.n811 vp_p.n810 0.001
R29443 vp_p.n2237 vp_p.n2236 0.001
R29444 vp_p.n3662 vp_p.n3661 0.001
R29445 vp_p.n5086 vp_p.n5085 0.001
R29446 vp_p.n6509 vp_p.n6508 0.001
R29447 vp_p.n7931 vp_p.n7930 0.001
R29448 vp_p.n15235 vp_p.n15234 0.001
R29449 vp_p.n16663 vp_p.n16662 0.001
R29450 vp_p.n18090 vp_p.n18089 0.001
R29451 vp_p.n19516 vp_p.n19515 0.001
R29452 vp_p.n20941 vp_p.n20940 0.001
R29453 vp_p.n22365 vp_p.n22364 0.001
R29454 vp_p.n23788 vp_p.n23787 0.001
R29455 vp_p.n25210 vp_p.n25209 0.001
R29456 vp_p.n26635 vp_p.n26634 0.001
R29457 vp_p.n12446 vp_p.n12445 0.001
R29458 vp_p.n11008 vp_p.n11007 0.001
R29459 vp_p.n9571 vp_p.n9570 0.001
R29460 vp_p.n825 vp_p.n824 0.001
R29461 vp_p.n2251 vp_p.n2250 0.001
R29462 vp_p.n3676 vp_p.n3675 0.001
R29463 vp_p.n5100 vp_p.n5099 0.001
R29464 vp_p.n6523 vp_p.n6522 0.001
R29465 vp_p.n7945 vp_p.n7944 0.001
R29466 vp_p.n15249 vp_p.n15248 0.001
R29467 vp_p.n16677 vp_p.n16676 0.001
R29468 vp_p.n18104 vp_p.n18103 0.001
R29469 vp_p.n19530 vp_p.n19529 0.001
R29470 vp_p.n20955 vp_p.n20954 0.001
R29471 vp_p.n22379 vp_p.n22378 0.001
R29472 vp_p.n23802 vp_p.n23801 0.001
R29473 vp_p.n25224 vp_p.n25223 0.001
R29474 vp_p.n26649 vp_p.n26648 0.001
R29475 vp_p.n12460 vp_p.n12459 0.001
R29476 vp_p.n11022 vp_p.n11021 0.001
R29477 vp_p.n9585 vp_p.n9584 0.001
R29478 vp_p.n839 vp_p.n838 0.001
R29479 vp_p.n2265 vp_p.n2264 0.001
R29480 vp_p.n3690 vp_p.n3689 0.001
R29481 vp_p.n5114 vp_p.n5113 0.001
R29482 vp_p.n6537 vp_p.n6536 0.001
R29483 vp_p.n7959 vp_p.n7958 0.001
R29484 vp_p.n15263 vp_p.n15262 0.001
R29485 vp_p.n16691 vp_p.n16690 0.001
R29486 vp_p.n18118 vp_p.n18117 0.001
R29487 vp_p.n19544 vp_p.n19543 0.001
R29488 vp_p.n20969 vp_p.n20968 0.001
R29489 vp_p.n22393 vp_p.n22392 0.001
R29490 vp_p.n23816 vp_p.n23815 0.001
R29491 vp_p.n25238 vp_p.n25237 0.001
R29492 vp_p.n26663 vp_p.n26662 0.001
R29493 vp_p.n12474 vp_p.n12473 0.001
R29494 vp_p.n11036 vp_p.n11035 0.001
R29495 vp_p.n9599 vp_p.n9598 0.001
R29496 vp_p.n853 vp_p.n852 0.001
R29497 vp_p.n2279 vp_p.n2278 0.001
R29498 vp_p.n3704 vp_p.n3703 0.001
R29499 vp_p.n5128 vp_p.n5127 0.001
R29500 vp_p.n6551 vp_p.n6550 0.001
R29501 vp_p.n7973 vp_p.n7972 0.001
R29502 vp_p.n15277 vp_p.n15276 0.001
R29503 vp_p.n16705 vp_p.n16704 0.001
R29504 vp_p.n18132 vp_p.n18131 0.001
R29505 vp_p.n19558 vp_p.n19557 0.001
R29506 vp_p.n20983 vp_p.n20982 0.001
R29507 vp_p.n22407 vp_p.n22406 0.001
R29508 vp_p.n23830 vp_p.n23829 0.001
R29509 vp_p.n25252 vp_p.n25251 0.001
R29510 vp_p.n26677 vp_p.n26676 0.001
R29511 vp_p.n12488 vp_p.n12487 0.001
R29512 vp_p.n11050 vp_p.n11049 0.001
R29513 vp_p.n9613 vp_p.n9612 0.001
R29514 vp_p.n867 vp_p.n866 0.001
R29515 vp_p.n2293 vp_p.n2292 0.001
R29516 vp_p.n3718 vp_p.n3717 0.001
R29517 vp_p.n5142 vp_p.n5141 0.001
R29518 vp_p.n6565 vp_p.n6564 0.001
R29519 vp_p.n7987 vp_p.n7986 0.001
R29520 vp_p.n15291 vp_p.n15290 0.001
R29521 vp_p.n16719 vp_p.n16718 0.001
R29522 vp_p.n18146 vp_p.n18145 0.001
R29523 vp_p.n19572 vp_p.n19571 0.001
R29524 vp_p.n20997 vp_p.n20996 0.001
R29525 vp_p.n22421 vp_p.n22420 0.001
R29526 vp_p.n23844 vp_p.n23843 0.001
R29527 vp_p.n25266 vp_p.n25265 0.001
R29528 vp_p.n26691 vp_p.n26690 0.001
R29529 vp_p.n12502 vp_p.n12501 0.001
R29530 vp_p.n11064 vp_p.n11063 0.001
R29531 vp_p.n9627 vp_p.n9626 0.001
R29532 vp_p.n881 vp_p.n880 0.001
R29533 vp_p.n2307 vp_p.n2306 0.001
R29534 vp_p.n3732 vp_p.n3731 0.001
R29535 vp_p.n5156 vp_p.n5155 0.001
R29536 vp_p.n6579 vp_p.n6578 0.001
R29537 vp_p.n8001 vp_p.n8000 0.001
R29538 vp_p.n15305 vp_p.n15304 0.001
R29539 vp_p.n16733 vp_p.n16732 0.001
R29540 vp_p.n18160 vp_p.n18159 0.001
R29541 vp_p.n19586 vp_p.n19585 0.001
R29542 vp_p.n21011 vp_p.n21010 0.001
R29543 vp_p.n22435 vp_p.n22434 0.001
R29544 vp_p.n23858 vp_p.n23857 0.001
R29545 vp_p.n25280 vp_p.n25279 0.001
R29546 vp_p.n26705 vp_p.n26704 0.001
R29547 vp_p.n12516 vp_p.n12515 0.001
R29548 vp_p.n11078 vp_p.n11077 0.001
R29549 vp_p.n9641 vp_p.n9640 0.001
R29550 vp_p.n895 vp_p.n894 0.001
R29551 vp_p.n2321 vp_p.n2320 0.001
R29552 vp_p.n3746 vp_p.n3745 0.001
R29553 vp_p.n5170 vp_p.n5169 0.001
R29554 vp_p.n6593 vp_p.n6592 0.001
R29555 vp_p.n8015 vp_p.n8014 0.001
R29556 vp_p.n15319 vp_p.n15318 0.001
R29557 vp_p.n16747 vp_p.n16746 0.001
R29558 vp_p.n18174 vp_p.n18173 0.001
R29559 vp_p.n19600 vp_p.n19599 0.001
R29560 vp_p.n21025 vp_p.n21024 0.001
R29561 vp_p.n22449 vp_p.n22448 0.001
R29562 vp_p.n23872 vp_p.n23871 0.001
R29563 vp_p.n25294 vp_p.n25293 0.001
R29564 vp_p.n26719 vp_p.n26718 0.001
R29565 vp_p.n12530 vp_p.n12529 0.001
R29566 vp_p.n11092 vp_p.n11091 0.001
R29567 vp_p.n9655 vp_p.n9654 0.001
R29568 vp_p.n909 vp_p.n908 0.001
R29569 vp_p.n2335 vp_p.n2334 0.001
R29570 vp_p.n3760 vp_p.n3759 0.001
R29571 vp_p.n5184 vp_p.n5183 0.001
R29572 vp_p.n6607 vp_p.n6606 0.001
R29573 vp_p.n8029 vp_p.n8028 0.001
R29574 vp_p.n15333 vp_p.n15332 0.001
R29575 vp_p.n16761 vp_p.n16760 0.001
R29576 vp_p.n18188 vp_p.n18187 0.001
R29577 vp_p.n19614 vp_p.n19613 0.001
R29578 vp_p.n21039 vp_p.n21038 0.001
R29579 vp_p.n22463 vp_p.n22462 0.001
R29580 vp_p.n23886 vp_p.n23885 0.001
R29581 vp_p.n25308 vp_p.n25307 0.001
R29582 vp_p.n26733 vp_p.n26732 0.001
R29583 vp_p.n12544 vp_p.n12543 0.001
R29584 vp_p.n11106 vp_p.n11105 0.001
R29585 vp_p.n9669 vp_p.n9668 0.001
R29586 vp_p.n923 vp_p.n922 0.001
R29587 vp_p.n2349 vp_p.n2348 0.001
R29588 vp_p.n3774 vp_p.n3773 0.001
R29589 vp_p.n5198 vp_p.n5197 0.001
R29590 vp_p.n6621 vp_p.n6620 0.001
R29591 vp_p.n8043 vp_p.n8042 0.001
R29592 vp_p.n15347 vp_p.n15346 0.001
R29593 vp_p.n16775 vp_p.n16774 0.001
R29594 vp_p.n18202 vp_p.n18201 0.001
R29595 vp_p.n19628 vp_p.n19627 0.001
R29596 vp_p.n21053 vp_p.n21052 0.001
R29597 vp_p.n22477 vp_p.n22476 0.001
R29598 vp_p.n23900 vp_p.n23899 0.001
R29599 vp_p.n25322 vp_p.n25321 0.001
R29600 vp_p.n26747 vp_p.n26746 0.001
R29601 vp_p.n12558 vp_p.n12557 0.001
R29602 vp_p.n11120 vp_p.n11119 0.001
R29603 vp_p.n9683 vp_p.n9682 0.001
R29604 vp_p.n937 vp_p.n936 0.001
R29605 vp_p.n2363 vp_p.n2362 0.001
R29606 vp_p.n3788 vp_p.n3787 0.001
R29607 vp_p.n5212 vp_p.n5211 0.001
R29608 vp_p.n6635 vp_p.n6634 0.001
R29609 vp_p.n8057 vp_p.n8056 0.001
R29610 vp_p.n15361 vp_p.n15360 0.001
R29611 vp_p.n16789 vp_p.n16788 0.001
R29612 vp_p.n18216 vp_p.n18215 0.001
R29613 vp_p.n19642 vp_p.n19641 0.001
R29614 vp_p.n21067 vp_p.n21066 0.001
R29615 vp_p.n22491 vp_p.n22490 0.001
R29616 vp_p.n23914 vp_p.n23913 0.001
R29617 vp_p.n25336 vp_p.n25335 0.001
R29618 vp_p.n26761 vp_p.n26760 0.001
R29619 vp_p.n12572 vp_p.n12571 0.001
R29620 vp_p.n11134 vp_p.n11133 0.001
R29621 vp_p.n9697 vp_p.n9696 0.001
R29622 vp_p.n951 vp_p.n950 0.001
R29623 vp_p.n2377 vp_p.n2376 0.001
R29624 vp_p.n3802 vp_p.n3801 0.001
R29625 vp_p.n5226 vp_p.n5225 0.001
R29626 vp_p.n6649 vp_p.n6648 0.001
R29627 vp_p.n8071 vp_p.n8070 0.001
R29628 vp_p.n15375 vp_p.n15374 0.001
R29629 vp_p.n16803 vp_p.n16802 0.001
R29630 vp_p.n18230 vp_p.n18229 0.001
R29631 vp_p.n19656 vp_p.n19655 0.001
R29632 vp_p.n21081 vp_p.n21080 0.001
R29633 vp_p.n22505 vp_p.n22504 0.001
R29634 vp_p.n23928 vp_p.n23927 0.001
R29635 vp_p.n25350 vp_p.n25349 0.001
R29636 vp_p.n26775 vp_p.n26774 0.001
R29637 vp_p.n12586 vp_p.n12585 0.001
R29638 vp_p.n11148 vp_p.n11147 0.001
R29639 vp_p.n9711 vp_p.n9710 0.001
R29640 vp_p.n965 vp_p.n964 0.001
R29641 vp_p.n2391 vp_p.n2390 0.001
R29642 vp_p.n3816 vp_p.n3815 0.001
R29643 vp_p.n5240 vp_p.n5239 0.001
R29644 vp_p.n6663 vp_p.n6662 0.001
R29645 vp_p.n8085 vp_p.n8084 0.001
R29646 vp_p.n15389 vp_p.n15388 0.001
R29647 vp_p.n16817 vp_p.n16816 0.001
R29648 vp_p.n18244 vp_p.n18243 0.001
R29649 vp_p.n19670 vp_p.n19669 0.001
R29650 vp_p.n21095 vp_p.n21094 0.001
R29651 vp_p.n22519 vp_p.n22518 0.001
R29652 vp_p.n23942 vp_p.n23941 0.001
R29653 vp_p.n25364 vp_p.n25363 0.001
R29654 vp_p.n26789 vp_p.n26788 0.001
R29655 vp_p.n12600 vp_p.n12599 0.001
R29656 vp_p.n11162 vp_p.n11161 0.001
R29657 vp_p.n9725 vp_p.n9724 0.001
R29658 vp_p.n979 vp_p.n978 0.001
R29659 vp_p.n2405 vp_p.n2404 0.001
R29660 vp_p.n3830 vp_p.n3829 0.001
R29661 vp_p.n5254 vp_p.n5253 0.001
R29662 vp_p.n6677 vp_p.n6676 0.001
R29663 vp_p.n8099 vp_p.n8098 0.001
R29664 vp_p.n15403 vp_p.n15402 0.001
R29665 vp_p.n16831 vp_p.n16830 0.001
R29666 vp_p.n18258 vp_p.n18257 0.001
R29667 vp_p.n19684 vp_p.n19683 0.001
R29668 vp_p.n21109 vp_p.n21108 0.001
R29669 vp_p.n22533 vp_p.n22532 0.001
R29670 vp_p.n23956 vp_p.n23955 0.001
R29671 vp_p.n25378 vp_p.n25377 0.001
R29672 vp_p.n26803 vp_p.n26802 0.001
R29673 vp_p.n12614 vp_p.n12613 0.001
R29674 vp_p.n11176 vp_p.n11175 0.001
R29675 vp_p.n9739 vp_p.n9738 0.001
R29676 vp_p.n993 vp_p.n992 0.001
R29677 vp_p.n2419 vp_p.n2418 0.001
R29678 vp_p.n3844 vp_p.n3843 0.001
R29679 vp_p.n5268 vp_p.n5267 0.001
R29680 vp_p.n6691 vp_p.n6690 0.001
R29681 vp_p.n8113 vp_p.n8112 0.001
R29682 vp_p.n15417 vp_p.n15416 0.001
R29683 vp_p.n16845 vp_p.n16844 0.001
R29684 vp_p.n18272 vp_p.n18271 0.001
R29685 vp_p.n19698 vp_p.n19697 0.001
R29686 vp_p.n21123 vp_p.n21122 0.001
R29687 vp_p.n22547 vp_p.n22546 0.001
R29688 vp_p.n23970 vp_p.n23969 0.001
R29689 vp_p.n25392 vp_p.n25391 0.001
R29690 vp_p.n26817 vp_p.n26816 0.001
R29691 vp_p.n12628 vp_p.n12627 0.001
R29692 vp_p.n11190 vp_p.n11189 0.001
R29693 vp_p.n9753 vp_p.n9752 0.001
R29694 vp_p.n1007 vp_p.n1006 0.001
R29695 vp_p.n2433 vp_p.n2432 0.001
R29696 vp_p.n3858 vp_p.n3857 0.001
R29697 vp_p.n5282 vp_p.n5281 0.001
R29698 vp_p.n6705 vp_p.n6704 0.001
R29699 vp_p.n8127 vp_p.n8126 0.001
R29700 vp_p.n15431 vp_p.n15430 0.001
R29701 vp_p.n16859 vp_p.n16858 0.001
R29702 vp_p.n18286 vp_p.n18285 0.001
R29703 vp_p.n19712 vp_p.n19711 0.001
R29704 vp_p.n21137 vp_p.n21136 0.001
R29705 vp_p.n22561 vp_p.n22560 0.001
R29706 vp_p.n23984 vp_p.n23983 0.001
R29707 vp_p.n25406 vp_p.n25405 0.001
R29708 vp_p.n26831 vp_p.n26830 0.001
R29709 vp_p.n12642 vp_p.n12641 0.001
R29710 vp_p.n11204 vp_p.n11203 0.001
R29711 vp_p.n9767 vp_p.n9766 0.001
R29712 vp_p.n1021 vp_p.n1020 0.001
R29713 vp_p.n2447 vp_p.n2446 0.001
R29714 vp_p.n3872 vp_p.n3871 0.001
R29715 vp_p.n5296 vp_p.n5295 0.001
R29716 vp_p.n6719 vp_p.n6718 0.001
R29717 vp_p.n8141 vp_p.n8140 0.001
R29718 vp_p.n15445 vp_p.n15444 0.001
R29719 vp_p.n16873 vp_p.n16872 0.001
R29720 vp_p.n18300 vp_p.n18299 0.001
R29721 vp_p.n19726 vp_p.n19725 0.001
R29722 vp_p.n21151 vp_p.n21150 0.001
R29723 vp_p.n22575 vp_p.n22574 0.001
R29724 vp_p.n23998 vp_p.n23997 0.001
R29725 vp_p.n25420 vp_p.n25419 0.001
R29726 vp_p.n26845 vp_p.n26844 0.001
R29727 vp_p.n12656 vp_p.n12655 0.001
R29728 vp_p.n11218 vp_p.n11217 0.001
R29729 vp_p.n9781 vp_p.n9780 0.001
R29730 vp_p.n1035 vp_p.n1034 0.001
R29731 vp_p.n2461 vp_p.n2460 0.001
R29732 vp_p.n3886 vp_p.n3885 0.001
R29733 vp_p.n5310 vp_p.n5309 0.001
R29734 vp_p.n6733 vp_p.n6732 0.001
R29735 vp_p.n8155 vp_p.n8154 0.001
R29736 vp_p.n15459 vp_p.n15458 0.001
R29737 vp_p.n16887 vp_p.n16886 0.001
R29738 vp_p.n18314 vp_p.n18313 0.001
R29739 vp_p.n19740 vp_p.n19739 0.001
R29740 vp_p.n21165 vp_p.n21164 0.001
R29741 vp_p.n22589 vp_p.n22588 0.001
R29742 vp_p.n24012 vp_p.n24011 0.001
R29743 vp_p.n25434 vp_p.n25433 0.001
R29744 vp_p.n26859 vp_p.n26858 0.001
R29745 vp_p.n12670 vp_p.n12669 0.001
R29746 vp_p.n11232 vp_p.n11231 0.001
R29747 vp_p.n9795 vp_p.n9794 0.001
R29748 vp_p.n1049 vp_p.n1048 0.001
R29749 vp_p.n2475 vp_p.n2474 0.001
R29750 vp_p.n3900 vp_p.n3899 0.001
R29751 vp_p.n5324 vp_p.n5323 0.001
R29752 vp_p.n6747 vp_p.n6746 0.001
R29753 vp_p.n8169 vp_p.n8168 0.001
R29754 vp_p.n15473 vp_p.n15472 0.001
R29755 vp_p.n16901 vp_p.n16900 0.001
R29756 vp_p.n18328 vp_p.n18327 0.001
R29757 vp_p.n19754 vp_p.n19753 0.001
R29758 vp_p.n21179 vp_p.n21178 0.001
R29759 vp_p.n22603 vp_p.n22602 0.001
R29760 vp_p.n24026 vp_p.n24025 0.001
R29761 vp_p.n25448 vp_p.n25447 0.001
R29762 vp_p.n26873 vp_p.n26872 0.001
R29763 vp_p.n12684 vp_p.n12683 0.001
R29764 vp_p.n11246 vp_p.n11245 0.001
R29765 vp_p.n9809 vp_p.n9808 0.001
R29766 vp_p.n1063 vp_p.n1062 0.001
R29767 vp_p.n2489 vp_p.n2488 0.001
R29768 vp_p.n3914 vp_p.n3913 0.001
R29769 vp_p.n5338 vp_p.n5337 0.001
R29770 vp_p.n6761 vp_p.n6760 0.001
R29771 vp_p.n8183 vp_p.n8182 0.001
R29772 vp_p.n15487 vp_p.n15486 0.001
R29773 vp_p.n16915 vp_p.n16914 0.001
R29774 vp_p.n18342 vp_p.n18341 0.001
R29775 vp_p.n19768 vp_p.n19767 0.001
R29776 vp_p.n21193 vp_p.n21192 0.001
R29777 vp_p.n22617 vp_p.n22616 0.001
R29778 vp_p.n24040 vp_p.n24039 0.001
R29779 vp_p.n25462 vp_p.n25461 0.001
R29780 vp_p.n26887 vp_p.n26886 0.001
R29781 vp_p.n12698 vp_p.n12697 0.001
R29782 vp_p.n11260 vp_p.n11259 0.001
R29783 vp_p.n9823 vp_p.n9822 0.001
R29784 vp_p.n1077 vp_p.n1076 0.001
R29785 vp_p.n2503 vp_p.n2502 0.001
R29786 vp_p.n3928 vp_p.n3927 0.001
R29787 vp_p.n5352 vp_p.n5351 0.001
R29788 vp_p.n6775 vp_p.n6774 0.001
R29789 vp_p.n8197 vp_p.n8196 0.001
R29790 vp_p.n15501 vp_p.n15500 0.001
R29791 vp_p.n16929 vp_p.n16928 0.001
R29792 vp_p.n18356 vp_p.n18355 0.001
R29793 vp_p.n19782 vp_p.n19781 0.001
R29794 vp_p.n21207 vp_p.n21206 0.001
R29795 vp_p.n22631 vp_p.n22630 0.001
R29796 vp_p.n24054 vp_p.n24053 0.001
R29797 vp_p.n25476 vp_p.n25475 0.001
R29798 vp_p.n26901 vp_p.n26900 0.001
R29799 vp_p.n12712 vp_p.n12711 0.001
R29800 vp_p.n11274 vp_p.n11273 0.001
R29801 vp_p.n9837 vp_p.n9836 0.001
R29802 vp_p.n1091 vp_p.n1090 0.001
R29803 vp_p.n2517 vp_p.n2516 0.001
R29804 vp_p.n3942 vp_p.n3941 0.001
R29805 vp_p.n5366 vp_p.n5365 0.001
R29806 vp_p.n6789 vp_p.n6788 0.001
R29807 vp_p.n8211 vp_p.n8210 0.001
R29808 vp_p.n15515 vp_p.n15514 0.001
R29809 vp_p.n16943 vp_p.n16942 0.001
R29810 vp_p.n18370 vp_p.n18369 0.001
R29811 vp_p.n19796 vp_p.n19795 0.001
R29812 vp_p.n21221 vp_p.n21220 0.001
R29813 vp_p.n22645 vp_p.n22644 0.001
R29814 vp_p.n24068 vp_p.n24067 0.001
R29815 vp_p.n25490 vp_p.n25489 0.001
R29816 vp_p.n26915 vp_p.n26914 0.001
R29817 vp_p.n12726 vp_p.n12725 0.001
R29818 vp_p.n11288 vp_p.n11287 0.001
R29819 vp_p.n9851 vp_p.n9850 0.001
R29820 vp_p.n1105 vp_p.n1104 0.001
R29821 vp_p.n2531 vp_p.n2530 0.001
R29822 vp_p.n3956 vp_p.n3955 0.001
R29823 vp_p.n5380 vp_p.n5379 0.001
R29824 vp_p.n6803 vp_p.n6802 0.001
R29825 vp_p.n8225 vp_p.n8224 0.001
R29826 vp_p.n15529 vp_p.n15528 0.001
R29827 vp_p.n16957 vp_p.n16956 0.001
R29828 vp_p.n18384 vp_p.n18383 0.001
R29829 vp_p.n19810 vp_p.n19809 0.001
R29830 vp_p.n21235 vp_p.n21234 0.001
R29831 vp_p.n22659 vp_p.n22658 0.001
R29832 vp_p.n24082 vp_p.n24081 0.001
R29833 vp_p.n25504 vp_p.n25503 0.001
R29834 vp_p.n26929 vp_p.n26928 0.001
R29835 vp_p.n12740 vp_p.n12739 0.001
R29836 vp_p.n11302 vp_p.n11301 0.001
R29837 vp_p.n9865 vp_p.n9864 0.001
R29838 vp_p.n1119 vp_p.n1118 0.001
R29839 vp_p.n2545 vp_p.n2544 0.001
R29840 vp_p.n3970 vp_p.n3969 0.001
R29841 vp_p.n5394 vp_p.n5393 0.001
R29842 vp_p.n6817 vp_p.n6816 0.001
R29843 vp_p.n8239 vp_p.n8238 0.001
R29844 vp_p.n15543 vp_p.n15542 0.001
R29845 vp_p.n16971 vp_p.n16970 0.001
R29846 vp_p.n18398 vp_p.n18397 0.001
R29847 vp_p.n19824 vp_p.n19823 0.001
R29848 vp_p.n21249 vp_p.n21248 0.001
R29849 vp_p.n22673 vp_p.n22672 0.001
R29850 vp_p.n24096 vp_p.n24095 0.001
R29851 vp_p.n25518 vp_p.n25517 0.001
R29852 vp_p.n26943 vp_p.n26942 0.001
R29853 vp_p.n12754 vp_p.n12753 0.001
R29854 vp_p.n11316 vp_p.n11315 0.001
R29855 vp_p.n9879 vp_p.n9878 0.001
R29856 vp_p.n1133 vp_p.n1132 0.001
R29857 vp_p.n2559 vp_p.n2558 0.001
R29858 vp_p.n3984 vp_p.n3983 0.001
R29859 vp_p.n5408 vp_p.n5407 0.001
R29860 vp_p.n6831 vp_p.n6830 0.001
R29861 vp_p.n8253 vp_p.n8252 0.001
R29862 vp_p.n15557 vp_p.n15556 0.001
R29863 vp_p.n16985 vp_p.n16984 0.001
R29864 vp_p.n18412 vp_p.n18411 0.001
R29865 vp_p.n19838 vp_p.n19837 0.001
R29866 vp_p.n21263 vp_p.n21262 0.001
R29867 vp_p.n22687 vp_p.n22686 0.001
R29868 vp_p.n24110 vp_p.n24109 0.001
R29869 vp_p.n25532 vp_p.n25531 0.001
R29870 vp_p.n26957 vp_p.n26956 0.001
R29871 vp_p.n12768 vp_p.n12767 0.001
R29872 vp_p.n11330 vp_p.n11329 0.001
R29873 vp_p.n9893 vp_p.n9892 0.001
R29874 vp_p.n1147 vp_p.n1146 0.001
R29875 vp_p.n2573 vp_p.n2572 0.001
R29876 vp_p.n3998 vp_p.n3997 0.001
R29877 vp_p.n5422 vp_p.n5421 0.001
R29878 vp_p.n6845 vp_p.n6844 0.001
R29879 vp_p.n8267 vp_p.n8266 0.001
R29880 vp_p.n15571 vp_p.n15570 0.001
R29881 vp_p.n16999 vp_p.n16998 0.001
R29882 vp_p.n18426 vp_p.n18425 0.001
R29883 vp_p.n19852 vp_p.n19851 0.001
R29884 vp_p.n21277 vp_p.n21276 0.001
R29885 vp_p.n22701 vp_p.n22700 0.001
R29886 vp_p.n24124 vp_p.n24123 0.001
R29887 vp_p.n25546 vp_p.n25545 0.001
R29888 vp_p.n26971 vp_p.n26970 0.001
R29889 vp_p.n12782 vp_p.n12781 0.001
R29890 vp_p.n11344 vp_p.n11343 0.001
R29891 vp_p.n9907 vp_p.n9906 0.001
R29892 vp_p.n1161 vp_p.n1160 0.001
R29893 vp_p.n2587 vp_p.n2586 0.001
R29894 vp_p.n4012 vp_p.n4011 0.001
R29895 vp_p.n5436 vp_p.n5435 0.001
R29896 vp_p.n6859 vp_p.n6858 0.001
R29897 vp_p.n8281 vp_p.n8280 0.001
R29898 vp_p.n15585 vp_p.n15584 0.001
R29899 vp_p.n17013 vp_p.n17012 0.001
R29900 vp_p.n18440 vp_p.n18439 0.001
R29901 vp_p.n19866 vp_p.n19865 0.001
R29902 vp_p.n21291 vp_p.n21290 0.001
R29903 vp_p.n22715 vp_p.n22714 0.001
R29904 vp_p.n24138 vp_p.n24137 0.001
R29905 vp_p.n25560 vp_p.n25559 0.001
R29906 vp_p.n26985 vp_p.n26984 0.001
R29907 vp_p.n12796 vp_p.n12795 0.001
R29908 vp_p.n11358 vp_p.n11357 0.001
R29909 vp_p.n9921 vp_p.n9920 0.001
R29910 vp_p.n1175 vp_p.n1174 0.001
R29911 vp_p.n2601 vp_p.n2600 0.001
R29912 vp_p.n4026 vp_p.n4025 0.001
R29913 vp_p.n5450 vp_p.n5449 0.001
R29914 vp_p.n6873 vp_p.n6872 0.001
R29915 vp_p.n8295 vp_p.n8294 0.001
R29916 vp_p.n15599 vp_p.n15598 0.001
R29917 vp_p.n17027 vp_p.n17026 0.001
R29918 vp_p.n18454 vp_p.n18453 0.001
R29919 vp_p.n19880 vp_p.n19879 0.001
R29920 vp_p.n21305 vp_p.n21304 0.001
R29921 vp_p.n22729 vp_p.n22728 0.001
R29922 vp_p.n24152 vp_p.n24151 0.001
R29923 vp_p.n25574 vp_p.n25573 0.001
R29924 vp_p.n26999 vp_p.n26998 0.001
R29925 vp_p.n12810 vp_p.n12809 0.001
R29926 vp_p.n11372 vp_p.n11371 0.001
R29927 vp_p.n9935 vp_p.n9934 0.001
R29928 vp_p.n1189 vp_p.n1188 0.001
R29929 vp_p.n2615 vp_p.n2614 0.001
R29930 vp_p.n4040 vp_p.n4039 0.001
R29931 vp_p.n5464 vp_p.n5463 0.001
R29932 vp_p.n6887 vp_p.n6886 0.001
R29933 vp_p.n8309 vp_p.n8308 0.001
R29934 vp_p.n15613 vp_p.n15612 0.001
R29935 vp_p.n17041 vp_p.n17040 0.001
R29936 vp_p.n18468 vp_p.n18467 0.001
R29937 vp_p.n19894 vp_p.n19893 0.001
R29938 vp_p.n21319 vp_p.n21318 0.001
R29939 vp_p.n22743 vp_p.n22742 0.001
R29940 vp_p.n24166 vp_p.n24165 0.001
R29941 vp_p.n25588 vp_p.n25587 0.001
R29942 vp_p.n27013 vp_p.n27012 0.001
R29943 vp_p.n12824 vp_p.n12823 0.001
R29944 vp_p.n11386 vp_p.n11385 0.001
R29945 vp_p.n9949 vp_p.n9948 0.001
R29946 vp_p.n1203 vp_p.n1202 0.001
R29947 vp_p.n2629 vp_p.n2628 0.001
R29948 vp_p.n4054 vp_p.n4053 0.001
R29949 vp_p.n5478 vp_p.n5477 0.001
R29950 vp_p.n6901 vp_p.n6900 0.001
R29951 vp_p.n8323 vp_p.n8322 0.001
R29952 vp_p.n15627 vp_p.n15626 0.001
R29953 vp_p.n17055 vp_p.n17054 0.001
R29954 vp_p.n18482 vp_p.n18481 0.001
R29955 vp_p.n19908 vp_p.n19907 0.001
R29956 vp_p.n21333 vp_p.n21332 0.001
R29957 vp_p.n22757 vp_p.n22756 0.001
R29958 vp_p.n24180 vp_p.n24179 0.001
R29959 vp_p.n25602 vp_p.n25601 0.001
R29960 vp_p.n27027 vp_p.n27026 0.001
R29961 vp_p.n12838 vp_p.n12837 0.001
R29962 vp_p.n11400 vp_p.n11399 0.001
R29963 vp_p.n9963 vp_p.n9962 0.001
R29964 vp_p.n1217 vp_p.n1216 0.001
R29965 vp_p.n2643 vp_p.n2642 0.001
R29966 vp_p.n4068 vp_p.n4067 0.001
R29967 vp_p.n5492 vp_p.n5491 0.001
R29968 vp_p.n6915 vp_p.n6914 0.001
R29969 vp_p.n8337 vp_p.n8336 0.001
R29970 vp_p.n15641 vp_p.n15640 0.001
R29971 vp_p.n17069 vp_p.n17068 0.001
R29972 vp_p.n18496 vp_p.n18495 0.001
R29973 vp_p.n19922 vp_p.n19921 0.001
R29974 vp_p.n21347 vp_p.n21346 0.001
R29975 vp_p.n22771 vp_p.n22770 0.001
R29976 vp_p.n24194 vp_p.n24193 0.001
R29977 vp_p.n25616 vp_p.n25615 0.001
R29978 vp_p.n27041 vp_p.n27040 0.001
R29979 vp_p.n12852 vp_p.n12851 0.001
R29980 vp_p.n11414 vp_p.n11413 0.001
R29981 vp_p.n9977 vp_p.n9976 0.001
R29982 vp_p.n1231 vp_p.n1230 0.001
R29983 vp_p.n2657 vp_p.n2656 0.001
R29984 vp_p.n4082 vp_p.n4081 0.001
R29985 vp_p.n5506 vp_p.n5505 0.001
R29986 vp_p.n6929 vp_p.n6928 0.001
R29987 vp_p.n8351 vp_p.n8350 0.001
R29988 vp_p.n15655 vp_p.n15654 0.001
R29989 vp_p.n17083 vp_p.n17082 0.001
R29990 vp_p.n18510 vp_p.n18509 0.001
R29991 vp_p.n19936 vp_p.n19935 0.001
R29992 vp_p.n21361 vp_p.n21360 0.001
R29993 vp_p.n22785 vp_p.n22784 0.001
R29994 vp_p.n24208 vp_p.n24207 0.001
R29995 vp_p.n25630 vp_p.n25629 0.001
R29996 vp_p.n27055 vp_p.n27054 0.001
R29997 vp_p.n12866 vp_p.n12865 0.001
R29998 vp_p.n11428 vp_p.n11427 0.001
R29999 vp_p.n9991 vp_p.n9990 0.001
R30000 vp_p.n1245 vp_p.n1244 0.001
R30001 vp_p.n2671 vp_p.n2670 0.001
R30002 vp_p.n4096 vp_p.n4095 0.001
R30003 vp_p.n5520 vp_p.n5519 0.001
R30004 vp_p.n6943 vp_p.n6942 0.001
R30005 vp_p.n8365 vp_p.n8364 0.001
R30006 vp_p.n15669 vp_p.n15668 0.001
R30007 vp_p.n17097 vp_p.n17096 0.001
R30008 vp_p.n18524 vp_p.n18523 0.001
R30009 vp_p.n19950 vp_p.n19949 0.001
R30010 vp_p.n21375 vp_p.n21374 0.001
R30011 vp_p.n22799 vp_p.n22798 0.001
R30012 vp_p.n24222 vp_p.n24221 0.001
R30013 vp_p.n25644 vp_p.n25643 0.001
R30014 vp_p.n27069 vp_p.n27068 0.001
R30015 vp_p.n12880 vp_p.n12879 0.001
R30016 vp_p.n11442 vp_p.n11441 0.001
R30017 vp_p.n10005 vp_p.n10004 0.001
R30018 vp_p.n1259 vp_p.n1258 0.001
R30019 vp_p.n2685 vp_p.n2684 0.001
R30020 vp_p.n4110 vp_p.n4109 0.001
R30021 vp_p.n5534 vp_p.n5533 0.001
R30022 vp_p.n6957 vp_p.n6956 0.001
R30023 vp_p.n8379 vp_p.n8378 0.001
R30024 vp_p.n15683 vp_p.n15682 0.001
R30025 vp_p.n17111 vp_p.n17110 0.001
R30026 vp_p.n18538 vp_p.n18537 0.001
R30027 vp_p.n19964 vp_p.n19963 0.001
R30028 vp_p.n21389 vp_p.n21388 0.001
R30029 vp_p.n22813 vp_p.n22812 0.001
R30030 vp_p.n24236 vp_p.n24235 0.001
R30031 vp_p.n25658 vp_p.n25657 0.001
R30032 vp_p.n27083 vp_p.n27082 0.001
R30033 vp_p.n12894 vp_p.n12893 0.001
R30034 vp_p.n11456 vp_p.n11455 0.001
R30035 vp_p.n10019 vp_p.n10018 0.001
R30036 vp_p.n1273 vp_p.n1272 0.001
R30037 vp_p.n2699 vp_p.n2698 0.001
R30038 vp_p.n4124 vp_p.n4123 0.001
R30039 vp_p.n5548 vp_p.n5547 0.001
R30040 vp_p.n6971 vp_p.n6970 0.001
R30041 vp_p.n8393 vp_p.n8392 0.001
R30042 vp_p.n15697 vp_p.n15696 0.001
R30043 vp_p.n17125 vp_p.n17124 0.001
R30044 vp_p.n18552 vp_p.n18551 0.001
R30045 vp_p.n19978 vp_p.n19977 0.001
R30046 vp_p.n21403 vp_p.n21402 0.001
R30047 vp_p.n22827 vp_p.n22826 0.001
R30048 vp_p.n24250 vp_p.n24249 0.001
R30049 vp_p.n25672 vp_p.n25671 0.001
R30050 vp_p.n27097 vp_p.n27096 0.001
R30051 vp_p.n12908 vp_p.n12907 0.001
R30052 vp_p.n11470 vp_p.n11469 0.001
R30053 vp_p.n10033 vp_p.n10032 0.001
R30054 vp_p.n1287 vp_p.n1286 0.001
R30055 vp_p.n2713 vp_p.n2712 0.001
R30056 vp_p.n4138 vp_p.n4137 0.001
R30057 vp_p.n5562 vp_p.n5561 0.001
R30058 vp_p.n6985 vp_p.n6984 0.001
R30059 vp_p.n8407 vp_p.n8406 0.001
R30060 vp_p.n15711 vp_p.n15710 0.001
R30061 vp_p.n17139 vp_p.n17138 0.001
R30062 vp_p.n18566 vp_p.n18565 0.001
R30063 vp_p.n19992 vp_p.n19991 0.001
R30064 vp_p.n21417 vp_p.n21416 0.001
R30065 vp_p.n22841 vp_p.n22840 0.001
R30066 vp_p.n24264 vp_p.n24263 0.001
R30067 vp_p.n25686 vp_p.n25685 0.001
R30068 vp_p.n27111 vp_p.n27110 0.001
R30069 vp_p.n12922 vp_p.n12921 0.001
R30070 vp_p.n11484 vp_p.n11483 0.001
R30071 vp_p.n10047 vp_p.n10046 0.001
R30072 vp_p.n1301 vp_p.n1300 0.001
R30073 vp_p.n2727 vp_p.n2726 0.001
R30074 vp_p.n4152 vp_p.n4151 0.001
R30075 vp_p.n5576 vp_p.n5575 0.001
R30076 vp_p.n6999 vp_p.n6998 0.001
R30077 vp_p.n8421 vp_p.n8420 0.001
R30078 vp_p.n15725 vp_p.n15724 0.001
R30079 vp_p.n17153 vp_p.n17152 0.001
R30080 vp_p.n18580 vp_p.n18579 0.001
R30081 vp_p.n20006 vp_p.n20005 0.001
R30082 vp_p.n21431 vp_p.n21430 0.001
R30083 vp_p.n22855 vp_p.n22854 0.001
R30084 vp_p.n24278 vp_p.n24277 0.001
R30085 vp_p.n25700 vp_p.n25699 0.001
R30086 vp_p.n27125 vp_p.n27124 0.001
R30087 vp_p.n12936 vp_p.n12935 0.001
R30088 vp_p.n11498 vp_p.n11497 0.001
R30089 vp_p.n10061 vp_p.n10060 0.001
R30090 vp_p.n1315 vp_p.n1314 0.001
R30091 vp_p.n2741 vp_p.n2740 0.001
R30092 vp_p.n4166 vp_p.n4165 0.001
R30093 vp_p.n5590 vp_p.n5589 0.001
R30094 vp_p.n7013 vp_p.n7012 0.001
R30095 vp_p.n8435 vp_p.n8434 0.001
R30096 vp_p.n15739 vp_p.n15738 0.001
R30097 vp_p.n17167 vp_p.n17166 0.001
R30098 vp_p.n18594 vp_p.n18593 0.001
R30099 vp_p.n20020 vp_p.n20019 0.001
R30100 vp_p.n21445 vp_p.n21444 0.001
R30101 vp_p.n22869 vp_p.n22868 0.001
R30102 vp_p.n24292 vp_p.n24291 0.001
R30103 vp_p.n25714 vp_p.n25713 0.001
R30104 vp_p.n27139 vp_p.n27138 0.001
R30105 vp_p.n12950 vp_p.n12949 0.001
R30106 vp_p.n11512 vp_p.n11511 0.001
R30107 vp_p.n10075 vp_p.n10074 0.001
R30108 vp_p.n1329 vp_p.n1328 0.001
R30109 vp_p.n2755 vp_p.n2754 0.001
R30110 vp_p.n4180 vp_p.n4179 0.001
R30111 vp_p.n5604 vp_p.n5603 0.001
R30112 vp_p.n7027 vp_p.n7026 0.001
R30113 vp_p.n8449 vp_p.n8448 0.001
R30114 vp_p.n15753 vp_p.n15752 0.001
R30115 vp_p.n17181 vp_p.n17180 0.001
R30116 vp_p.n18608 vp_p.n18607 0.001
R30117 vp_p.n20034 vp_p.n20033 0.001
R30118 vp_p.n21459 vp_p.n21458 0.001
R30119 vp_p.n22883 vp_p.n22882 0.001
R30120 vp_p.n24306 vp_p.n24305 0.001
R30121 vp_p.n25728 vp_p.n25727 0.001
R30122 vp_p.n27153 vp_p.n27152 0.001
R30123 vp_p.n12964 vp_p.n12963 0.001
R30124 vp_p.n11526 vp_p.n11525 0.001
R30125 vp_p.n10089 vp_p.n10088 0.001
R30126 vp_p.n1343 vp_p.n1342 0.001
R30127 vp_p.n2769 vp_p.n2768 0.001
R30128 vp_p.n4194 vp_p.n4193 0.001
R30129 vp_p.n5618 vp_p.n5617 0.001
R30130 vp_p.n7041 vp_p.n7040 0.001
R30131 vp_p.n8463 vp_p.n8462 0.001
R30132 vp_p.n15767 vp_p.n15766 0.001
R30133 vp_p.n17195 vp_p.n17194 0.001
R30134 vp_p.n18622 vp_p.n18621 0.001
R30135 vp_p.n20048 vp_p.n20047 0.001
R30136 vp_p.n21473 vp_p.n21472 0.001
R30137 vp_p.n22897 vp_p.n22896 0.001
R30138 vp_p.n24320 vp_p.n24319 0.001
R30139 vp_p.n25742 vp_p.n25741 0.001
R30140 vp_p.n27167 vp_p.n27166 0.001
R30141 vp_p.n12978 vp_p.n12977 0.001
R30142 vp_p.n11540 vp_p.n11539 0.001
R30143 vp_p.n10103 vp_p.n10102 0.001
R30144 vp_p.n1357 vp_p.n1356 0.001
R30145 vp_p.n2783 vp_p.n2782 0.001
R30146 vp_p.n4208 vp_p.n4207 0.001
R30147 vp_p.n5632 vp_p.n5631 0.001
R30148 vp_p.n7055 vp_p.n7054 0.001
R30149 vp_p.n8477 vp_p.n8476 0.001
R30150 vp_p.n15781 vp_p.n15780 0.001
R30151 vp_p.n17209 vp_p.n17208 0.001
R30152 vp_p.n18636 vp_p.n18635 0.001
R30153 vp_p.n20062 vp_p.n20061 0.001
R30154 vp_p.n21487 vp_p.n21486 0.001
R30155 vp_p.n22911 vp_p.n22910 0.001
R30156 vp_p.n24334 vp_p.n24333 0.001
R30157 vp_p.n25756 vp_p.n25755 0.001
R30158 vp_p.n27181 vp_p.n27180 0.001
R30159 vp_p.n12992 vp_p.n12991 0.001
R30160 vp_p.n11554 vp_p.n11553 0.001
R30161 vp_p.n10117 vp_p.n10116 0.001
R30162 vp_p.n1371 vp_p.n1370 0.001
R30163 vp_p.n2797 vp_p.n2796 0.001
R30164 vp_p.n4222 vp_p.n4221 0.001
R30165 vp_p.n5646 vp_p.n5645 0.001
R30166 vp_p.n7069 vp_p.n7068 0.001
R30167 vp_p.n8491 vp_p.n8490 0.001
R30168 vp_p.n15795 vp_p.n15794 0.001
R30169 vp_p.n17223 vp_p.n17222 0.001
R30170 vp_p.n18650 vp_p.n18649 0.001
R30171 vp_p.n20076 vp_p.n20075 0.001
R30172 vp_p.n21501 vp_p.n21500 0.001
R30173 vp_p.n22925 vp_p.n22924 0.001
R30174 vp_p.n24348 vp_p.n24347 0.001
R30175 vp_p.n25770 vp_p.n25769 0.001
R30176 vp_p.n27195 vp_p.n27194 0.001
R30177 vp_p.n13006 vp_p.n13005 0.001
R30178 vp_p.n11568 vp_p.n11567 0.001
R30179 vp_p.n10131 vp_p.n10130 0.001
R30180 vp_p.n1385 vp_p.n1384 0.001
R30181 vp_p.n2811 vp_p.n2810 0.001
R30182 vp_p.n4236 vp_p.n4235 0.001
R30183 vp_p.n5660 vp_p.n5659 0.001
R30184 vp_p.n7083 vp_p.n7082 0.001
R30185 vp_p.n8505 vp_p.n8504 0.001
R30186 vp_p.n15809 vp_p.n15808 0.001
R30187 vp_p.n17237 vp_p.n17236 0.001
R30188 vp_p.n18664 vp_p.n18663 0.001
R30189 vp_p.n20090 vp_p.n20089 0.001
R30190 vp_p.n21515 vp_p.n21514 0.001
R30191 vp_p.n22939 vp_p.n22938 0.001
R30192 vp_p.n24362 vp_p.n24361 0.001
R30193 vp_p.n25784 vp_p.n25783 0.001
R30194 vp_p.n27209 vp_p.n27208 0.001
R30195 vp_p.n11582 vp_p.n11581 0.001
R30196 vp_p.n10145 vp_p.n10144 0.001
R30197 vp_p.n1399 vp_p.n1398 0.001
R30198 vp_p.n2825 vp_p.n2824 0.001
R30199 vp_p.n4250 vp_p.n4249 0.001
R30200 vp_p.n5674 vp_p.n5673 0.001
R30201 vp_p.n7097 vp_p.n7096 0.001
R30202 vp_p.n8519 vp_p.n8518 0.001
R30203 vp_p.n17251 vp_p.n17250 0.001
R30204 vp_p.n18678 vp_p.n18677 0.001
R30205 vp_p.n20104 vp_p.n20103 0.001
R30206 vp_p.n21529 vp_p.n21528 0.001
R30207 vp_p.n22953 vp_p.n22952 0.001
R30208 vp_p.n24376 vp_p.n24375 0.001
R30209 vp_p.n25798 vp_p.n25797 0.001
R30210 vp_p.n27223 vp_p.n27222 0.001
R30211 vp_p.n10159 vp_p.n10158 0.001
R30212 vp_p.n1413 vp_p.n1412 0.001
R30213 vp_p.n2839 vp_p.n2838 0.001
R30214 vp_p.n4264 vp_p.n4263 0.001
R30215 vp_p.n5688 vp_p.n5687 0.001
R30216 vp_p.n7111 vp_p.n7110 0.001
R30217 vp_p.n8533 vp_p.n8532 0.001
R30218 vp_p.n18692 vp_p.n18691 0.001
R30219 vp_p.n20118 vp_p.n20117 0.001
R30220 vp_p.n21543 vp_p.n21542 0.001
R30221 vp_p.n22967 vp_p.n22966 0.001
R30222 vp_p.n24390 vp_p.n24389 0.001
R30223 vp_p.n25812 vp_p.n25811 0.001
R30224 vp_p.n27237 vp_p.n27236 0.001
R30225 vp_p.n1427 vp_p.n1426 0.001
R30226 vp_p.n2853 vp_p.n2852 0.001
R30227 vp_p.n4278 vp_p.n4277 0.001
R30228 vp_p.n5702 vp_p.n5701 0.001
R30229 vp_p.n7125 vp_p.n7124 0.001
R30230 vp_p.n8547 vp_p.n8546 0.001
R30231 vp_p.n20132 vp_p.n20131 0.001
R30232 vp_p.n21557 vp_p.n21556 0.001
R30233 vp_p.n22981 vp_p.n22980 0.001
R30234 vp_p.n24404 vp_p.n24403 0.001
R30235 vp_p.n25826 vp_p.n25825 0.001
R30236 vp_p.n27251 vp_p.n27250 0.001
R30237 vp_p.n2867 vp_p.n2866 0.001
R30238 vp_p.n4292 vp_p.n4291 0.001
R30239 vp_p.n5716 vp_p.n5715 0.001
R30240 vp_p.n7139 vp_p.n7138 0.001
R30241 vp_p.n8561 vp_p.n8560 0.001
R30242 vp_p.n21571 vp_p.n21570 0.001
R30243 vp_p.n22995 vp_p.n22994 0.001
R30244 vp_p.n24418 vp_p.n24417 0.001
R30245 vp_p.n25840 vp_p.n25839 0.001
R30246 vp_p.n27265 vp_p.n27264 0.001
R30247 vp_p.n4306 vp_p.n4305 0.001
R30248 vp_p.n5730 vp_p.n5729 0.001
R30249 vp_p.n7153 vp_p.n7152 0.001
R30250 vp_p.n8575 vp_p.n8574 0.001
R30251 vp_p.n23009 vp_p.n23008 0.001
R30252 vp_p.n24432 vp_p.n24431 0.001
R30253 vp_p.n25854 vp_p.n25853 0.001
R30254 vp_p.n27279 vp_p.n27278 0.001
R30255 vp_p.n5744 vp_p.n5743 0.001
R30256 vp_p.n7167 vp_p.n7166 0.001
R30257 vp_p.n8589 vp_p.n8588 0.001
R30258 vp_p.n24446 vp_p.n24445 0.001
R30259 vp_p.n25868 vp_p.n25867 0.001
R30260 vp_p.n27293 vp_p.n27292 0.001
R30261 vp_p.n7181 vp_p.n7180 0.001
R30262 vp_p.n8603 vp_p.n8602 0.001
R30263 vp_p.n25882 vp_p.n25881 0.001
R30264 vp_p.n27307 vp_p.n27306 0.001
R30265 vp_p.n8617 vp_p.n8616 0.001
R30266 vp_p.n27321 vp_p.n27320 0.001
R30267 vp_p.n14464 vp_p.n13102 0.001
R30268 vp_p.n14459 vp_p.n13107 0.001
R30269 vp_p.n14454 vp_p.n13112 0.001
R30270 vp_p.n14449 vp_p.n13117 0.001
R30271 vp_p.n14444 vp_p.n13122 0.001
R30272 vp_p.n14439 vp_p.n13127 0.001
R30273 vp_p.n14434 vp_p.n13132 0.001
R30274 vp_p.n14429 vp_p.n13137 0.001
R30275 vp_p.n14424 vp_p.n13142 0.001
R30276 vp_p.n14419 vp_p.n13147 0.001
R30277 vp_p.n14414 vp_p.n13152 0.001
R30278 vp_p.n14409 vp_p.n13157 0.001
R30279 vp_p.n14404 vp_p.n13162 0.001
R30280 vp_p.n14399 vp_p.n13167 0.001
R30281 vp_p.n14394 vp_p.n13172 0.001
R30282 vp_p.n14389 vp_p.n13177 0.001
R30283 vp_p.n13850 vp_p.n13837 0.001
R30284 vp_p.n13845 vp_p.n13842 0.001
R30285 vp_p.n13095 vp_p.n11668 0.001
R30286 vp_p.n13090 vp_p.n11673 0.001
R30287 vp_p.n13085 vp_p.n11678 0.001
R30288 vp_p.n13080 vp_p.n11683 0.001
R30289 vp_p.n13075 vp_p.n11688 0.001
R30290 vp_p.n13070 vp_p.n11693 0.001
R30291 vp_p.n13065 vp_p.n11698 0.001
R30292 vp_p.n13060 vp_p.n11703 0.001
R30293 vp_p.n13055 vp_p.n11708 0.001
R30294 vp_p.n13050 vp_p.n11713 0.001
R30295 vp_p.n13045 vp_p.n11718 0.001
R30296 vp_p.n13040 vp_p.n11723 0.001
R30297 vp_p.n13035 vp_p.n11728 0.001
R30298 vp_p.n13030 vp_p.n11733 0.001
R30299 vp_p.n13025 vp_p.n11738 0.001
R30300 vp_p.n12086 vp_p.n12073 0.001
R30301 vp_p.n12081 vp_p.n12078 0.001
R30302 vp_p.n15897 vp_p.n14471 0.001
R30303 vp_p.n15892 vp_p.n14476 0.001
R30304 vp_p.n15887 vp_p.n14481 0.001
R30305 vp_p.n15882 vp_p.n14486 0.001
R30306 vp_p.n15877 vp_p.n14491 0.001
R30307 vp_p.n15872 vp_p.n14496 0.001
R30308 vp_p.n15867 vp_p.n14501 0.001
R30309 vp_p.n15862 vp_p.n14506 0.001
R30310 vp_p.n15857 vp_p.n14511 0.001
R30311 vp_p.n15852 vp_p.n14516 0.001
R30312 vp_p.n15847 vp_p.n14521 0.001
R30313 vp_p.n15842 vp_p.n14526 0.001
R30314 vp_p.n15837 vp_p.n14531 0.001
R30315 vp_p.n15832 vp_p.n14536 0.001
R30316 vp_p.n14889 vp_p.n14876 0.001
R30317 vp_p.n14884 vp_p.n14881 0.001
R30318 vp_p.n11661 vp_p.n10235 0.001
R30319 vp_p.n11656 vp_p.n10240 0.001
R30320 vp_p.n11651 vp_p.n10245 0.001
R30321 vp_p.n11646 vp_p.n10250 0.001
R30322 vp_p.n11641 vp_p.n10255 0.001
R30323 vp_p.n11636 vp_p.n10260 0.001
R30324 vp_p.n11631 vp_p.n10265 0.001
R30325 vp_p.n11626 vp_p.n10270 0.001
R30326 vp_p.n11621 vp_p.n10275 0.001
R30327 vp_p.n11616 vp_p.n10280 0.001
R30328 vp_p.n11611 vp_p.n10285 0.001
R30329 vp_p.n11606 vp_p.n10290 0.001
R30330 vp_p.n11601 vp_p.n10295 0.001
R30331 vp_p.n10648 vp_p.n10635 0.001
R30332 vp_p.n10643 vp_p.n10640 0.001
R30333 vp_p.n17329 vp_p.n15904 0.001
R30334 vp_p.n17324 vp_p.n15909 0.001
R30335 vp_p.n17319 vp_p.n15914 0.001
R30336 vp_p.n17314 vp_p.n15919 0.001
R30337 vp_p.n17309 vp_p.n15924 0.001
R30338 vp_p.n17304 vp_p.n15929 0.001
R30339 vp_p.n17299 vp_p.n15934 0.001
R30340 vp_p.n17294 vp_p.n15939 0.001
R30341 vp_p.n17289 vp_p.n15944 0.001
R30342 vp_p.n17284 vp_p.n15949 0.001
R30343 vp_p.n17279 vp_p.n15954 0.001
R30344 vp_p.n17274 vp_p.n15959 0.001
R30345 vp_p.n16317 vp_p.n16304 0.001
R30346 vp_p.n16312 vp_p.n16309 0.001
R30347 vp_p.n10228 vp_p.n8738 0.001
R30348 vp_p.n10223 vp_p.n8743 0.001
R30349 vp_p.n10218 vp_p.n8748 0.001
R30350 vp_p.n10213 vp_p.n8753 0.001
R30351 vp_p.n10208 vp_p.n8758 0.001
R30352 vp_p.n10203 vp_p.n8763 0.001
R30353 vp_p.n10198 vp_p.n8768 0.001
R30354 vp_p.n10193 vp_p.n8773 0.001
R30355 vp_p.n10188 vp_p.n8778 0.001
R30356 vp_p.n10183 vp_p.n8783 0.001
R30357 vp_p.n10178 vp_p.n8788 0.001
R30358 vp_p.n9211 vp_p.n9133 0.001
R30359 vp_p.n9206 vp_p.n9138 0.001
R30360 vp_p.n18760 vp_p.n17336 0.001
R30361 vp_p.n18755 vp_p.n17341 0.001
R30362 vp_p.n18750 vp_p.n17346 0.001
R30363 vp_p.n18745 vp_p.n17351 0.001
R30364 vp_p.n18740 vp_p.n17356 0.001
R30365 vp_p.n18735 vp_p.n17361 0.001
R30366 vp_p.n18730 vp_p.n17366 0.001
R30367 vp_p.n18725 vp_p.n17371 0.001
R30368 vp_p.n18720 vp_p.n17376 0.001
R30369 vp_p.n18715 vp_p.n17381 0.001
R30370 vp_p.n17744 vp_p.n17731 0.001
R30371 vp_p.n17739 vp_p.n17736 0.001
R30372 vp_p.n1486 vp_p.n4 0.001
R30373 vp_p.n1481 vp_p.n9 0.001
R30374 vp_p.n1476 vp_p.n14 0.001
R30375 vp_p.n1471 vp_p.n19 0.001
R30376 vp_p.n1466 vp_p.n24 0.001
R30377 vp_p.n1461 vp_p.n29 0.001
R30378 vp_p.n1456 vp_p.n34 0.001
R30379 vp_p.n1451 vp_p.n39 0.001
R30380 vp_p.n1446 vp_p.n44 0.001
R30381 vp_p.n465 vp_p.n394 0.001
R30382 vp_p.n460 vp_p.n399 0.001
R30383 vp_p.n20190 vp_p.n18767 0.001
R30384 vp_p.n20185 vp_p.n18772 0.001
R30385 vp_p.n20180 vp_p.n18777 0.001
R30386 vp_p.n20175 vp_p.n18782 0.001
R30387 vp_p.n20170 vp_p.n18787 0.001
R30388 vp_p.n20165 vp_p.n18792 0.001
R30389 vp_p.n20160 vp_p.n18797 0.001
R30390 vp_p.n20155 vp_p.n18802 0.001
R30391 vp_p.n19170 vp_p.n19157 0.001
R30392 vp_p.n19165 vp_p.n19162 0.001
R30393 vp_p.n2916 vp_p.n1493 0.001
R30394 vp_p.n2911 vp_p.n1498 0.001
R30395 vp_p.n2906 vp_p.n1503 0.001
R30396 vp_p.n2901 vp_p.n1508 0.001
R30397 vp_p.n2896 vp_p.n1513 0.001
R30398 vp_p.n2891 vp_p.n1518 0.001
R30399 vp_p.n2886 vp_p.n1523 0.001
R30400 vp_p.n1891 vp_p.n1878 0.001
R30401 vp_p.n1886 vp_p.n1883 0.001
R30402 vp_p.n21619 vp_p.n20197 0.001
R30403 vp_p.n21614 vp_p.n20202 0.001
R30404 vp_p.n21609 vp_p.n20207 0.001
R30405 vp_p.n21604 vp_p.n20212 0.001
R30406 vp_p.n21599 vp_p.n20217 0.001
R30407 vp_p.n21594 vp_p.n20222 0.001
R30408 vp_p.n20595 vp_p.n20582 0.001
R30409 vp_p.n20590 vp_p.n20587 0.001
R30410 vp_p.n4345 vp_p.n2923 0.001
R30411 vp_p.n4340 vp_p.n2928 0.001
R30412 vp_p.n4335 vp_p.n2933 0.001
R30413 vp_p.n4330 vp_p.n2938 0.001
R30414 vp_p.n4325 vp_p.n2943 0.001
R30415 vp_p.n3316 vp_p.n3303 0.001
R30416 vp_p.n3311 vp_p.n3308 0.001
R30417 vp_p.n23047 vp_p.n21626 0.001
R30418 vp_p.n23042 vp_p.n21631 0.001
R30419 vp_p.n23037 vp_p.n21636 0.001
R30420 vp_p.n23032 vp_p.n21641 0.001
R30421 vp_p.n22019 vp_p.n22006 0.001
R30422 vp_p.n22014 vp_p.n22011 0.001
R30423 vp_p.n5773 vp_p.n4352 0.001
R30424 vp_p.n5768 vp_p.n4357 0.001
R30425 vp_p.n5763 vp_p.n4362 0.001
R30426 vp_p.n4740 vp_p.n4727 0.001
R30427 vp_p.n4735 vp_p.n4732 0.001
R30428 vp_p.n24474 vp_p.n23054 0.001
R30429 vp_p.n24469 vp_p.n23059 0.001
R30430 vp_p.n23442 vp_p.n23429 0.001
R30431 vp_p.n23437 vp_p.n23434 0.001
R30432 vp_p.n7200 vp_p.n5780 0.001
R30433 vp_p.n6163 vp_p.n6150 0.001
R30434 vp_p.n6158 vp_p.n6155 0.001
R30435 vp_p.n24864 vp_p.n24851 0.001
R30436 vp_p.n24859 vp_p.n24856 0.001
R30437 vp_p.n7575 vp_p.n7572 0.001
R30438 vp_p.n8627 vp_p.n8626 0.001
R30439 out_p.n768 out_p.t1615 7.173
R30440 out_p.n768 out_p.t1035 7.173
R30441 out_p.n767 out_p.t1773 7.173
R30442 out_p.n767 out_p.t2760 7.173
R30443 out_p.n766 out_p.t2277 7.173
R30444 out_p.n766 out_p.t2997 7.173
R30445 out_p.n765 out_p.t1037 7.173
R30446 out_p.n765 out_p.t2154 7.173
R30447 out_p.n764 out_p.t558 7.173
R30448 out_p.n764 out_p.t2081 7.173
R30449 out_p.n763 out_p.t3001 7.173
R30450 out_p.n763 out_p.t497 7.173
R30451 out_p.n762 out_p.t2157 7.173
R30452 out_p.n762 out_p.t2943 7.173
R30453 out_p.n761 out_p.t3195 7.173
R30454 out_p.n761 out_p.t2197 7.173
R30455 out_p.n760 out_p.t1599 7.173
R30456 out_p.n760 out_p.t1049 7.173
R30457 out_p.n759 out_p.t2461 7.173
R30458 out_p.n759 out_p.t2641 7.173
R30459 out_p.n758 out_p.t1619 7.173
R30460 out_p.n758 out_p.t902 7.173
R30461 out_p.n757 out_p.t2742 7.173
R30462 out_p.n757 out_p.t2004 7.173
R30463 out_p.n756 out_p.t3213 7.173
R30464 out_p.n756 out_p.t2280 7.173
R30465 out_p.n755 out_p.t766 7.173
R30466 out_p.n755 out_p.t3418 7.173
R30467 out_p.n754 out_p.t534 7.173
R30468 out_p.n754 out_p.t3175 7.173
R30469 out_p.n753 out_p.t1837 7.173
R30470 out_p.n753 out_p.t2761 7.173
R30471 out_p.n752 out_p.t3291 7.173
R30472 out_p.n752 out_p.t1279 7.173
R30473 out_p.n751 out_p.t3037 7.173
R30474 out_p.n751 out_p.t1659 7.173
R30475 out_p.n750 out_p.t2562 7.173
R30476 out_p.n750 out_p.t1550 7.173
R30477 out_p.n749 out_p.t1021 7.173
R30478 out_p.n749 out_p.t2106 7.173
R30479 out_p.n739 out_p.t2454 7.173
R30480 out_p.n739 out_p.t2308 7.173
R30481 out_p.n738 out_p.t846 7.173
R30482 out_p.n738 out_p.t1746 7.173
R30483 out_p.n737 out_p.t1076 7.173
R30484 out_p.n737 out_p.t2239 7.173
R30485 out_p.n736 out_p.t1229 7.173
R30486 out_p.n736 out_p.t1026 7.173
R30487 out_p.n735 out_p.t3051 7.173
R30488 out_p.n735 out_p.t540 7.173
R30489 out_p.n734 out_p.t2250 7.173
R30490 out_p.n734 out_p.t2983 7.173
R30491 out_p.n733 out_p.t1030 7.173
R30492 out_p.n733 out_p.t2123 7.173
R30493 out_p.n732 out_p.t567 7.173
R30494 out_p.n732 out_p.t3211 7.173
R30495 out_p.n731 out_p.t967 7.173
R30496 out_p.n731 out_p.t1424 7.173
R30497 out_p.n730 out_p.t2976 7.173
R30498 out_p.n730 out_p.t1407 7.173
R30499 out_p.n729 out_p.t2554 7.173
R30500 out_p.n729 out_p.t1642 7.173
R30501 out_p.n728 out_p.t1848 7.173
R30502 out_p.n728 out_p.t2765 7.173
R30503 out_p.n727 out_p.t592 7.173
R30504 out_p.n727 out_p.t3239 7.173
R30505 out_p.n726 out_p.t1430 7.173
R30506 out_p.n726 out_p.t794 7.173
R30507 out_p.n725 out_p.t2219 7.173
R30508 out_p.n725 out_p.t551 7.173
R30509 out_p.n724 out_p.t3110 7.173
R30510 out_p.n724 out_p.t1940 7.173
R30511 out_p.n723 out_p.t669 7.173
R30512 out_p.n723 out_p.t3315 7.173
R30513 out_p.n722 out_p.t2449 7.173
R30514 out_p.n722 out_p.t3065 7.173
R30515 out_p.n721 out_p.t1421 7.173
R30516 out_p.n721 out_p.t2539 7.173
R30517 out_p.n720 out_p.t2124 7.173
R30518 out_p.n720 out_p.t1006 7.173
R30519 out_p.n715 out_p.t2667 7.173
R30520 out_p.n715 out_p.t739 7.173
R30521 out_p.n714 out_p.t3074 7.173
R30522 out_p.n714 out_p.t1141 7.173
R30523 out_p.n713 out_p.t3329 7.173
R30524 out_p.n713 out_p.t2709 7.173
R30525 out_p.n712 out_p.t1974 7.173
R30526 out_p.n712 out_p.t1576 7.173
R30527 out_p.n711 out_p.t1805 7.173
R30528 out_p.n711 out_p.t3370 7.173
R30529 out_p.n710 out_p.t815 7.173
R30530 out_p.n710 out_p.t2160 7.173
R30531 out_p.n709 out_p.t3255 7.173
R30532 out_p.n709 out_p.t2658 7.173
R30533 out_p.n708 out_p.t1198 7.173
R30534 out_p.n708 out_p.t1621 7.173
R30535 out_p.n707 out_p.t3008 7.173
R30536 out_p.n707 out_p.t2919 7.173
R30537 out_p.n706 out_p.t1227 7.173
R30538 out_p.n706 out_p.t680 7.173
R30539 out_p.n705 out_p.t2299 7.173
R30540 out_p.n705 out_p.t1347 7.173
R30541 out_p.n704 out_p.t3083 7.173
R30542 out_p.n704 out_p.t430 7.173
R30543 out_p.n703 out_p.t1481 7.173
R30544 out_p.n703 out_p.t1666 7.173
R30545 out_p.n702 out_p.t1100 7.173
R30546 out_p.n702 out_p.t2775 7.173
R30547 out_p.n701 out_p.t868 7.173
R30548 out_p.n701 out_p.t2519 7.173
R30549 out_p.n700 out_p.t463 7.173
R30550 out_p.n700 out_p.t807 7.173
R30551 out_p.n699 out_p.t1964 7.173
R30552 out_p.n699 out_p.t1795 7.173
R30553 out_p.n698 out_p.t3383 7.173
R30554 out_p.n698 out_p.t2505 7.173
R30555 out_p.n697 out_p.t1282 7.173
R30556 out_p.n697 out_p.t1994 7.173
R30557 out_p.n696 out_p.t1891 7.173
R30558 out_p.n696 out_p.t1540 7.173
R30559 out_p.n691 out_p.t1567 7.173
R30560 out_p.n691 out_p.t917 7.173
R30561 out_p.n690 out_p.t2383 7.173
R30562 out_p.n690 out_p.t2650 7.173
R30563 out_p.n689 out_p.t2135 7.173
R30564 out_p.n689 out_p.t2883 7.173
R30565 out_p.n688 out_p.t2652 7.173
R30566 out_p.n688 out_p.t1898 7.173
R30567 out_p.n687 out_p.t857 7.173
R30568 out_p.n687 out_p.t1614 7.173
R30569 out_p.n686 out_p.t3310 7.173
R30570 out_p.n686 out_p.t1273 7.173
R30571 out_p.n685 out_p.t1917 7.173
R30572 out_p.n685 out_p.t2820 7.173
R30573 out_p.n684 out_p.t905 7.173
R30574 out_p.n684 out_p.t3325 7.173
R30575 out_p.n683 out_p.t1767 7.173
R30576 out_p.n683 out_p.t1202 7.173
R30577 out_p.n682 out_p.t3328 7.173
R30578 out_p.n682 out_p.t1832 7.173
R30579 out_p.n681 out_p.t2902 7.173
R30580 out_p.n681 out_p.t1855 7.173
R30581 out_p.n680 out_p.t464 7.173
R30582 out_p.n680 out_p.t2861 7.173
R30583 out_p.n679 out_p.t943 7.173
R30584 out_p.n679 out_p.t3345 7.173
R30585 out_p.n678 out_p.t2075 7.173
R30586 out_p.n678 out_p.t891 7.173
R30587 out_p.n677 out_p.t1598 7.173
R30588 out_p.n677 out_p.t663 7.173
R30589 out_p.n676 out_p.t1414 7.173
R30590 out_p.n676 out_p.t2225 7.173
R30591 out_p.n675 out_p.t1010 7.173
R30592 out_p.n675 out_p.t3404 7.173
R30593 out_p.n674 out_p.t761 7.173
R30594 out_p.n674 out_p.t3163 7.173
R30595 out_p.n673 out_p.t2862 7.173
R30596 out_p.n673 out_p.t2349 7.173
R30597 out_p.n672 out_p.t2628 7.173
R30598 out_p.n672 out_p.t1851 7.173
R30599 out_p.n667 out_p.t717 7.173
R30600 out_p.n667 out_p.t2203 7.173
R30601 out_p.n666 out_p.t1130 7.173
R30602 out_p.n666 out_p.t2380 7.173
R30603 out_p.n665 out_p.t2692 7.173
R30604 out_p.n665 out_p.t525 7.173
R30605 out_p.n664 out_p.t1542 7.173
R30606 out_p.n664 out_p.t2965 7.173
R30607 out_p.n663 out_p.t3354 7.173
R30608 out_p.n663 out_p.t1157 7.173
R30609 out_p.n662 out_p.t2068 7.173
R30610 out_p.n662 out_p.t1905 7.173
R30611 out_p.n661 out_p.t2635 7.173
R30612 out_p.n661 out_p.t2497 7.173
R30613 out_p.n660 out_p.t1654 7.173
R30614 out_p.n660 out_p.t2313 7.173
R30615 out_p.n659 out_p.t2814 7.173
R30616 out_p.n659 out_p.t745 7.173
R30617 out_p.n658 out_p.t698 7.173
R30618 out_p.n658 out_p.t1025 7.173
R30619 out_p.n657 out_p.t2429 7.173
R30620 out_p.n657 out_p.t600 7.173
R30621 out_p.n656 out_p.t1383 7.173
R30622 out_p.n656 out_p.t1450 7.173
R30623 out_p.n655 out_p.t1712 7.173
R30624 out_p.n655 out_p.t2364 7.173
R30625 out_p.n654 out_p.t2795 7.173
R30626 out_p.n654 out_p.t3118 7.173
R30627 out_p.n653 out_p.t2541 7.173
R30628 out_p.n653 out_p.t2864 7.173
R30629 out_p.n652 out_p.t831 7.173
R30630 out_p.n652 out_p.t1132 7.173
R30631 out_p.n651 out_p.t1840 7.173
R30632 out_p.n651 out_p.t1444 7.173
R30633 out_p.n650 out_p.t1413 7.173
R30634 out_p.n650 out_p.t1993 7.173
R30635 out_p.n649 out_p.t1959 7.173
R30636 out_p.n649 out_p.t3187 7.173
R30637 out_p.n648 out_p.t1518 7.173
R30638 out_p.n648 out_p.t2949 7.173
R30639 out_p.n643 out_p.t890 7.173
R30640 out_p.n643 out_p.t1047 7.173
R30641 out_p.n642 out_p.t2627 7.173
R30642 out_p.n642 out_p.t2774 7.173
R30643 out_p.n641 out_p.t2857 7.173
R30644 out_p.n641 out_p.t3010 7.173
R30645 out_p.n640 out_p.t1854 7.173
R30646 out_p.n640 out_p.t2179 7.173
R30647 out_p.n639 out_p.t2232 7.173
R30648 out_p.n639 out_p.t2151 7.173
R30649 out_p.n638 out_p.t1302 7.173
R30650 out_p.n638 out_p.t511 7.173
R30651 out_p.n637 out_p.t2802 7.173
R30652 out_p.n637 out_p.t2953 7.173
R30653 out_p.n636 out_p.t3342 7.173
R30654 out_p.n636 out_p.t2909 7.173
R30655 out_p.n635 out_p.t435 7.173
R30656 out_p.n635 out_p.t1425 7.173
R30657 out_p.n634 out_p.t1938 7.173
R30658 out_p.n634 out_p.t1874 7.173
R30659 out_p.n633 out_p.t1900 7.173
R30660 out_p.n633 out_p.t1717 7.173
R30661 out_p.n632 out_p.t2886 7.173
R30662 out_p.n632 out_p.t1134 7.173
R30663 out_p.n631 out_p.t3363 7.173
R30664 out_p.n631 out_p.t2942 7.173
R30665 out_p.n630 out_p.t919 7.173
R30666 out_p.n630 out_p.t499 7.173
R30667 out_p.n629 out_p.t684 7.173
R30668 out_p.n629 out_p.t2261 7.173
R30669 out_p.n628 out_p.t1250 7.173
R30670 out_p.n628 out_p.t2153 7.173
R30671 out_p.n627 out_p.t440 7.173
R30672 out_p.n627 out_p.t2996 7.173
R30673 out_p.n626 out_p.t3193 7.173
R30674 out_p.n626 out_p.t2759 7.173
R30675 out_p.n625 out_p.t2307 7.173
R30676 out_p.n625 out_p.t1596 7.173
R30677 out_p.n624 out_p.t1806 7.173
R30678 out_p.n624 out_p.t2142 7.173
R30679 out_p.n619 out_p.t1370 7.173
R30680 out_p.n619 out_p.t2518 7.173
R30681 out_p.n618 out_p.t2177 7.173
R30682 out_p.n618 out_p.t2947 7.173
R30683 out_p.n617 out_p.t1705 7.173
R30684 out_p.n617 out_p.t3186 7.173
R30685 out_p.n616 out_p.t2521 7.173
R30686 out_p.n616 out_p.t1446 7.173
R30687 out_p.n615 out_p.t736 7.173
R30688 out_p.n615 out_p.t1565 7.173
R30689 out_p.n614 out_p.t3191 7.173
R30690 out_p.n614 out_p.t677 7.173
R30691 out_p.n613 out_p.t1449 7.173
R30692 out_p.n613 out_p.t3124 7.173
R30693 out_p.n612 out_p.t1865 7.173
R30694 out_p.n612 out_p.t1039 7.173
R30695 out_p.n611 out_p.t2584 7.173
R30696 out_p.n611 out_p.t2013 7.173
R30697 out_p.n610 out_p.t805 7.173
R30698 out_p.n610 out_p.t455 7.173
R30699 out_p.n609 out_p.t1263 7.173
R30700 out_p.n609 out_p.t3024 7.173
R30701 out_p.n608 out_p.t1417 7.173
R30702 out_p.n608 out_p.t583 7.173
R30703 out_p.n607 out_p.t1922 7.173
R30704 out_p.n607 out_p.t1057 7.173
R30705 out_p.n606 out_p.t2896 7.173
R30706 out_p.n606 out_p.t2331 7.173
R30707 out_p.n605 out_p.t2664 7.173
R30708 out_p.n605 out_p.t1831 7.173
R30709 out_p.n604 out_p.t929 7.173
R30710 out_p.n604 out_p.t1583 7.173
R30711 out_p.n603 out_p.t2060 7.173
R30712 out_p.n603 out_p.t1117 7.173
R30713 out_p.n602 out_p.t1579 7.173
R30714 out_p.n602 out_p.t882 7.173
R30715 out_p.n601 out_p.t2749 7.173
R30716 out_p.n601 out_p.t2222 7.173
R30717 out_p.n600 out_p.t1175 7.173
R30718 out_p.n600 out_p.t2469 7.173
R30719 out_p.n595 out_p.t2675 7.173
R30720 out_p.n595 out_p.t2417 7.173
R30721 out_p.n594 out_p.t3088 7.173
R30722 out_p.n594 out_p.t2133 7.173
R30723 out_p.n593 out_p.t3338 7.173
R30724 out_p.n593 out_p.t1594 7.173
R30725 out_p.n592 out_p.t2019 7.173
R30726 out_p.n592 out_p.t1174 7.173
R30727 out_p.n591 out_p.t1838 7.173
R30728 out_p.n591 out_p.t715 7.173
R30729 out_p.n590 out_p.t827 7.173
R30730 out_p.n590 out_p.t3165 7.173
R30731 out_p.n589 out_p.t3270 7.173
R30732 out_p.n589 out_p.t2472 7.173
R30733 out_p.n588 out_p.t608 7.173
R30734 out_p.n588 out_p.t1911 7.173
R30735 out_p.n587 out_p.t2074 7.173
R30736 out_p.n587 out_p.t1156 7.173
R30737 out_p.n586 out_p.t3012 7.173
R30738 out_p.n586 out_p.t830 7.173
R30739 out_p.n585 out_p.t2600 7.173
R30740 out_p.n585 out_p.t2516 7.173
R30741 out_p.n584 out_p.t1996 7.173
R30742 out_p.n584 out_p.t1607 7.173
R30743 out_p.n583 out_p.t639 7.173
R30744 out_p.n583 out_p.t1960 7.173
R30745 out_p.n582 out_p.t1504 7.173
R30746 out_p.n582 out_p.t2925 7.173
R30747 out_p.n581 out_p.t1460 7.173
R30748 out_p.n581 out_p.t2680 7.173
R30749 out_p.n580 out_p.t3148 7.173
R30750 out_p.n580 out_p.t959 7.173
R30751 out_p.n579 out_p.t700 7.173
R30752 out_p.n579 out_p.t2129 7.173
R30753 out_p.n578 out_p.t459 7.173
R30754 out_p.n578 out_p.t1618 7.173
R30755 out_p.n577 out_p.t1262 7.173
R30756 out_p.n577 out_p.t2727 7.173
R30757 out_p.n576 out_p.t1951 7.173
R30758 out_p.n576 out_p.t1159 7.173
R30759 out_p.n571 out_p.t2838 7.173
R30760 out_p.n571 out_p.t3181 7.173
R30761 out_p.n570 out_p.t3265 7.173
R30762 out_p.n570 out_p.t1754 7.173
R30763 out_p.n569 out_p.t2008 7.173
R30764 out_p.n569 out_p.t1563 7.173
R30765 out_p.n568 out_p.t1280 7.173
R30766 out_p.n568 out_p.t675 7.173
R30767 out_p.n567 out_p.t2193 7.173
R30768 out_p.n567 out_p.t2115 7.173
R30769 out_p.n566 out_p.t999 7.173
R30770 out_p.n566 out_p.t2647 7.173
R30771 out_p.n565 out_p.t431 7.173
R30772 out_p.n565 out_p.t1455 7.173
R30773 out_p.n564 out_p.t1524 7.173
R30774 out_p.n564 out_p.t1062 7.173
R30775 out_p.n563 out_p.t1318 7.173
R30776 out_p.n563 out_p.t590 7.173
R30777 out_p.n562 out_p.t1129 7.173
R30778 out_p.n562 out_p.t1738 7.173
R30779 out_p.n561 out_p.t716 7.173
R30780 out_p.n561 out_p.t3060 7.173
R30781 out_p.n560 out_p.t1640 7.173
R30782 out_p.n560 out_p.t621 7.173
R30783 out_p.n559 out_p.t1636 7.173
R30784 out_p.n559 out_p.t1078 7.173
R30785 out_p.n558 out_p.t3238 7.173
R30786 out_p.n558 out_p.t2382 7.173
R30787 out_p.n557 out_p.t2993 7.173
R30788 out_p.n557 out_p.t1888 7.173
R30789 out_p.n556 out_p.t2576 7.173
R30790 out_p.n556 out_p.t1801 7.173
R30791 out_p.n555 out_p.t1939 7.173
R30792 out_p.n555 out_p.t1140 7.173
R30793 out_p.n554 out_p.t2265 7.173
R30794 out_p.n554 out_p.t912 7.173
R30795 out_p.n553 out_p.t554 7.173
R30796 out_p.n553 out_p.t886 7.173
R30797 out_p.n552 out_p.t1286 7.173
R30798 out_p.n552 out_p.t657 7.173
R30799 out_p.n547 out_p.t1011 7.173
R30800 out_p.n547 out_p.t1941 7.173
R30801 out_p.n546 out_p.t2725 7.173
R30802 out_p.n546 out_p.t553 7.173
R30803 out_p.n545 out_p.t2972 7.173
R30804 out_p.n545 out_p.t800 7.173
R30805 out_p.n544 out_p.t2083 7.173
R30806 out_p.n544 out_p.t3242 7.173
R30807 out_p.n543 out_p.t1966 7.173
R30808 out_p.n543 out_p.t2767 7.173
R30809 out_p.n542 out_p.t467 7.173
R30810 out_p.n542 out_p.t1651 7.173
R30811 out_p.n541 out_p.t2906 7.173
R30812 out_p.n541 out_p.t721 7.173
R30813 out_p.n540 out_p.t2694 7.173
R30814 out_p.n540 out_p.t3017 7.173
R30815 out_p.n539 out_p.t2169 7.173
R30816 out_p.n539 out_p.t3390 7.173
R30817 out_p.n538 out_p.t1494 7.173
R30818 out_p.n538 out_p.t2110 7.173
R30819 out_p.n537 out_p.t3379 7.173
R30820 out_p.n537 out_p.t2356 7.173
R30821 out_p.n536 out_p.t942 7.173
R30822 out_p.n536 out_p.t2561 7.173
R30823 out_p.n535 out_p.t2716 7.173
R30824 out_p.n535 out_p.t3043 7.173
R30825 out_p.n534 out_p.t2434 7.173
R30826 out_p.n534 out_p.t597 7.173
R30827 out_p.n533 out_p.t1511 7.173
R30828 out_p.n533 out_p.t1308 7.173
R30829 out_p.n532 out_p.t1709 7.173
R30830 out_p.n532 out_p.t2358 7.173
R30831 out_p.n531 out_p.t2790 7.173
R30832 out_p.n531 out_p.t3116 7.173
R30833 out_p.n530 out_p.t2536 7.173
R30834 out_p.n530 out_p.t2856 7.173
R30835 out_p.n529 out_p.t1509 7.173
R30836 out_p.n529 out_p.t1603 7.173
R30837 out_p.n528 out_p.t2029 7.173
R30838 out_p.n528 out_p.t3219 7.173
R30839 out_p.n523 out_p.t1215 7.173
R30840 out_p.n523 out_p.t2644 7.173
R30841 out_p.n522 out_p.t1686 7.173
R30842 out_p.n522 out_p.t3046 7.173
R30843 out_p.n521 out_p.t2192 7.173
R30844 out_p.n521 out_p.t3300 7.173
R30845 out_p.n520 out_p.t998 7.173
R30846 out_p.n520 out_p.t1868 7.173
R30847 out_p.n519 out_p.t521 7.173
R30848 out_p.n519 out_p.t1758 7.173
R30849 out_p.n518 out_p.t2963 7.173
R30850 out_p.n518 out_p.t779 7.173
R30851 out_p.n517 out_p.t2049 7.173
R30852 out_p.n517 out_p.t3223 7.173
R30853 out_p.n516 out_p.t1660 7.173
R30854 out_p.n516 out_p.t1359 7.173
R30855 out_p.n515 out_p.t2540 7.173
R30856 out_p.n515 out_p.t496 7.173
R30857 out_p.n514 out_p.t1150 7.173
R30858 out_p.n514 out_p.t2809 7.173
R30859 out_p.n513 out_p.t755 7.173
R30860 out_p.n513 out_p.t1071 7.173
R30861 out_p.n512 out_p.t1711 7.173
R30862 out_p.n512 out_p.t2363 7.173
R30863 out_p.n511 out_p.t1762 7.173
R30864 out_p.n511 out_p.t1313 7.173
R30865 out_p.n510 out_p.t3273 7.173
R30866 out_p.n510 out_p.t1695 7.173
R30867 out_p.n509 out_p.t3021 7.173
R30868 out_p.n509 out_p.t3349 7.173
R30869 out_p.n508 out_p.t2615 7.173
R30870 out_p.n508 out_p.t2938 7.173
R30871 out_p.n507 out_p.t2021 7.173
R30872 out_p.n507 out_p.t494 7.173
R30873 out_p.n506 out_p.t2319 7.173
R30874 out_p.n506 out_p.t2257 7.173
R30875 out_p.n505 out_p.t1190 7.173
R30876 out_p.n505 out_p.t2441 7.173
R30877 out_p.n504 out_p.t976 7.173
R30878 out_p.n504 out_p.t1766 7.173
R30879 out_p.n499 out_p.t1244 7.173
R30880 out_p.n499 out_p.t1532 7.173
R30881 out_p.n498 out_p.t803 7.173
R30882 out_p.n498 out_p.t2335 7.173
R30883 out_p.n497 out_p.t1044 7.173
R30884 out_p.n497 out_p.t2043 7.173
R30885 out_p.n496 out_p.t1212 7.173
R30886 out_p.n496 out_p.t2625 7.173
R30887 out_p.n495 out_p.t3007 7.173
R30888 out_p.n495 out_p.t839 7.173
R30889 out_p.n494 out_p.t2167 7.173
R30890 out_p.n494 out_p.t3283 7.173
R30891 out_p.n493 out_p.t983 7.173
R30892 out_p.n493 out_p.t1809 7.173
R30893 out_p.n492 out_p.t3066 7.173
R30894 out_p.n492 out_p.t3384 7.173
R30895 out_p.n491 out_p.t1756 7.173
R30896 out_p.n491 out_p.t3199 7.173
R30897 out_p.n490 out_p.t2201 7.173
R30898 out_p.n490 out_p.t2046 7.173
R30899 out_p.n489 out_p.t1410 7.173
R30900 out_p.n489 out_p.t1982 7.173
R30901 out_p.n488 out_p.t2619 7.173
R30902 out_p.n488 out_p.t2941 7.173
R30903 out_p.n487 out_p.t3090 7.173
R30904 out_p.n487 out_p.t3403 7.173
R30905 out_p.n486 out_p.t652 7.173
R30906 out_p.n486 out_p.t972 7.173
R30907 out_p.n485 out_p.t1338 7.173
R30908 out_p.n485 out_p.t714 7.173
R30909 out_p.n484 out_p.t2458 7.173
R30910 out_p.n484 out_p.t1298 7.173
R30911 out_p.n483 out_p.t3160 7.173
R30912 out_p.n483 out_p.t1774 7.173
R30913 out_p.n482 out_p.t2915 7.173
R30914 out_p.n482 out_p.t3235 7.173
R30915 out_p.n481 out_p.t2416 7.173
R30916 out_p.n481 out_p.t2836 7.173
R30917 out_p.n480 out_p.t1622 7.173
R30918 out_p.n480 out_p.t2598 7.173
R30919 out_p.n475 out_p.t2621 7.173
R30920 out_p.n475 out_p.t702 7.173
R30921 out_p.n474 out_p.t3023 7.173
R30922 out_p.n474 out_p.t1099 7.173
R30923 out_p.n473 out_p.t3277 7.173
R30924 out_p.n473 out_p.t2673 7.173
R30925 out_p.n472 out_p.t1765 7.173
R30926 out_p.n472 out_p.t1506 7.173
R30927 out_p.n471 out_p.t1721 7.173
R30928 out_p.n471 out_p.t3334 7.173
R30929 out_p.n470 out_p.t762 7.173
R30930 out_p.n470 out_p.t1999 7.173
R30931 out_p.n469 out_p.t3205 7.173
R30932 out_p.n469 out_p.t2604 7.173
R30933 out_p.n468 out_p.t2482 7.173
R30934 out_p.n468 out_p.t760 7.173
R30935 out_p.n467 out_p.t1246 7.173
R30936 out_p.n467 out_p.t2431 7.173
R30937 out_p.n466 out_p.t2827 7.173
R30938 out_p.n466 out_p.t3168 7.173
R30939 out_p.n465 out_p.t1085 7.173
R30940 out_p.n465 out_p.t2752 7.173
R30941 out_p.n464 out_p.t2394 7.173
R30942 out_p.n464 out_p.t1259 7.173
R30943 out_p.n463 out_p.t1341 7.173
R30944 out_p.n463 out_p.t782 7.173
R30945 out_p.n462 out_p.t1859 7.173
R30946 out_p.n462 out_p.t1769 7.173
R30947 out_p.n461 out_p.t3365 7.173
R30948 out_p.n461 out_p.t2419 7.173
R30949 out_p.n460 out_p.t2958 7.173
R30950 out_p.n460 out_p.t3304 7.173
R30951 out_p.n459 out_p.t516 7.173
R30952 out_p.n459 out_p.t855 7.173
R30953 out_p.n458 out_p.t1325 7.173
R30954 out_p.n458 out_p.t614 7.173
R30955 out_p.n457 out_p.t1240 7.173
R30956 out_p.n457 out_p.t1909 7.173
R30957 out_p.n456 out_p.t1684 7.173
R30958 out_p.n456 out_p.t1476 7.173
R30959 out_p.n451 out_p.t1503 7.173
R30960 out_p.n451 out_p.t867 7.173
R30961 out_p.n450 out_p.t2296 7.173
R30962 out_p.n450 out_p.t2594 7.173
R30963 out_p.n449 out_p.t1978 7.173
R30964 out_p.n449 out_p.t2834 7.173
R30965 out_p.n448 out_p.t2597 7.173
R30966 out_p.n448 out_p.t1797 7.173
R30967 out_p.n447 out_p.t818 7.173
R30968 out_p.n447 out_p.t1926 7.173
R30969 out_p.n446 out_p.t3263 7.173
R30970 out_p.n446 out_p.t2381 7.173
R30971 out_p.n445 out_p.t1726 7.173
R30972 out_p.n445 out_p.t2777 7.173
R30973 out_p.n444 out_p.t3400 7.173
R30974 out_p.n444 out_p.t2117 7.173
R30975 out_p.n443 out_p.t3093 7.173
R30976 out_p.n443 out_p.t909 7.173
R30977 out_p.n442 out_p.t2137 7.173
R30978 out_p.n442 out_p.t2607 7.173
R30979 out_p.n441 out_p.t2037 7.173
R30980 out_p.n441 out_p.t874 7.173
R30981 out_p.n440 out_p.t2959 7.173
R30982 out_p.n440 out_p.t1958 7.173
R30983 out_p.n439 out_p.t437 7.173
R30984 out_p.n439 out_p.t2196 7.173
R30985 out_p.n438 out_p.t995 7.173
R30986 out_p.n438 out_p.t3389 7.173
R30987 out_p.n437 out_p.t738 7.173
R30988 out_p.n437 out_p.t3156 7.173
R30989 out_p.n436 out_p.t2475 7.173
R30990 out_p.n436 out_p.t2732 7.173
R30991 out_p.n435 out_p.t1985 7.173
R30992 out_p.n435 out_p.t2444 7.173
R30993 out_p.n434 out_p.t3261 7.173
R30994 out_p.n434 out_p.t1545 7.173
R30995 out_p.n433 out_p.t2823 7.173
R30996 out_p.n433 out_p.t2254 7.173
R30997 out_p.n432 out_p.t2571 7.173
R30998 out_p.n432 out_p.t1759 7.173
R30999 out_p.n427 out_p.t1029 7.173
R31000 out_p.n427 out_p.t2122 7.173
R31001 out_p.n426 out_p.t2744 7.173
R31002 out_p.n426 out_p.t2209 7.173
R31003 out_p.n425 out_p.t2987 7.173
R31004 out_p.n425 out_p.t480 7.173
R31005 out_p.n424 out_p.t2131 7.173
R31006 out_p.n424 out_p.t2924 7.173
R31007 out_p.n423 out_p.t2055 7.173
R31008 out_p.n423 out_p.t1118 7.173
R31009 out_p.n422 out_p.t482 7.173
R31010 out_p.n422 out_p.t1605 7.173
R31011 out_p.n421 out_p.t2926 7.173
R31012 out_p.n421 out_p.t1253 7.173
R31013 out_p.n420 out_p.t1992 7.173
R31014 out_p.n420 out_p.t1090 7.173
R31015 out_p.n419 out_p.t946 7.173
R31016 out_p.n419 out_p.t1384 7.173
R31017 out_p.n418 out_p.t863 7.173
R31018 out_p.n418 out_p.t2147 7.173
R31019 out_p.n417 out_p.t2499 7.173
R31020 out_p.n417 out_p.t3097 7.173
R31021 out_p.n416 out_p.t1906 7.173
R31022 out_p.n416 out_p.t659 7.173
R31023 out_p.n415 out_p.t2052 7.173
R31024 out_p.n415 out_p.t1116 7.173
R31025 out_p.n414 out_p.t2964 7.173
R31026 out_p.n414 out_p.t2470 7.173
R31027 out_p.n413 out_p.t2712 7.173
R31028 out_p.n413 out_p.t1968 7.173
R31029 out_p.n412 out_p.t1002 7.173
R31030 out_p.n412 out_p.t2012 7.173
R31031 out_p.n411 out_p.t2202 7.173
R31032 out_p.n411 out_p.t1173 7.173
R31033 out_p.n410 out_p.t1700 7.173
R31034 out_p.n410 out_p.t962 7.173
R31035 out_p.n409 out_p.t1522 7.173
R31036 out_p.n409 out_p.t3145 7.173
R31037 out_p.n408 out_p.t2064 7.173
R31038 out_p.n408 out_p.t2895 7.173
R31039 out_p.n403 out_p.t1169 7.173
R31040 out_p.n403 out_p.t1008 7.173
R31041 out_p.n402 out_p.t2922 7.173
R31042 out_p.n402 out_p.t2719 7.173
R31043 out_p.n401 out_p.t3161 7.173
R31044 out_p.n401 out_p.t2968 7.173
R31045 out_p.n400 out_p.t2462 7.173
R31046 out_p.n400 out_p.t2072 7.173
R31047 out_p.n399 out_p.t1530 7.173
R31048 out_p.n399 out_p.t1963 7.173
R31049 out_p.n398 out_p.t653 7.173
R31050 out_p.n398 out_p.t462 7.173
R31051 out_p.n397 out_p.t3091 7.173
R31052 out_p.n397 out_p.t2901 7.173
R31053 out_p.n396 out_p.t1217 7.173
R31054 out_p.n396 out_p.t2050 7.173
R31055 out_p.n395 out_p.t2863 7.173
R31056 out_p.n395 out_p.t840 7.173
R31057 out_p.n394 out_p.t2485 7.173
R31058 out_p.n394 out_p.t883 7.173
R31059 out_p.n393 out_p.t2252 7.173
R31060 out_p.n393 out_p.t481 7.173
R31061 out_p.n392 out_p.t3059 7.173
R31062 out_p.n392 out_p.t2035 7.173
R31063 out_p.n391 out_p.t1201 7.173
R31064 out_p.n391 out_p.t2121 7.173
R31065 out_p.n390 out_p.t1077 7.173
R31066 out_p.n390 out_p.t2982 7.173
R31067 out_p.n389 out_p.t850 7.173
R31068 out_p.n389 out_p.t2741 7.173
R31069 out_p.n388 out_p.t1264 7.173
R31070 out_p.n388 out_p.t1024 7.173
R31071 out_p.n387 out_p.t1800 7.173
R31072 out_p.n387 out_p.t2238 7.173
R31073 out_p.n386 out_p.t3359 7.173
R31074 out_p.n386 out_p.t1745 7.173
R31075 out_p.n385 out_p.t2171 7.173
R31076 out_p.n385 out_p.t1468 7.173
R31077 out_p.n384 out_p.t2398 7.173
R31078 out_p.n384 out_p.t2017 7.173
R31079 out_p.n379 out_p.t2236 7.173
R31080 out_p.n379 out_p.t1149 7.173
R31081 out_p.n378 out_p.t2062 7.173
R31082 out_p.n378 out_p.t2893 7.173
R31083 out_p.n377 out_p.t1514 7.173
R31084 out_p.n377 out_p.t3144 7.173
R31085 out_p.n376 out_p.t1155 7.173
R31086 out_p.n376 out_p.t2397 7.173
R31087 out_p.n375 out_p.t699 7.173
R31088 out_p.n375 out_p.t1496 7.173
R31089 out_p.n374 out_p.t3147 7.173
R31090 out_p.n374 out_p.t635 7.173
R31091 out_p.n373 out_p.t2413 7.173
R31092 out_p.n373 out_p.t3070 7.173
R31093 out_p.n372 out_p.t881 7.173
R31094 out_p.n372 out_p.t2463 7.173
R31095 out_p.n371 out_p.t2393 7.173
R31096 out_p.n371 out_p.t2769 7.173
R31097 out_p.n370 out_p.t3302 7.173
R31098 out_p.n370 out_p.t1236 7.173
R31099 out_p.n369 out_p.t2876 7.173
R31100 out_p.n369 out_p.t2290 7.173
R31101 out_p.n368 out_p.t1348 7.173
R31102 out_p.n368 out_p.t3078 7.173
R31103 out_p.n367 out_p.t908 7.173
R31104 out_p.n367 out_p.t1459 7.173
R31105 out_p.n366 out_p.t2016 7.173
R31106 out_p.n366 out_p.t1098 7.173
R31107 out_p.n365 out_p.t1562 7.173
R31108 out_p.n365 out_p.t866 7.173
R31109 out_p.n364 out_p.t3422 7.173
R31110 out_p.n364 out_p.t458 7.173
R31111 out_p.n363 out_p.t988 7.173
R31112 out_p.n363 out_p.t1928 7.173
R31113 out_p.n362 out_p.t729 7.173
R31114 out_p.n362 out_p.t3381 7.173
R31115 out_p.n361 out_p.t2701 7.173
R31116 out_p.n361 out_p.t2090 7.173
R31117 out_p.n360 out_p.t1136 7.173
R31118 out_p.n360 out_p.t2367 7.173
R31119 out_p.n355 out_p.t2634 7.173
R31120 out_p.n355 out_p.t1862 7.173
R31121 out_p.n354 out_p.t3042 7.173
R31122 out_p.n354 out_p.t1836 7.173
R31123 out_p.n353 out_p.t3294 7.173
R31124 out_p.n353 out_p.t1310 7.173
R31125 out_p.n352 out_p.t1847 7.173
R31126 out_p.n352 out_p.t2807 7.173
R31127 out_p.n351 out_p.t1748 7.173
R31128 out_p.n351 out_p.t1023 7.173
R31129 out_p.n350 out_p.t771 7.173
R31130 out_p.n350 out_p.t1204 7.173
R31131 out_p.n349 out_p.t3217 7.173
R31132 out_p.n349 out_p.t2440 7.173
R31133 out_p.n348 out_p.t3104 7.173
R31134 out_p.n348 out_p.t2264 7.173
R31135 out_p.n347 out_p.t2793 7.173
R31136 out_p.n347 out_p.t617 7.173
R31137 out_p.n346 out_p.t2266 7.173
R31138 out_p.n346 out_p.t1000 7.173
R31139 out_p.n345 out_p.t1477 7.173
R31140 out_p.n345 out_p.t575 7.173
R31141 out_p.n344 out_p.t2659 7.173
R31142 out_p.n344 out_p.t1409 7.173
R31143 out_p.n343 out_p.t3135 7.173
R31144 out_p.n343 out_p.t2306 7.173
R31145 out_p.n342 out_p.t687 7.173
R31146 out_p.n342 out_p.t3087 7.173
R31147 out_p.n341 out_p.t1351 7.173
R31148 out_p.n341 out_p.t2840 7.173
R31149 out_p.n340 out_p.t1470 7.173
R31150 out_p.n340 out_p.t1105 7.173
R31151 out_p.n339 out_p.t3197 7.173
R31152 out_p.n339 out_p.t2457 7.173
R31153 out_p.n338 out_p.t2956 7.173
R31154 out_p.n338 out_p.t1944 7.173
R31155 out_p.n337 out_p.t1337 7.173
R31156 out_p.n337 out_p.t3020 7.173
R31157 out_p.n336 out_p.t1741 7.173
R31158 out_p.n336 out_p.t2781 7.173
R31159 out_p.n331 out_p.t2801 7.173
R31160 out_p.n331 out_p.t879 7.173
R31161 out_p.n330 out_p.t3210 7.173
R31162 out_p.n330 out_p.t2614 7.173
R31163 out_p.n329 out_p.t1191 7.173
R31164 out_p.n329 out_p.t2845 7.173
R31165 out_p.n328 out_p.t2430 7.173
R31166 out_p.n328 out_p.t1829 7.173
R31167 out_p.n327 out_p.t2105 7.173
R31168 out_p.n327 out_p.t2100 7.173
R31169 out_p.n326 out_p.t952 7.173
R31170 out_p.n326 out_p.t1260 7.173
R31171 out_p.n325 out_p.t3387 7.173
R31172 out_p.n325 out_p.t2786 7.173
R31173 out_p.n324 out_p.t2527 7.173
R31174 out_p.n324 out_p.t2882 7.173
R31175 out_p.n323 out_p.t3410 7.173
R31176 out_p.n323 out_p.t3330 7.173
R31177 out_p.n322 out_p.t2011 7.173
R31178 out_p.n322 out_p.t1808 7.173
R31179 out_p.n321 out_p.t3220 7.173
R31180 out_p.n321 out_p.t1535 7.173
R31181 out_p.n320 out_p.t776 7.173
R31182 out_p.n320 out_p.t1109 7.173
R31183 out_p.n319 out_p.t2558 7.173
R31184 out_p.n319 out_p.t2910 7.173
R31185 out_p.n318 out_p.t1849 7.173
R31186 out_p.n318 out_p.t469 7.173
R31187 out_p.n317 out_p.t2230 7.173
R31188 out_p.n317 out_p.t2195 7.173
R31189 out_p.n316 out_p.t1441 7.173
R31190 out_p.n316 out_p.t2086 7.173
R31191 out_p.n315 out_p.t2640 7.173
R31192 out_p.n315 out_p.t2975 7.173
R31193 out_p.n314 out_p.t1070 7.173
R31194 out_p.n314 out_p.t2731 7.173
R31195 out_p.n313 out_p.t517 7.173
R31196 out_p.n313 out_p.t2286 7.173
R31197 out_p.n312 out_p.t1270 7.173
R31198 out_p.n312 out_p.t1783 7.173
R31199 out_p.n307 out_p.t1815 7.173
R31200 out_p.n307 out_p.t3123 7.173
R31201 out_p.n306 out_p.t1740 7.173
R31202 out_p.n306 out_p.t2415 7.173
R31203 out_p.n305 out_p.t1272 7.173
R31204 out_p.n305 out_p.t1462 7.173
R31205 out_p.n304 out_p.t2783 7.173
R31206 out_p.n304 out_p.t607 7.173
R31207 out_p.n303 out_p.t1005 7.173
R31208 out_p.n303 out_p.t1896 7.173
R31209 out_p.n302 out_p.t444 7.173
R31210 out_p.n302 out_p.t2569 7.173
R31211 out_p.n301 out_p.t1225 7.173
R31212 out_p.n301 out_p.t2392 7.173
R31213 out_p.n300 out_p.t2301 7.173
R31214 out_p.n300 out_p.t2221 7.173
R31215 out_p.n299 out_p.t515 7.173
R31216 out_p.n299 out_p.t1971 7.173
R31217 out_p.n298 out_p.t1020 7.173
R31218 out_p.n298 out_p.t2653 7.173
R31219 out_p.n297 out_p.t598 7.173
R31220 out_p.n297 out_p.t918 7.173
R31221 out_p.n296 out_p.t1443 7.173
R31222 out_p.n296 out_p.t2036 7.173
R31223 out_p.n295 out_p.t2359 7.173
R31224 out_p.n295 out_p.t1309 7.173
R31225 out_p.n294 out_p.t3115 7.173
R31226 out_p.n294 out_p.t438 7.173
R31227 out_p.n293 out_p.t2860 7.173
R31228 out_p.n293 out_p.t3190 7.173
R31229 out_p.n292 out_p.t1128 7.173
R31230 out_p.n292 out_p.t2776 7.173
R31231 out_p.n291 out_p.t1405 7.173
R31232 out_p.n291 out_p.t2455 7.173
R31233 out_p.n290 out_p.t1984 7.173
R31234 out_p.n290 out_p.t1704 7.173
R31235 out_p.n289 out_p.t3002 7.173
R31236 out_p.n289 out_p.t835 7.173
R31237 out_p.n288 out_p.t2763 7.173
R31238 out_p.n288 out_p.t582 7.173
R31239 out_p.n283 out_p.t1192 7.173
R31240 out_p.n283 out_p.t2583 7.173
R31241 out_p.n282 out_p.t1610 7.173
R31242 out_p.n282 out_p.t3000 7.173
R31243 out_p.n281 out_p.t2099 7.173
R31244 out_p.n281 out_p.t3248 7.173
R31245 out_p.n280 out_p.t951 7.173
R31246 out_p.n280 out_p.t1681 7.173
R31247 out_p.n279 out_p.t474 7.173
R31248 out_p.n279 out_p.t1665 7.173
R31249 out_p.n278 out_p.t2914 7.173
R31250 out_p.n278 out_p.t728 7.173
R31251 out_p.n277 out_p.t1943 7.173
R31252 out_p.n277 out_p.t3179 7.173
R31253 out_p.n276 out_p.t2563 7.173
R31254 out_p.n276 out_p.t2885 7.173
R31255 out_p.n275 out_p.t2330 7.173
R31256 out_p.n275 out_p.t1798 7.173
R31257 out_p.n274 out_p.t2128 7.173
R31258 out_p.n274 out_p.t1828 7.173
R31259 out_p.n273 out_p.t3254 7.173
R31260 out_p.n273 out_p.t1561 7.173
R31261 out_p.n272 out_p.t814 7.173
R31262 out_p.n272 out_p.t1112 7.173
R31263 out_p.n271 out_p.t2590 7.173
R31264 out_p.n271 out_p.t2918 7.173
R31265 out_p.n270 out_p.t1973 7.173
R31266 out_p.n270 out_p.t479 7.173
R31267 out_p.n269 out_p.t2288 7.173
R31268 out_p.n269 out_p.t2207 7.173
R31269 out_p.n268 out_p.t1493 7.173
R31270 out_p.n268 out_p.t2109 7.173
R31271 out_p.n267 out_p.t2668 7.173
R31272 out_p.n267 out_p.t2981 7.173
R31273 out_p.n266 out_p.t1097 7.173
R31274 out_p.n266 out_p.t2738 7.173
R31275 out_p.n265 out_p.t1146 7.173
R31276 out_p.n265 out_p.t2442 7.173
R31277 out_p.n264 out_p.t925 7.173
R31278 out_p.n264 out_p.t1570 7.173
R31279 out_p.n259 out_p.t1780 7.173
R31280 out_p.n259 out_p.t1454 7.173
R31281 out_p.n258 out_p.t1662 7.173
R31282 out_p.n258 out_p.t2249 7.173
R31283 out_p.n257 out_p.t1275 7.173
R31284 out_p.n257 out_p.t1895 7.173
R31285 out_p.n256 out_p.t2762 7.173
R31286 out_p.n256 out_p.t2565 7.173
R31287 out_p.n255 out_p.t986 7.173
R31288 out_p.n255 out_p.t788 7.173
R31289 out_p.n254 out_p.t3420 7.173
R31290 out_p.n254 out_p.t3231 7.173
R31291 out_p.n253 out_p.t2283 7.173
R31292 out_p.n253 out_p.t1592 7.173
R31293 out_p.n252 out_p.t1817 7.173
R31294 out_p.n252 out_p.t1329 7.173
R31295 out_p.n251 out_p.t2613 7.173
R31296 out_p.n251 out_p.t571 7.173
R31297 out_p.n250 out_p.t778 7.173
R31298 out_p.n250 out_p.t2678 7.173
R31299 out_p.n249 out_p.t1237 7.173
R31300 out_p.n249 out_p.t958 7.173
R31301 out_p.n248 out_p.t1200 7.173
R31302 out_p.n248 out_p.t2120 7.173
R31303 out_p.n247 out_p.t1879 7.173
R31304 out_p.n247 out_p.t2443 7.173
R31305 out_p.n246 out_p.t2873 7.173
R31306 out_p.n246 out_p.t1534 7.173
R31307 out_p.n245 out_p.t2643 7.173
R31308 out_p.n245 out_p.t3215 7.173
R31309 out_p.n244 out_p.t903 7.173
R31310 out_p.n244 out_p.t2808 7.173
R31311 out_p.n243 out_p.t2006 7.173
R31312 out_p.n243 out_p.t1315 7.173
R31313 out_p.n242 out_p.t1555 7.173
R31314 out_p.n242 out_p.t1835 7.173
R31315 out_p.n241 out_p.t2984 7.173
R31316 out_p.n241 out_p.t2799 7.173
R31317 out_p.n240 out_p.t2740 7.173
R31318 out_p.n240 out_p.t2543 7.173
R31319 out_p.n235 out_p.t2905 7.173
R31320 out_p.n235 out_p.t1747 7.173
R31321 out_p.n234 out_p.t3331 7.173
R31322 out_p.n234 out_p.t1569 7.173
R31323 out_p.n233 out_p.t1501 7.173
R31324 out_p.n233 out_p.t2432 7.173
R31325 out_p.n232 out_p.t1353 7.173
R31326 out_p.n232 out_p.t2743 7.173
R31327 out_p.n231 out_p.t2315 7.173
R31328 out_p.n231 out_p.t963 7.173
R31329 out_p.n230 out_p.t1050 7.173
R31330 out_p.n230 out_p.t3395 7.173
R31331 out_p.n229 out_p.t1962 7.173
R31332 out_p.n229 out_p.t2210 7.173
R31333 out_p.n228 out_p.t585 7.173
R31334 out_p.n228 out_p.t1867 7.173
R31335 out_p.n227 out_p.t2141 7.173
R31336 out_p.n227 out_p.t1172 7.173
R31337 out_p.n226 out_p.t2992 7.173
R31338 out_p.n226 out_p.t811 7.173
R31339 out_p.n225 out_p.t2573 7.173
R31340 out_p.n225 out_p.t1241 7.173
R31341 out_p.n224 out_p.t1937 7.173
R31342 out_p.n224 out_p.t1458 7.173
R31343 out_p.n223 out_p.t616 7.173
R31344 out_p.n223 out_p.t1924 7.173
R31345 out_p.n222 out_p.t1474 7.173
R31346 out_p.n222 out_p.t2897 7.173
R31347 out_p.n221 out_p.t1207 7.173
R31348 out_p.n221 out_p.t2665 7.173
R31349 out_p.n220 out_p.t3131 7.173
R31350 out_p.n220 out_p.t935 7.173
R31351 out_p.n219 out_p.t685 7.173
R31352 out_p.n219 out_p.t2061 7.173
R31353 out_p.n218 out_p.t1267 7.173
R31354 out_p.n218 out_p.t1589 7.173
R31355 out_p.n217 out_p.t623 7.173
R31356 out_p.n217 out_p.t2967 7.173
R31357 out_p.n216 out_p.t1328 7.173
R31358 out_p.n216 out_p.t2717 7.173
R31359 out_p.n211 out_p.t2048 7.173
R31360 out_p.n211 out_p.t833 7.173
R31361 out_p.n210 out_p.t2159 7.173
R31362 out_p.n210 out_p.t2544 7.173
R31363 out_p.n209 out_p.t1343 7.173
R31364 out_p.n209 out_p.t2796 7.173
R31365 out_p.n208 out_p.t2889 7.173
R31366 out_p.n208 out_p.t1713 7.173
R31367 out_p.n207 out_p.t1089 7.173
R31368 out_p.n207 out_p.t1401 7.173
R31369 out_p.n206 out_p.t2343 7.173
R31370 out_p.n206 out_p.t2407 7.173
R31371 out_p.n205 out_p.t1333 7.173
R31372 out_p.n205 out_p.t2720 7.173
R31373 out_p.n204 out_p.t1623 7.173
R31374 out_p.n204 out_p.t2693 7.173
R31375 out_p.n203 out_p.t2522 7.173
R31376 out_p.n203 out_p.t1655 7.173
R31377 out_p.n202 out_p.t1281 7.173
R31378 out_p.n202 out_p.t1488 7.173
R31379 out_p.n201 out_p.t2379 7.173
R31380 out_p.n201 out_p.t3375 7.173
R31381 out_p.n200 out_p.t3134 7.173
R31382 out_p.n200 out_p.t939 7.173
R31383 out_p.n199 out_p.t1799 7.173
R31384 out_p.n199 out_p.t2713 7.173
R31385 out_p.n198 out_p.t1139 7.173
R31386 out_p.n198 out_p.t2401 7.173
R31387 out_p.n197 out_p.t911 7.173
R31388 out_p.n197 out_p.t1510 7.173
R31389 out_p.n196 out_p.t506 7.173
R31390 out_p.n196 out_p.t1701 7.173
R31391 out_p.n195 out_p.t2149 7.173
R31392 out_p.n195 out_p.t2789 7.173
R31393 out_p.n194 out_p.t434 7.173
R31394 out_p.n194 out_p.t2533 7.173
R31395 out_p.n193 out_p.t3119 7.173
R31396 out_p.n193 out_p.t2180 7.173
R31397 out_p.n192 out_p.t2865 7.173
R31398 out_p.n192 out_p.t1675 7.173
R31399 out_p.n187 out_p.t2386 7.173
R31400 out_p.n187 out_p.t1995 7.173
R31401 out_p.n186 out_p.t1274 7.173
R31402 out_p.n186 out_p.t2069 7.173
R31403 out_p.n185 out_p.t624 7.173
R31404 out_p.n185 out_p.t2452 7.173
R31405 out_p.n184 out_p.t3062 7.173
R31406 out_p.n184 out_p.t2868 7.173
R31407 out_p.n183 out_p.t2579 7.173
R31408 out_p.n183 out_p.t1075 7.173
R31409 out_p.n182 out_p.t1434 7.173
R31410 out_p.n182 out_p.t2342 7.173
R31411 out_p.n181 out_p.t548 7.173
R31412 out_p.n181 out_p.t1320 7.173
R31413 out_p.n180 out_p.t3013 7.173
R31414 out_p.n180 out_p.t1775 7.173
R31415 out_p.n179 out_p.t3157 7.173
R31416 out_p.n179 out_p.t1102 7.173
R31417 out_p.n178 out_p.t2107 7.173
R31418 out_p.n178 out_p.t1352 7.173
R31419 out_p.n177 out_p.t2328 7.173
R31420 out_p.n177 out_p.t2420 7.173
R31421 out_p.n176 out_p.t2557 7.173
R31422 out_p.n176 out_p.t3153 7.173
R31423 out_p.n175 out_p.t3036 7.173
R31424 out_p.n175 out_p.t1929 7.173
R31425 out_p.n174 out_p.t594 7.173
R31426 out_p.n174 out_p.t1161 7.173
R31427 out_p.n173 out_p.t1299 7.173
R31428 out_p.n173 out_p.t944 7.173
R31429 out_p.n172 out_p.t2350 7.173
R31430 out_p.n172 out_p.t529 7.173
R31431 out_p.n171 out_p.t3111 7.173
R31432 out_p.n171 out_p.t2293 7.173
R31433 out_p.n170 out_p.t2855 7.173
R31434 out_p.n170 out_p.t1432 7.173
R31435 out_p.n169 out_p.t3292 7.173
R31436 out_p.n169 out_p.t3095 7.173
R31437 out_p.n168 out_p.t3038 7.173
R31438 out_p.n168 out_p.t2843 7.173
R31439 out_p.n163 out_p.t1131 7.173
R31440 out_p.n163 out_p.t2402 7.173
R31441 out_p.n162 out_p.t2866 7.173
R31442 out_p.n162 out_p.t694 7.173
R31443 out_p.n161 out_p.t3120 7.173
R31444 out_p.n161 out_p.t945 7.173
R31445 out_p.n160 out_p.t2365 7.173
R31446 out_p.n160 out_p.t3378 7.173
R31447 out_p.n159 out_p.t1451 7.173
R31448 out_p.n159 out_p.t2903 7.173
R31449 out_p.n158 out_p.t601 7.173
R31450 out_p.n158 out_p.t1931 7.173
R31451 out_p.n157 out_p.t3044 7.173
R31452 out_p.n157 out_p.t864 7.173
R31453 out_p.n156 out_p.t2486 7.173
R31454 out_p.n156 out_p.t707 7.173
R31455 out_p.n155 out_p.t2262 7.173
R31456 out_p.n155 out_p.t1505 7.173
R31457 out_p.n154 out_p.t2804 7.173
R31458 out_p.n154 out_p.t3129 7.173
R31459 out_p.n153 out_p.t1069 7.173
R31460 out_p.n153 out_p.t2700 7.173
R31461 out_p.n152 out_p.t2360 7.173
R31462 out_p.n152 out_p.t1300 7.173
R31463 out_p.n151 out_p.t1304 7.173
R31464 out_p.n151 out_p.t731 7.173
R31465 out_p.n150 out_p.t1673 7.173
R31466 out_p.n150 out_p.t1668 7.173
R31467 out_p.n149 out_p.t3347 7.173
R31468 out_p.n149 out_p.t2126 7.173
R31469 out_p.n148 out_p.t2935 7.173
R31470 out_p.n148 out_p.t3250 7.173
R31471 out_p.n147 out_p.t493 7.173
R31472 out_p.n147 out_p.t812 7.173
R31473 out_p.n146 out_p.t2243 7.173
R31474 out_p.n146 out_p.t561 7.173
R31475 out_p.n145 out_p.t2022 7.173
R31476 out_p.n145 out_p.t1802 7.173
R31477 out_p.n144 out_p.t2320 7.173
R31478 out_p.n144 out_p.t3356 7.173
R31479 out_p.n139 out_p.t2032 7.173
R31480 out_p.n139 out_p.t2778 7.173
R31481 out_p.n138 out_p.t1967 7.173
R31482 out_p.n138 out_p.t3192 7.173
R31483 out_p.n137 out_p.t2471 7.173
R31484 out_p.n137 out_p.t429 7.173
R31485 out_p.n136 out_p.t1113 7.173
R31486 out_p.n136 out_p.t1301 7.173
R31487 out_p.n135 out_p.t660 7.173
R31488 out_p.n135 out_p.t2038 7.173
R31489 out_p.n134 out_p.t3098 7.173
R31490 out_p.n134 out_p.t920 7.173
R31491 out_p.n133 out_p.t2332 7.173
R31492 out_p.n133 out_p.t3364 7.173
R31493 out_p.n132 out_p.t3382 7.173
R31494 out_p.n132 out_p.t2371 7.173
R31495 out_p.n131 out_p.t2960 7.173
R31496 out_p.n131 out_p.t888 7.173
R31497 out_p.n130 out_p.t2044 7.173
R31498 out_p.n130 out_p.t504 7.173
R31499 out_p.n129 out_p.t1981 7.173
R31500 out_p.n129 out_p.t1685 7.173
R31501 out_p.n128 out_p.t2940 7.173
R31502 out_p.n128 out_p.t3256 7.173
R31503 out_p.n127 out_p.t3401 7.173
R31504 out_p.n127 out_p.t2506 7.173
R31505 out_p.n126 out_p.t970 7.173
R31506 out_p.n126 out_p.t2591 7.173
R31507 out_p.n125 out_p.t713 7.173
R31508 out_p.n125 out_p.t1043 7.173
R31509 out_p.n124 out_p.t2427 7.173
R31510 out_p.n124 out_p.t631 7.173
R31511 out_p.n123 out_p.t1656 7.173
R31512 out_p.n123 out_p.t1490 7.173
R31513 out_p.n122 out_p.t3232 7.173
R31514 out_p.n122 out_p.t1392 7.173
R31515 out_p.n121 out_p.t2669 7.173
R31516 out_p.n121 out_p.t491 7.173
R31517 out_p.n120 out_p.t1095 7.173
R31518 out_p.n120 out_p.t2244 7.173
R31519 out_p.n115 out_p.t452 7.173
R31520 out_p.n115 out_p.t1770 7.173
R31521 out_p.n114 out_p.t678 7.173
R31522 out_p.n114 out_p.t1637 7.173
R31523 out_p.n113 out_p.t913 7.173
R31524 out_p.n113 out_p.t1311 7.173
R31525 out_p.n112 out_p.t3360 7.173
R31526 out_p.n112 out_p.t2755 7.173
R31527 out_p.n111 out_p.t2880 7.173
R31528 out_p.n111 out_p.t978 7.173
R31529 out_p.n110 out_p.t1889 7.173
R31530 out_p.n110 out_p.t3411 7.173
R31531 out_p.n109 out_p.t851 7.173
R31532 out_p.n109 out_p.t2258 7.173
R31533 out_p.n108 out_p.t724 7.173
R31534 out_p.n108 out_p.t1072 7.173
R31535 out_p.n107 out_p.t2312 7.173
R31536 out_p.n107 out_p.t1822 7.173
R31537 out_p.n106 out_p.t3149 7.173
R31538 out_p.n106 out_p.t1857 7.173
R31539 out_p.n105 out_p.t2721 7.173
R31540 out_p.n105 out_p.t3071 7.173
R31541 out_p.n104 out_p.t2405 7.173
R31542 out_p.n104 out_p.t637 7.173
R31543 out_p.n103 out_p.t757 7.173
R31544 out_p.n103 out_p.t1091 7.173
R31545 out_p.n102 out_p.t1714 7.173
R31546 out_p.n102 out_p.t2411 7.173
R31547 out_p.n101 out_p.t2272 7.173
R31548 out_p.n101 out_p.t1923 7.173
R31549 out_p.n100 out_p.t3276 7.173
R31550 out_p.n100 out_p.t1861 7.173
R31551 out_p.n99 out_p.t834 7.173
R31552 out_p.n99 out_p.t1151 7.173
R31553 out_p.n98 out_p.t580 7.173
R31554 out_p.n98 out_p.t934 7.173
R31555 out_p.n97 out_p.t1648 7.173
R31556 out_p.n97 out_p.t2978 7.173
R31557 out_p.n96 out_p.t3343 7.173
R31558 out_p.n96 out_p.t2733 7.173
R31559 out_p.n91 out_p.t2750 7.173
R31560 out_p.n91 out_p.t2143 7.173
R31561 out_p.n90 out_p.t3166 7.173
R31562 out_p.n90 out_p.t2245 7.173
R31563 out_p.n89 out_p.t3406 7.173
R31564 out_p.n89 out_p.t492 7.173
R31565 out_p.n88 out_p.t2247 7.173
R31566 out_p.n88 out_p.t2934 7.173
R31567 out_p.n87 out_p.t1990 7.173
R31568 out_p.n87 out_p.t1126 7.173
R31569 out_p.n86 out_p.t893 7.173
R31570 out_p.n86 out_p.t1671 7.173
R31571 out_p.n85 out_p.t3348 7.173
R31572 out_p.n85 out_p.t2483 7.173
R31573 out_p.n84 out_p.t2510 7.173
R31574 out_p.n84 out_p.t526 7.173
R31575 out_p.n83 out_p.t791 7.173
R31576 out_p.n83 out_p.t2316 7.173
R31577 out_p.n82 out_p.t528 7.173
R31578 out_p.n82 out_p.t2932 7.173
R31579 out_p.n81 out_p.t1787 7.173
R31580 out_p.n81 out_p.t1178 7.173
R31581 out_p.n80 out_p.t3279 7.173
R31582 out_p.n80 out_p.t1633 7.173
R31583 out_p.n79 out_p.t1419 7.173
R31584 out_p.n79 out_p.t543 7.173
R31585 out_p.n78 out_p.t2623 7.173
R31586 out_p.n78 out_p.t2464 7.173
R31587 out_p.n77 out_p.t1058 7.173
R31588 out_p.n77 out_p.t1208 7.173
R31589 out_p.n76 out_p.t654 7.173
R31590 out_p.n76 out_p.t3052 7.173
R31591 out_p.n75 out_p.t1531 7.173
R31592 out_p.n75 out_p.t615 7.173
R31593 out_p.n74 out_p.t1584 7.173
R31594 out_p.n74 out_p.t2515 7.173
R31595 out_p.n73 out_p.t468 7.173
R31596 out_p.n73 out_p.t3154 7.173
R31597 out_p.n72 out_p.t2194 7.173
R31598 out_p.n72 out_p.t2907 7.173
R31599 out_p.n67 out_p.t2414 7.173
R31600 out_p.n67 out_p.t3069 7.173
R31601 out_p.n66 out_p.t1242 7.173
R31602 out_p.n66 out_p.t1844 7.173
R31603 out_p.n65 out_p.t640 7.173
R31604 out_p.n65 out_p.t1367 7.173
R31605 out_p.n64 out_p.t3075 7.173
R31606 out_p.n64 out_p.t560 7.173
R31607 out_p.n63 out_p.t2599 7.173
R31608 out_p.n63 out_p.t1703 7.173
R31609 out_p.n62 out_p.t1379 7.173
R31610 out_p.n62 out_p.t2520 7.173
R31611 out_p.n61 out_p.t563 7.173
R31612 out_p.n61 out_p.t2125 7.173
R31613 out_p.n60 out_p.t1707 7.173
R31614 out_p.n60 out_p.t2726 7.173
R31615 out_p.n59 out_p.t2366 7.173
R31616 out_p.n59 out_p.t2746 7.173
R31617 out_p.n58 out_p.t1164 7.173
R31618 out_p.n58 out_p.t1551 7.173
R31619 out_p.n57 out_p.t764 7.173
R31620 out_p.n57 out_p.t3413 7.173
R31621 out_p.n56 out_p.t1725 7.173
R31622 out_p.n56 out_p.t979 7.173
R31623 out_p.n55 out_p.t1812 7.173
R31624 out_p.n55 out_p.t2756 7.173
R31625 out_p.n54 out_p.t3287 7.173
R31626 out_p.n54 out_p.t1316 7.173
R31627 out_p.n53 out_p.t3034 7.173
R31628 out_p.n53 out_p.t1638 7.173
R31629 out_p.n52 out_p.t2629 7.173
R31630 out_p.n52 out_p.t1771 7.173
R31631 out_p.n51 out_p.t2047 7.173
R31632 out_p.n51 out_p.t2824 7.173
R31633 out_p.n50 out_p.t2347 7.173
R31634 out_p.n50 out_p.t2577 7.173
R31635 out_p.n49 out_p.t3305 7.173
R31636 out_p.n49 out_p.t780 7.173
R31637 out_p.n48 out_p.t3053 7.173
R31638 out_p.n48 out_p.t541 7.173
R31639 out_p.n43 out_p.t1952 7.173
R31640 out_p.n43 out_p.t2376 7.173
R31641 out_p.n42 out_p.t556 7.173
R31642 out_p.n42 out_p.t1292 7.173
R31643 out_p.n41 out_p.t808 7.173
R31644 out_p.n41 out_p.t618 7.173
R31645 out_p.n40 out_p.t3246 7.173
R31646 out_p.n40 out_p.t3055 7.173
R31647 out_p.n39 out_p.t2771 7.173
R31648 out_p.n39 out_p.t2574 7.173
R31649 out_p.n38 out_p.t1663 7.173
R31650 out_p.n38 out_p.t2465 7.173
R31651 out_p.n37 out_p.t725 7.173
R31652 out_p.n37 out_p.t545 7.173
R31653 out_p.n36 out_p.t1543 7.173
R31654 out_p.n36 out_p.t1810 7.173
R31655 out_p.n35 out_p.t566 7.173
R31656 out_p.n35 out_p.t2168 7.173
R31657 out_p.n34 out_p.t628 7.173
R31658 out_p.n34 out_p.t1184 7.173
R31659 out_p.n33 out_p.t2162 7.173
R31660 out_p.n33 out_p.t792 7.173
R31661 out_p.n32 out_p.t3376 7.173
R31662 out_p.n32 out_p.t1772 7.173
R31663 out_p.n31 out_p.t1585 7.173
R31664 out_p.n31 out_p.t1918 7.173
R31665 out_p.n30 out_p.t2714 7.173
R31666 out_p.n30 out_p.t3311 7.173
R31667 out_p.n29 out_p.t1144 7.173
R31668 out_p.n29 out_p.t3061 7.173
R31669 out_p.n28 out_p.t746 7.173
R31670 out_p.n28 out_p.t2654 7.173
R31671 out_p.n27 out_p.t1691 7.173
R31672 out_p.n27 out_p.t2138 7.173
R31673 out_p.n26 out_p.t2186 7.173
R31674 out_p.n26 out_p.t2385 7.173
R31675 out_p.n25 out_p.t1669 7.173
R31676 out_p.n25 out_p.t3285 7.173
R31677 out_p.n24 out_p.t3221 7.173
R31678 out_p.n24 out_p.t3030 7.173
R31679 out_p.n19 out_p.t2645 7.173
R31680 out_p.n19 out_p.t2706 7.173
R31681 out_p.n18 out_p.t3049 7.173
R31682 out_p.n18 out_p.t3137 7.173
R31683 out_p.n17 out_p.t3303 7.173
R31684 out_p.n17 out_p.t3367 7.173
R31685 out_p.n16 out_p.t1870 7.173
R31686 out_p.n16 out_p.t2139 7.173
R31687 out_p.n15 out_p.t1760 7.173
R31688 out_p.n15 out_p.t1913 7.173
R31689 out_p.n14 out_p.t783 7.173
R31690 out_p.n14 out_p.t858 7.173
R31691 out_p.n13 out_p.t3226 7.173
R31692 out_p.n13 out_p.t3312 7.173
R31693 out_p.n12 out_p.t1183 7.173
R31694 out_p.n12 out_p.t2170 7.173
R31695 out_p.n11 out_p.t3280 7.173
R31696 out_p.n11 out_p.t2791 7.173
R31697 out_p.n10 out_p.t1860 7.173
R31698 out_p.n10 out_p.t1297 7.173
R31699 out_p.n9 out_p.t3200 7.173
R31700 out_p.n9 out_p.t2263 7.173
R31701 out_p.n8 out_p.t753 7.173
R31702 out_p.n8 out_p.t3063 7.173
R31703 out_p.n7 out_p.t2528 7.173
R31704 out_p.n7 out_p.t1205 7.173
R31705 out_p.n6 out_p.t1742 7.173
R31706 out_p.n6 out_p.t1080 7.173
R31707 out_p.n5 out_p.t2190 7.173
R31708 out_p.n5 out_p.t854 7.173
R31709 out_p.n4 out_p.t1386 7.173
R31710 out_p.n4 out_p.t1266 7.173
R31711 out_p.n3 out_p.t2608 7.173
R31712 out_p.n3 out_p.t1823 7.173
R31713 out_p.n2 out_p.t1051 7.173
R31714 out_p.n2 out_p.t3361 7.173
R31715 out_p.n1 out_p.t2477 7.173
R31716 out_p.n1 out_p.t1255 7.173
R31717 out_p.n0 out_p.t1788 7.173
R31718 out_p.n0 out_p.t2065 7.173
R31719 out_p.n824 out_p.t2849 7.173
R31720 out_p.n824 out_p.t2337 7.173
R31721 out_p.n823 out_p.t3284 7.173
R31722 out_p.n823 out_p.t2484 7.173
R31723 out_p.n822 out_p.t1221 7.173
R31724 out_p.n822 out_p.t589 7.173
R31725 out_p.n821 out_p.t2513 7.173
R31726 out_p.n821 out_p.t3031 7.173
R31727 out_p.n820 out_p.t2217 7.173
R31728 out_p.n820 out_p.t2551 7.173
R31729 out_p.n819 out_p.t1013 7.173
R31730 out_p.n819 out_p.t2309 7.173
R31731 out_p.n818 out_p.t1196 7.173
R31732 out_p.n818 out_p.t532 7.173
R31733 out_p.n817 out_p.t3080 7.173
R31734 out_p.n817 out_p.t2218 7.173
R31735 out_p.n816 out_p.t2815 7.173
R31736 out_p.n816 out_p.t641 7.173
R31737 out_p.n815 out_p.t2227 7.173
R31738 out_p.n815 out_p.t980 7.173
R31739 out_p.n814 out_p.t1438 7.173
R31740 out_p.n814 out_p.t557 7.173
R31741 out_p.n813 out_p.t2639 7.173
R31742 out_p.n813 out_p.t2504 7.173
R31743 out_p.n812 out_p.t3112 7.173
R31744 out_p.n812 out_p.t2276 7.173
R31745 out_p.n811 out_p.t670 7.173
R31746 out_p.n811 out_p.t3068 7.173
R31747 out_p.n810 out_p.t1317 7.173
R31748 out_p.n810 out_p.t2828 7.173
R31749 out_p.n809 out_p.t1403 7.173
R31750 out_p.n809 out_p.t1087 7.173
R31751 out_p.n808 out_p.t3172 7.173
R31752 out_p.n808 out_p.t2395 7.173
R31753 out_p.n807 out_p.t2939 7.173
R31754 out_p.n807 out_p.t1912 7.173
R31755 out_p.n806 out_p.t568 7.173
R31756 out_p.n806 out_p.t3264 7.173
R31757 out_p.n805 out_p.t1295 7.173
R31758 out_p.n805 out_p.t3014 7.173
R31759 out_p.n844 out_p.t3028 7.173
R31760 out_p.n844 out_p.t1104 7.173
R31761 out_p.n843 out_p.t1456 7.173
R31762 out_p.n843 out_p.t2839 7.173
R31763 out_p.n842 out_p.t2294 7.173
R31764 out_p.n842 out_p.t3086 7.173
R31765 out_p.n841 out_p.t530 7.173
R31766 out_p.n841 out_p.t2305 7.173
R31767 out_p.n840 out_p.t1525 7.173
R31768 out_p.n840 out_p.t1398 7.173
R31769 out_p.n839 out_p.t1160 7.173
R31770 out_p.n839 out_p.t573 7.173
R31771 out_p.n838 out_p.t1907 7.173
R31772 out_p.n838 out_p.t3018 7.173
R31773 out_p.n837 out_p.t1187 7.173
R31774 out_p.n837 out_p.t2858 7.173
R31775 out_p.n836 out_p.t442 7.173
R31776 out_p.n836 out_p.t3346 7.173
R31777 out_p.n835 out_p.t1904 7.173
R31778 out_p.n835 out_p.t1781 7.173
R31779 out_p.n834 out_p.t3202 7.173
R31780 out_p.n834 out_p.t2344 7.173
R31781 out_p.n833 out_p.t758 7.173
R31782 out_p.n833 out_p.t1092 7.173
R31783 out_p.n832 out_p.t2534 7.173
R31784 out_p.n832 out_p.t2890 7.173
R31785 out_p.n831 out_p.t1763 7.173
R31786 out_p.n831 out_p.t1344 7.173
R31787 out_p.n830 out_p.t2200 7.173
R31788 out_p.n830 out_p.t2140 7.173
R31789 out_p.n829 out_p.t1408 7.173
R31790 out_p.n829 out_p.t2039 7.173
R31791 out_p.n828 out_p.t2617 7.173
R31792 out_p.n828 out_p.t2961 7.173
R31793 out_p.n827 out_p.t1055 7.173
R31794 out_p.n827 out_p.t2707 7.173
R31795 out_p.n826 out_p.t737 7.173
R31796 out_p.n826 out_p.t1942 7.173
R31797 out_p.n825 out_p.t508 7.173
R31798 out_p.n825 out_p.t2267 7.173
R31799 out_p.n868 out_p.t2297 7.173
R31800 out_p.n868 out_p.t3351 7.173
R31801 out_p.n867 out_p.t1291 7.173
R31802 out_p.n867 out_p.t1439 7.173
R31803 out_p.n866 out_p.t569 7.173
R31804 out_p.n866 out_p.t1876 7.173
R31805 out_p.n865 out_p.t3015 7.173
R31806 out_p.n865 out_p.t843 7.173
R31807 out_p.n864 out_p.t2529 7.173
R31808 out_p.n864 out_p.t1251 7.173
R31809 out_p.n863 out_p.t2184 7.173
R31810 out_p.n863 out_p.t2812 7.173
R31811 out_p.n862 out_p.t513 7.173
R31812 out_p.n862 out_p.t1734 7.173
R31813 out_p.n861 out_p.t2268 7.173
R31814 out_p.n861 out_p.t2174 7.173
R31815 out_p.n860 out_p.t535 7.173
R31816 out_p.n860 out_p.t2025 7.173
R31817 out_p.n859 out_p.t1003 7.173
R31818 out_p.n859 out_p.t2633 7.173
R31819 out_p.n858 out_p.t577 7.173
R31820 out_p.n858 out_p.t894 7.173
R31821 out_p.n857 out_p.t1412 7.173
R31822 out_p.n857 out_p.t1991 7.173
R31823 out_p.n856 out_p.t2318 7.173
R31824 out_p.n856 out_p.t2248 7.173
R31825 out_p.n855 out_p.t3092 7.173
R31826 out_p.n855 out_p.t3407 7.173
R31827 out_p.n854 out_p.t2841 7.173
R31828 out_p.n854 out_p.t3167 7.173
R31829 out_p.n853 out_p.t1110 7.173
R31830 out_p.n853 out_p.t2751 7.173
R31831 out_p.n852 out_p.t2468 7.173
R31832 out_p.n852 out_p.t1303 7.173
R31833 out_p.n851 out_p.t1948 7.173
R31834 out_p.n851 out_p.t1634 7.173
R31835 out_p.n850 out_p.t3240 7.173
R31836 out_p.n850 out_p.t1059 7.173
R31837 out_p.n849 out_p.t2994 7.173
R31838 out_p.n849 out_p.t823 7.173
R31839 out_p.n892 out_p.t1084 7.173
R31840 out_p.n892 out_p.t2211 7.173
R31841 out_p.n891 out_p.t2825 7.173
R31842 out_p.n891 out_p.t655 7.173
R31843 out_p.n890 out_p.t3067 7.173
R31844 out_p.n890 out_p.t884 7.173
R31845 out_p.n889 out_p.t2274 7.173
R31846 out_p.n889 out_p.t3339 7.173
R31847 out_p.n888 out_p.t2511 7.173
R31848 out_p.n888 out_p.t2847 7.173
R31849 out_p.n887 out_p.t555 7.173
R31850 out_p.n887 out_p.t1841 7.173
R31851 out_p.n886 out_p.t2998 7.173
R31852 out_p.n886 out_p.t832 7.173
R31853 out_p.n885 out_p.t2884 7.173
R31854 out_p.n885 out_p.t3206 7.173
R31855 out_p.n884 out_p.t3237 7.173
R31856 out_p.n884 out_p.t1158 7.173
R31857 out_p.n883 out_p.t1818 7.173
R31858 out_p.n883 out_p.t1362 7.173
R31859 out_p.n882 out_p.t1558 7.173
R31860 out_p.n882 out_p.t1631 7.173
R31861 out_p.n881 out_p.t1111 7.173
R31862 out_p.n881 out_p.t2757 7.173
R31863 out_p.n880 out_p.t2916 7.173
R31864 out_p.n880 out_p.t3233 7.173
R31865 out_p.n879 out_p.t475 7.173
R31866 out_p.n879 out_p.t790 7.173
R31867 out_p.n878 out_p.t2198 7.173
R31868 out_p.n878 out_p.t547 7.173
R31869 out_p.n877 out_p.t2095 7.173
R31870 out_p.n877 out_p.t1914 7.173
R31871 out_p.n876 out_p.t2979 7.173
R31872 out_p.n876 out_p.t3309 7.173
R31873 out_p.n875 out_p.t2734 7.173
R31874 out_p.n875 out_p.t3056 7.173
R31875 out_p.n874 out_p.t1850 7.173
R31876 out_p.n874 out_p.t1457 7.173
R31877 out_p.n873 out_p.t2228 7.173
R31878 out_p.n873 out_p.t3321 7.173
R31879 out_p.n916 out_p.t1718 7.173
R31880 out_p.n916 out_p.t2722 7.173
R31881 out_p.n915 out_p.t1877 7.173
R31882 out_p.n915 out_p.t3150 7.173
R31883 out_p.n914 out_p.t2368 7.173
R31884 out_p.n914 out_p.t3385 7.173
R31885 out_p.n913 out_p.t1073 7.173
R31886 out_p.n913 out_p.t2172 7.173
R31887 out_p.n912 out_p.t610 7.173
R31888 out_p.n912 out_p.t1934 7.173
R31889 out_p.n911 out_p.t3048 7.173
R31890 out_p.n911 out_p.t869 7.173
R31891 out_p.n910 out_p.t2240 7.173
R31892 out_p.n910 out_p.t3326 7.173
R31893 out_p.n909 out_p.t1278 7.173
R31894 out_p.n909 out_p.t581 7.173
R31895 out_p.n908 out_p.t1277 7.173
R31896 out_p.n908 out_p.t1627 7.173
R31897 out_p.n907 out_p.t2676 7.173
R31898 out_p.n907 out_p.t2991 7.173
R31899 out_p.n906 out_p.t954 7.173
R31900 out_p.n906 out_p.t2572 7.173
R31901 out_p.n905 out_p.t2119 7.173
R31902 out_p.n905 out_p.t1919 7.173
R31903 out_p.n904 out_p.t2450 7.173
R31904 out_p.n904 out_p.t612 7.173
R31905 out_p.n903 out_p.t1467 7.173
R31906 out_p.n903 out_p.t1466 7.173
R31907 out_p.n902 out_p.t3212 7.173
R31908 out_p.n902 out_p.t1206 7.173
R31909 out_p.n901 out_p.t2805 7.173
R31910 out_p.n901 out_p.t3130 7.173
R31911 out_p.n900 out_p.t1307 7.173
R31912 out_p.n900 out_p.t683 7.173
R31913 out_p.n899 out_p.t1833 7.173
R31914 out_p.n899 out_p.t1265 7.173
R31915 out_p.n898 out_p.t2622 7.173
R31916 out_p.n898 out_p.t1349 7.173
R31917 out_p.n897 out_p.t1060 7.173
R31918 out_p.n897 out_p.t2112 7.173
R31919 out_p.n940 out_p.t549 7.173
R31920 out_p.n940 out_p.t1678 7.173
R31921 out_p.n939 out_p.t973 7.173
R31922 out_p.n939 out_p.t1471 7.173
R31923 out_p.n938 out_p.t1185 7.173
R31924 out_p.n938 out_p.t1249 7.173
R31925 out_p.n937 out_p.t2078 7.173
R31926 out_p.n937 out_p.t2704 7.173
R31927 out_p.n936 out_p.t3176 7.173
R31928 out_p.n936 out_p.t926 7.173
R31929 out_p.n935 out_p.t1404 7.173
R31930 out_p.n935 out_p.t3366 7.173
R31931 out_p.n934 out_p.t1127 7.173
R31932 out_p.n934 out_p.t2136 7.173
R31933 out_p.n933 out_p.t899 7.173
R31934 out_p.n933 out_p.t1606 7.173
R31935 out_p.n932 out_p.t3140 7.173
R31936 out_p.n932 out_p.t989 7.173
R31937 out_p.n931 out_p.t3322 7.173
R31938 out_p.n931 out_p.t1293 7.173
R31939 out_p.n930 out_p.t2898 7.173
R31940 out_p.n930 out_p.t2377 7.173
R31941 out_p.n929 out_p.t2501 7.173
R31942 out_p.n929 out_p.t3132 7.173
R31943 out_p.n928 out_p.t936 7.173
R31944 out_p.n928 out_p.t1776 7.173
R31945 out_p.n927 out_p.t2063 7.173
R31946 out_p.n927 out_p.t1138 7.173
R31947 out_p.n926 out_p.t1588 7.173
R31948 out_p.n926 out_p.t910 7.173
R31949 out_p.n925 out_p.t445 7.173
R31950 out_p.n925 out_p.t505 7.173
R31951 out_p.n924 out_p.t1007 7.173
R31952 out_p.n924 out_p.t2148 7.173
R31953 out_p.n923 out_p.t752 7.173
R31954 out_p.n923 out_p.t3426 7.173
R31955 out_p.n922 out_p.t1617 7.173
R31956 out_p.n922 out_p.t2944 7.173
R31957 out_p.n921 out_p.t1986 7.173
R31958 out_p.n921 out_p.t2690 7.173
R31959 out_p.n964 out_p.t3045 7.173
R31960 out_p.n964 out_p.t2018 7.173
R31961 out_p.n963 out_p.t1508 7.173
R31962 out_p.n963 out_p.t2113 7.173
R31963 out_p.n962 out_p.t2372 7.173
R31964 out_p.n962 out_p.t1350 7.173
R31965 out_p.n961 out_p.t538 7.173
R31966 out_p.n961 out_p.t2879 7.173
R31967 out_p.n960 out_p.t1571 7.173
R31968 out_p.n960 out_p.t1081 7.173
R31969 out_p.n959 out_p.t1170 7.173
R31970 out_p.n959 out_p.t1203 7.173
R31971 out_p.n958 out_p.t2009 7.173
R31972 out_p.n958 out_p.t1289 7.173
R31973 out_p.n957 out_p.t1639 7.173
R31974 out_p.n957 out_p.t3011 7.173
R31975 out_p.n956 out_p.t2208 7.173
R31976 out_p.n956 out_p.t2911 7.173
R31977 out_p.n955 out_p.t692 7.173
R31978 out_p.n955 out_p.t2087 7.173
R31979 out_p.n954 out_p.t2406 7.173
R31980 out_p.n954 out_p.t2326 7.173
R31981 out_p.n953 out_p.t454 7.173
R31982 out_p.n953 out_p.t2555 7.173
R31983 out_p.n952 out_p.t1697 7.173
R31984 out_p.n952 out_p.t3035 7.173
R31985 out_p.n951 out_p.t2787 7.173
R31986 out_p.n951 out_p.t593 7.173
R31987 out_p.n950 out_p.t2532 7.173
R31988 out_p.n950 out_p.t2514 7.173
R31989 out_p.n949 out_p.t824 7.173
R31990 out_p.n949 out_p.t2338 7.173
R31991 out_p.n948 out_p.t1830 7.173
R31992 out_p.n948 out_p.t3105 7.173
R31993 out_p.n947 out_p.t1399 7.173
R31994 out_p.n947 out_p.t2850 7.173
R31995 out_p.n946 out_p.t756 7.173
R31996 out_p.n946 out_p.t3106 7.173
R31997 out_p.n945 out_p.t522 7.173
R31998 out_p.n945 out_p.t2851 7.173
R31999 out_p.n988 out_p.t2333 7.173
R32000 out_p.n988 out_p.t3022 7.173
R32001 out_p.n987 out_p.t1232 7.173
R32002 out_p.n987 out_p.t448 7.173
R32003 out_p.n986 out_p.t584 7.173
R32004 out_p.n986 out_p.t2270 7.173
R32005 out_p.n985 out_p.t3025 7.173
R32006 out_p.n985 out_p.t524 7.173
R32007 out_p.n984 out_p.t2545 7.173
R32008 out_p.n984 out_p.t1513 7.173
R32009 out_p.n983 out_p.t2273 7.173
R32010 out_p.n983 out_p.t1153 7.173
R32011 out_p.n982 out_p.t527 7.173
R32012 out_p.n982 out_p.t1883 7.173
R32013 out_p.n981 out_p.t2578 7.173
R32014 out_p.n981 out_p.t1687 7.173
R32015 out_p.n980 out_p.t2945 7.173
R32016 out_p.n980 out_p.t1869 7.173
R32017 out_p.n979 out_p.t2233 7.173
R32018 out_p.n979 out_p.t708 7.173
R32019 out_p.n978 out_p.t3271 7.173
R32020 out_p.n978 out_p.t2437 7.173
R32021 out_p.n977 out_p.t828 7.173
R32022 out_p.n977 out_p.t1645 7.173
R32023 out_p.n976 out_p.t2609 7.173
R32024 out_p.n976 out_p.t1735 7.173
R32025 out_p.n975 out_p.t2020 7.173
R32026 out_p.n975 out_p.t2813 7.173
R32027 out_p.n974 out_p.t2317 7.173
R32028 out_p.n974 out_p.t2559 7.173
R32029 out_p.n973 out_p.t1519 7.173
R32030 out_p.n973 out_p.t844 7.173
R32031 out_p.n972 out_p.t2679 7.173
R32032 out_p.n972 out_p.t1878 7.173
R32033 out_p.n971 out_p.t1106 7.173
R32034 out_p.n971 out_p.t1442 7.173
R32035 out_p.n970 out_p.t3257 7.173
R32036 out_p.n970 out_p.t732 7.173
R32037 out_p.n969 out_p.t3009 7.173
R32038 out_p.n969 out_p.t502 7.173
R32039 out_p.n1012 out_p.t1743 7.173
R32040 out_p.n1012 out_p.t2259 7.173
R32041 out_p.n1011 out_p.t519 7.173
R32042 out_p.n1011 out_p.t667 7.173
R32043 out_p.n1010 out_p.t754 7.173
R32044 out_p.n1010 out_p.t896 7.173
R32045 out_p.n1009 out_p.t3201 7.173
R32046 out_p.n1009 out_p.t3350 7.173
R32047 out_p.n1008 out_p.t2718 7.173
R32048 out_p.n1008 out_p.t2869 7.173
R32049 out_p.n1007 out_p.t1590 7.173
R32050 out_p.n1007 out_p.t1866 7.173
R32051 out_p.n1006 out_p.t691 7.173
R32052 out_p.n1006 out_p.t841 7.173
R32053 out_p.n1005 out_p.t704 7.173
R32054 out_p.n1005 out_p.t2399 7.173
R32055 out_p.n1004 out_p.t1482 7.173
R32056 out_p.n1004 out_p.t1649 7.173
R32057 out_p.n1003 out_p.t3127 7.173
R32058 out_p.n1003 out_p.t2686 7.173
R32059 out_p.n1002 out_p.t2699 7.173
R32060 out_p.n1002 out_p.t971 7.173
R32061 out_p.n1001 out_p.t1354 7.173
R32062 out_p.n1001 out_p.t2152 7.173
R32063 out_p.n1000 out_p.t726 7.173
R32064 out_p.n1000 out_p.t2488 7.173
R32065 out_p.n999 out_p.t1667 7.173
R32066 out_p.n999 out_p.t1715 7.173
R32067 out_p.n998 out_p.t2104 7.173
R32068 out_p.n998 out_p.t3227 7.173
R32069 out_p.n997 out_p.t3247 7.173
R32070 out_p.n997 out_p.t2817 7.173
R32071 out_p.n996 out_p.t809 7.173
R32072 out_p.n996 out_p.t1284 7.173
R32073 out_p.n995 out_p.t559 7.173
R32074 out_p.n995 out_p.t1892 7.173
R32075 out_p.n994 out_p.t3421 7.173
R32076 out_p.n994 out_p.t1559 7.173
R32077 out_p.n993 out_p.t3177 7.173
R32078 out_p.n993 out_p.t3332 7.173
R32079 out_p.n1036 out_p.t2588 7.173
R32080 out_p.n1036 out_p.t2448 7.173
R32081 out_p.n1035 out_p.t3005 7.173
R32082 out_p.n1035 out_p.t837 7.173
R32083 out_p.n1034 out_p.t3253 7.173
R32084 out_p.n1034 out_p.t1068 7.173
R32085 out_p.n1033 out_p.t1683 7.173
R32086 out_p.n1033 out_p.t1220 7.173
R32087 out_p.n1032 out_p.t1676 7.173
R32088 out_p.n1032 out_p.t3039 7.173
R32089 out_p.n1031 out_p.t734 7.173
R32090 out_p.n1031 out_p.t2213 7.173
R32091 out_p.n1030 out_p.t3182 7.173
R32092 out_p.n1030 out_p.t1012 7.173
R32093 out_p.n1029 out_p.t2370 7.173
R32094 out_p.n1029 out_p.t1899 7.173
R32095 out_p.n1028 out_p.t661 7.173
R32096 out_p.n1028 out_p.t2278 7.173
R32097 out_p.n1027 out_p.t503 7.173
R32098 out_p.n1027 out_p.t820 7.173
R32099 out_p.n1026 out_p.t1682 7.173
R32100 out_p.n1026 out_p.t1331 7.173
R32101 out_p.n1025 out_p.t3251 7.173
R32102 out_p.n1025 out_p.t1560 7.173
R32103 out_p.n1024 out_p.t2502 7.173
R32104 out_p.n1024 out_p.t1935 7.173
R32105 out_p.n1023 out_p.t2587 7.173
R32106 out_p.n1023 out_p.t2912 7.173
R32107 out_p.n1022 out_p.t1040 7.173
R32108 out_p.n1022 out_p.t2671 7.173
R32109 out_p.n1021 out_p.t629 7.173
R32110 out_p.n1021 out_p.t948 7.173
R32111 out_p.n1020 out_p.t1489 7.173
R32112 out_p.n1020 out_p.t2096 7.173
R32113 out_p.n1019 out_p.t1375 7.173
R32114 out_p.n1019 out_p.t1609 7.173
R32115 out_p.n1018 out_p.t2403 7.173
R32116 out_p.n1018 out_p.t1385 7.173
R32117 out_p.n1017 out_p.t1572 7.173
R32118 out_p.n1017 out_p.t1211 7.173
R32119 out_p.n1060 out_p.t2199 7.173
R32120 out_p.n1060 out_p.t2913 7.173
R32121 out_p.n1059 out_p.t647 7.173
R32122 out_p.n1059 out_p.t3333 7.173
R32123 out_p.n1058 out_p.t876 7.173
R32124 out_p.n1058 out_p.t1537 7.173
R32125 out_p.n1057 out_p.t3335 7.173
R32126 out_p.n1057 out_p.t1330 7.173
R32127 out_p.n1056 out_p.t2844 7.173
R32128 out_p.n1056 out_p.t2321 7.173
R32129 out_p.n1055 out_p.t1819 7.173
R32130 out_p.n1055 out_p.t1053 7.173
R32131 out_p.n1054 out_p.t821 7.173
R32132 out_p.n1054 out_p.t2031 7.173
R32133 out_p.n1053 out_p.t2474 7.173
R32134 out_p.n1053 out_p.t2702 7.173
R32135 out_p.n1052 out_p.t1785 7.173
R32136 out_p.n1052 out_p.t2616 7.173
R32137 out_p.n1051 out_p.t2703 7.173
R32138 out_p.n1051 out_p.t1516 7.173
R32139 out_p.n1050 out_p.t993 7.173
R32140 out_p.n1050 out_p.t3388 7.173
R32141 out_p.n1049 out_p.t2182 7.173
R32142 out_p.n1049 out_p.t955 7.173
R32143 out_p.n1048 out_p.t439 7.173
R32144 out_p.n1048 out_p.t2728 7.173
R32145 out_p.n1047 out_p.t1214 7.173
R32146 out_p.n1047 out_p.t2426 7.173
R32147 out_p.n1046 out_p.t3258 7.173
R32148 out_p.n1046 out_p.t1526 7.173
R32149 out_p.n1045 out_p.t2833 7.173
R32150 out_p.n1045 out_p.t1722 7.173
R32151 out_p.n1044 out_p.t2487 7.173
R32152 out_p.n1044 out_p.t2806 7.173
R32153 out_p.n1043 out_p.t1975 7.173
R32154 out_p.n1043 out_p.t2546 7.173
R32155 out_p.n1042 out_p.t1376 7.173
R32156 out_p.n1042 out_p.t627 7.173
R32157 out_p.n1041 out_p.t3316 7.173
R32158 out_p.n1041 out_p.t1334 7.173
R32159 out_p.n1084 out_p.t2985 7.173
R32160 out_p.n1084 out_p.t1066 7.173
R32161 out_p.n1083 out_p.t3398 7.173
R32162 out_p.n1083 out_p.t2803 7.173
R32163 out_p.n1082 out_p.t2056 7.173
R32164 out_p.n1082 out_p.t3040 7.173
R32165 out_p.n1081 out_p.t483 7.173
R32166 out_p.n1081 out_p.t2214 7.173
R32167 out_p.n1080 out_p.t2473 7.173
R32168 out_p.n1080 out_p.t2353 7.173
R32169 out_p.n1079 out_p.t1119 7.173
R32170 out_p.n1079 out_p.t536 7.173
R32171 out_p.n1078 out_p.t1624 7.173
R32172 out_p.n1078 out_p.t2973 7.173
R32173 out_p.n1077 out_p.t2389 7.173
R32174 out_p.n1077 out_p.t1956 7.173
R32175 out_p.n1076 out_p.t817 7.173
R32176 out_p.n1076 out_p.t712 7.173
R32177 out_p.n1075 out_p.t509 7.173
R32178 out_p.n1075 out_p.t849 7.173
R32179 out_p.n1074 out_p.t1706 7.173
R32180 out_p.n1074 out_p.t2490 7.173
R32181 out_p.n1073 out_p.t3259 7.173
R32182 out_p.n1073 out_p.t1777 7.173
R32183 out_p.n1072 out_p.t1368 7.173
R32184 out_p.n1072 out_p.t2002 7.173
R32185 out_p.n1071 out_p.t2592 7.173
R32186 out_p.n1071 out_p.t2948 7.173
R32187 out_p.n1070 out_p.t1045 7.173
R32188 out_p.n1070 out_p.t2696 7.173
R32189 out_p.n1069 out_p.t636 7.173
R32190 out_p.n1069 out_p.t981 7.173
R32191 out_p.n1068 out_p.t1502 7.173
R32192 out_p.n1068 out_p.t2165 7.173
R32193 out_p.n1067 out_p.t1418 7.173
R32194 out_p.n1067 out_p.t1652 7.173
R32195 out_p.n1066 out_p.t701 7.173
R32196 out_p.n1066 out_p.t1731 7.173
R32197 out_p.n1065 out_p.t460 7.173
R32198 out_p.n1065 out_p.t2188 7.173
R32199 out_p.n1108 out_p.t2161 7.173
R32200 out_p.n1108 out_p.t3313 7.173
R32201 out_p.n1107 out_p.t626 7.173
R32202 out_p.n1107 out_p.t1435 7.173
R32203 out_p.n1106 out_p.t861 7.173
R32204 out_p.n1106 out_p.t1779 7.173
R32205 out_p.n1105 out_p.t3317 7.173
R32206 out_p.n1105 out_p.t793 7.173
R32207 out_p.n1104 out_p.t2832 7.173
R32208 out_p.n1104 out_p.t1324 7.173
R32209 out_p.n1103 out_p.t1784 7.173
R32210 out_p.n1103 out_p.t2764 7.173
R32211 out_p.n1102 out_p.t801 7.173
R32212 out_p.n1102 out_p.t1641 7.173
R32213 out_p.n1101 out_p.t1635 7.173
R32214 out_p.n1101 out_p.t2705 7.173
R32215 out_p.n1100 out_p.t2409 7.173
R32216 out_p.n1100 out_p.t2772 7.173
R32217 out_p.n1099 out_p.t1145 7.173
R32218 out_p.n1099 out_p.t1520 7.173
R32219 out_p.n1098 out_p.t747 7.173
R32220 out_p.n1098 out_p.t3391 7.173
R32221 out_p.n1097 out_p.t1698 7.173
R32222 out_p.n1097 out_p.t960 7.173
R32223 out_p.n1096 out_p.t1730 7.173
R32224 out_p.n1096 out_p.t2736 7.173
R32225 out_p.n1095 out_p.t3268 7.173
R32226 out_p.n1095 out_p.t2447 7.173
R32227 out_p.n1094 out_p.t3019 7.173
R32228 out_p.n1094 out_p.t1548 7.173
R32229 out_p.n1093 out_p.t2605 7.173
R32230 out_p.n1093 out_p.t1732 7.173
R32231 out_p.n1092 out_p.t2000 7.173
R32232 out_p.n1092 out_p.t2811 7.173
R32233 out_p.n1091 out_p.t2302 7.173
R32234 out_p.n1091 out_p.t2556 7.173
R32235 out_p.n1090 out_p.t2388 7.173
R32236 out_p.n1090 out_p.t1022 7.173
R32237 out_p.n1089 out_p.t3295 7.173
R32238 out_p.n1089 out_p.t767 7.173
R32239 out_p.n1132 out_p.t2698 7.173
R32240 out_p.n1132 out_p.t2088 7.173
R32241 out_p.n1131 out_p.t3122 7.173
R32242 out_p.n1131 out_p.t602 7.173
R32243 out_p.n1130 out_p.t3357 7.173
R32244 out_p.n1130 out_p.t847 7.173
R32245 out_p.n1129 out_p.t2089 7.173
R32246 out_p.n1129 out_p.t3297 7.173
R32247 out_p.n1128 out_p.t1890 7.173
R32248 out_p.n1128 out_p.t2816 7.173
R32249 out_p.n1127 out_p.t852 7.173
R32250 out_p.n1127 out_p.t1750 7.173
R32251 out_p.n1126 out_p.t3301 7.173
R32252 out_p.n1126 out_p.t773 7.173
R32253 out_p.n1125 out_p.t3058 7.173
R32254 out_p.n1125 out_p.t1727 7.173
R32255 out_p.n1124 out_p.t2681 7.173
R32256 out_p.n1124 out_p.t2204 7.173
R32257 out_p.n1123 out_p.t2191 7.173
R32258 out_p.n1123 out_p.t1166 7.173
R32259 out_p.n1122 out_p.t1387 7.173
R32260 out_p.n1122 out_p.t768 7.173
R32261 out_p.n1121 out_p.t2610 7.173
R32262 out_p.n1121 out_p.t1736 7.173
R32263 out_p.n1120 out_p.t3081 7.173
R32264 out_p.n1120 out_p.t1845 7.173
R32265 out_p.n1119 out_p.t644 7.173
R32266 out_p.n1119 out_p.t3293 7.173
R32267 out_p.n1118 out_p.t1355 7.173
R32268 out_p.n1118 out_p.t3041 7.173
R32269 out_p.n1117 out_p.t2422 7.173
R32270 out_p.n1117 out_p.t2631 7.173
R32271 out_p.n1116 out_p.t3155 7.173
R32272 out_p.n1116 out_p.t2066 7.173
R32273 out_p.n1115 out_p.t2908 7.173
R32274 out_p.n1115 out_p.t2351 7.173
R32275 out_p.n1114 out_p.t2480 7.173
R32276 out_p.n1114 out_p.t2111 7.173
R32277 out_p.n1113 out_p.t2023 7.173
R32278 out_p.n1113 out_p.t3274 7.173
R32279 out_p.n1156 out_p.t2870 7.173
R32280 out_p.n1156 out_p.t2683 7.173
R32281 out_p.n1155 out_p.t3296 7.173
R32282 out_p.n1155 out_p.t3099 7.173
R32283 out_p.n1154 out_p.t2352 7.173
R32284 out_p.n1154 out_p.t3344 7.173
R32285 out_p.n1153 out_p.t1336 7.173
R32286 out_p.n1153 out_p.t2024 7.173
R32287 out_p.n1152 out_p.t2241 7.173
R32288 out_p.n1152 out_p.t1842 7.173
R32289 out_p.n1151 out_p.t1027 7.173
R32290 out_p.n1151 out_p.t836 7.173
R32291 out_p.n1150 out_p.t1557 7.173
R32292 out_p.n1150 out_p.t3278 7.173
R32293 out_p.n1149 out_p.t1165 7.173
R32294 out_p.n1149 out_p.t3077 7.173
R32295 out_p.n1148 out_p.t3306 7.173
R32296 out_p.n1148 out_p.t2566 7.173
R32297 out_p.n1147 out_p.t1719 7.173
R32298 out_p.n1147 out_p.t2226 7.173
R32299 out_p.n1146 out_p.t3178 7.173
R32300 out_p.n1146 out_p.t1431 7.173
R32301 out_p.n1145 out_p.t727 7.173
R32302 out_p.n1145 out_p.t2638 7.173
R32303 out_p.n1144 out_p.t1188 7.173
R32304 out_p.n1144 out_p.t3107 7.173
R32305 out_p.n1143 out_p.t1680 7.173
R32306 out_p.n1143 out_p.t668 7.173
R32307 out_p.n1142 out_p.t2164 7.173
R32308 out_p.n1142 out_p.t1305 7.173
R32309 out_p.n1141 out_p.t1437 7.173
R32310 out_p.n1141 out_p.t1363 7.173
R32311 out_p.n1140 out_p.t2585 7.173
R32312 out_p.n1140 out_p.t3170 7.173
R32313 out_p.n1139 out_p.t1038 7.173
R32314 out_p.n1139 out_p.t2936 7.173
R32315 out_p.n1138 out_p.t578 7.173
R32316 out_p.n1138 out_p.t1358 7.173
R32317 out_p.n1137 out_p.t1248 7.173
R32318 out_p.n1137 out_p.t1976 7.173
R32319 out_p.n1180 out_p.t514 7.173
R32320 out_p.n1180 out_p.t3194 7.173
R32321 out_p.n1179 out_p.t921 7.173
R32322 out_p.n1179 out_p.t1824 7.173
R32323 out_p.n1178 out_p.t1142 7.173
R32324 out_p.n1178 out_p.t1574 7.173
R32325 out_p.n1177 out_p.t1858 7.173
R32326 out_p.n1177 out_p.t686 7.173
R32327 out_p.n1176 out_p.t3138 7.173
R32328 out_p.n1176 out_p.t2158 7.173
R32329 out_p.n1175 out_p.t2387 7.173
R32330 out_p.n1175 out_p.t2655 7.173
R32331 out_p.n1174 out_p.t1082 7.173
R32332 out_p.n1174 out_p.t1475 7.173
R32333 out_p.n1173 out_p.t3394 7.173
R32334 out_p.n1173 out_p.t2092 7.173
R32335 out_p.n1172 out_p.t518 7.173
R32336 out_p.n1172 out_p.t1749 7.173
R32337 out_p.n1171 out_p.t2114 7.173
R32338 out_p.n1171 out_p.t2601 7.173
R32339 out_p.n1170 out_p.t2026 7.173
R32340 out_p.n1170 out_p.t871 7.173
R32341 out_p.n1169 out_p.t2955 7.173
R32342 out_p.n1169 out_p.t1936 7.173
R32343 out_p.n1168 out_p.t3427 7.173
R32344 out_p.n1168 out_p.t2175 7.173
R32345 out_p.n1167 out_p.t991 7.173
R32346 out_p.n1167 out_p.t3386 7.173
R32347 out_p.n1166 out_p.t733 7.173
R32348 out_p.n1166 out_p.t3152 7.173
R32349 out_p.n1165 out_p.t1340 7.173
R32350 out_p.n1165 out_p.t2723 7.173
R32351 out_p.n1164 out_p.t1903 7.173
R32352 out_p.n1164 out_p.t2446 7.173
R32353 out_p.n1163 out_p.t3252 7.173
R32354 out_p.n1163 out_p.t1523 7.173
R32355 out_p.n1162 out_p.t1544 7.173
R32356 out_p.n1162 out_p.t895 7.173
R32357 out_p.n1161 out_p.t1693 7.173
R32358 out_p.n1161 out_p.t665 7.173
R32359 out_p.n1204 out_p.t2999 7.173
R32360 out_p.n1204 out_p.t1657 7.173
R32361 out_p.n1203 out_p.t3414 7.173
R32362 out_p.n1203 out_p.t495 7.173
R32363 out_p.n1202 out_p.t2101 7.173
R32364 out_p.n1202 out_p.t722 7.173
R32365 out_p.n1201 out_p.t498 7.173
R32366 out_p.n1201 out_p.t3173 7.173
R32367 out_p.n1200 out_p.t1445 7.173
R32368 out_p.n1200 out_p.t2697 7.173
R32369 out_p.n1199 out_p.t1133 7.173
R32370 out_p.n1199 out_p.t1552 7.173
R32371 out_p.n1198 out_p.t1696 7.173
R32372 out_p.n1198 out_p.t671 7.173
R32373 out_p.n1197 out_p.t774 7.173
R32374 out_p.n1197 out_p.t3183 7.173
R32375 out_p.n1196 out_p.t3218 7.173
R32376 out_p.n1196 out_p.t1041 7.173
R32377 out_p.n1195 out_p.t3188 7.173
R32378 out_p.n1195 out_p.t2421 7.173
R32379 out_p.n1194 out_p.t2773 7.173
R32380 out_p.n1194 out_p.t1602 7.173
R32381 out_p.n1193 out_p.t1247 7.173
R32382 out_p.n1193 out_p.t2729 7.173
R32383 out_p.n1192 out_p.t810 7.173
R32384 out_p.n1192 out_p.t3207 7.173
R32385 out_p.n1191 out_p.t1796 7.173
R32386 out_p.n1191 out_p.t763 7.173
R32387 out_p.n1190 out_p.t1366 7.173
R32388 out_p.n1190 out_p.t531 7.173
R32389 out_p.n1189 out_p.t3323 7.173
R32390 out_p.n1189 out_p.t1789 7.173
R32391 out_p.n1188 out_p.t865 7.173
R32392 out_p.n1188 out_p.t3281 7.173
R32393 out_p.n1187 out_p.t633 7.173
R32394 out_p.n1187 out_p.t3029 7.173
R32395 out_p.n1186 out_p.t706 7.173
R32396 out_p.n1186 out_p.t3392 7.173
R32397 out_p.n1185 out_p.t476 7.173
R32398 out_p.n1185 out_p.t3158 7.173
R32399 out_p.n1228 out_p.t3169 7.173
R32400 out_p.n1228 out_p.t3327 7.173
R32401 out_p.n1227 out_p.t1672 7.173
R32402 out_p.n1227 out_p.t1380 7.173
R32403 out_p.n1226 out_p.t1541 7.173
R32404 out_p.n1226 out_p.t1804 7.173
R32405 out_p.n1225 out_p.t666 7.173
R32406 out_p.n1225 out_p.t813 7.173
R32407 out_p.n1224 out_p.t2067 7.173
R32408 out_p.n1224 out_p.t1283 7.173
R32409 out_p.n1223 out_p.t2636 7.173
R32410 out_p.n1223 out_p.t2779 7.173
R32411 out_p.n1222 out_p.t1428 7.173
R32412 out_p.n1222 out_p.t1677 7.173
R32413 out_p.n1221 out_p.t2173 7.173
R32414 out_p.n1221 out_p.t2030 7.173
R32415 out_p.n1220 out_p.t1564 7.173
R32416 out_p.n1220 out_p.t1601 7.173
R32417 out_p.n1219 out_p.t2630 7.173
R32418 out_p.n1219 out_p.t875 7.173
R32419 out_p.n1218 out_p.t892 7.173
R32420 out_p.n1218 out_p.t471 7.173
R32421 out_p.n1217 out_p.t1983 7.173
R32422 out_p.n1217 out_p.t2010 7.173
R32423 out_p.n1216 out_p.t2246 7.173
R32424 out_p.n1216 out_p.t2097 7.173
R32425 out_p.n1215 out_p.t3405 7.173
R32426 out_p.n1215 out_p.t2980 7.173
R32427 out_p.n1214 out_p.t3164 7.173
R32428 out_p.n1214 out_p.t2735 7.173
R32429 out_p.n1213 out_p.t2748 7.173
R32430 out_p.n1213 out_p.t1016 7.173
R32431 out_p.n1212 out_p.t1296 7.173
R32432 out_p.n1212 out_p.t2229 7.173
R32433 out_p.n1211 out_p.t1593 7.173
R32434 out_p.n1211 out_p.t1724 7.173
R32435 out_p.n1210 out_p.t872 7.173
R32436 out_p.n1210 out_p.t1034 7.173
R32437 out_p.n1209 out_p.t645 7.173
R32438 out_p.n1209 out_p.t784 7.173
R32439 out_p.n1252 out_p.t1549 7.173
R32440 out_p.n1252 out_p.t1880 7.173
R32441 out_p.n1251 out_p.t472 7.173
R32442 out_p.n1251 out_p.t1664 7.173
R32443 out_p.n1250 out_p.t705 7.173
R32444 out_p.n1250 out_p.t2178 7.173
R32445 out_p.n1249 out_p.t3159 7.173
R32446 out_p.n1249 out_p.t987 7.173
R32447 out_p.n1248 out_p.t2682 7.173
R32448 out_p.n1248 out_p.t510 7.173
R32449 out_p.n1247 out_p.t1529 7.173
R32450 out_p.n1247 out_p.t2952 7.173
R32451 out_p.n1246 out_p.t649 7.173
R32452 out_p.n1246 out_p.t2014 7.173
R32453 out_p.n1245 out_p.t3203 7.173
R32454 out_p.n1245 out_p.t2291 7.173
R32455 out_p.n1244 out_p.t940 7.173
R32456 out_p.n1244 out_p.t2070 7.173
R32457 out_p.n1243 out_p.t1360 7.173
R32458 out_p.n1243 out_p.t1335 7.173
R32459 out_p.n1242 out_p.t1629 7.173
R32460 out_p.n1242 out_p.t2287 7.173
R32461 out_p.n1241 out_p.t2753 7.173
R32462 out_p.n1241 out_p.t3076 7.173
R32463 out_p.n1240 out_p.t3228 7.173
R32464 out_p.n1240 out_p.t1393 7.173
R32465 out_p.n1239 out_p.t785 7.173
R32466 out_p.n1239 out_p.t1096 7.173
R32467 out_p.n1238 out_p.t544 7.173
R32468 out_p.n1238 out_p.t860 7.173
R32469 out_p.n1237 out_p.t1893 7.173
R32470 out_p.n1237 out_p.t1346 7.173
R32471 out_p.n1236 out_p.t3307 7.173
R32472 out_p.n1236 out_p.t1884 7.173
R32473 out_p.n1235 out_p.t3054 7.173
R32474 out_p.n1235 out_p.t3372 7.173
R32475 out_p.n1234 out_p.t3373 7.173
R32476 out_p.n1234 out_p.t1176 7.173
R32477 out_p.n1233 out_p.t3139 7.173
R32478 out_p.n1233 out_p.t964 7.173
R32479 out_p.n1276 out_p.t2538 7.173
R32480 out_p.n1276 out_p.t1285 7.173
R32481 out_p.n1275 out_p.t2966 7.173
R32482 out_p.n1275 out_p.t786 7.173
R32483 out_p.n1274 out_p.t3204 7.173
R32484 out_p.n1274 out_p.t1033 7.173
R32485 out_p.n1273 out_p.t1512 7.173
R32486 out_p.n1273 out_p.t1692 7.173
R32487 out_p.n1272 out_p.t1600 7.173
R32488 out_p.n1272 out_p.t2995 7.173
R32489 out_p.n1271 out_p.t697 7.173
R32490 out_p.n1271 out_p.t2145 7.173
R32491 out_p.n1270 out_p.t3142 7.173
R32492 out_p.n1270 out_p.t968 7.173
R32493 out_p.n1269 out_p.t579 7.173
R32494 out_p.n1269 out_p.t897 7.173
R32495 out_p.n1268 out_p.t2033 7.173
R32496 out_p.n1268 out_p.t2891 7.173
R32497 out_p.n1267 out_p.t2989 7.173
R32498 out_p.n1267 out_p.t3319 7.173
R32499 out_p.n1266 out_p.t2570 7.173
R32500 out_p.n1266 out_p.t2894 7.173
R32501 out_p.n1265 out_p.t1915 7.173
R32502 out_p.n1265 out_p.t2498 7.173
R32503 out_p.n1264 out_p.t611 7.173
R32504 out_p.n1264 out_p.t930 7.173
R32505 out_p.n1263 out_p.t1465 7.173
R32506 out_p.n1263 out_p.t2053 7.173
R32507 out_p.n1262 out_p.t1199 7.173
R32508 out_p.n1262 out_p.t1586 7.173
R32509 out_p.n1261 out_p.t3128 7.173
R32510 out_p.n1261 out_p.t428 7.173
R32511 out_p.n1260 out_p.t681 7.173
R32512 out_p.n1260 out_p.t1004 7.173
R32513 out_p.n1259 out_p.t2493 7.173
R32514 out_p.n1259 out_p.t750 7.173
R32515 out_p.n1258 out_p.t457 7.173
R32516 out_p.n1258 out_p.t2311 7.173
R32517 out_p.n1257 out_p.t1447 7.173
R32518 out_p.n1257 out_p.t1195 7.173
R32519 out_p.n1300 out_p.t1517 7.173
R32520 out_p.n1300 out_p.t2859 7.173
R32521 out_p.n1299 out_p.t2314 7.173
R32522 out_p.n1299 out_p.t3288 7.173
R32523 out_p.n1298 out_p.t2001 7.173
R32524 out_p.n1298 out_p.t2255 7.173
R32525 out_p.n1297 out_p.t2606 7.173
R32526 out_p.n1297 out_p.t1306 7.173
R32527 out_p.n1296 out_p.t826 7.173
R32528 out_p.n1296 out_p.t2231 7.173
R32529 out_p.n1295 out_p.t3269 7.173
R32530 out_p.n1295 out_p.t1018 7.173
R32531 out_p.n1294 out_p.t1739 7.173
R32532 out_p.n1294 out_p.t1197 7.173
R32533 out_p.n1293 out_p.t2524 7.173
R32534 out_p.n1293 out_p.t1632 7.173
R32535 out_p.n1292 out_p.t838 7.173
R32536 out_p.n1292 out_p.t2459 7.173
R32537 out_p.n1291 out_p.t1987 7.173
R32538 out_p.n1291 out_p.t689 7.173
R32539 out_p.n1290 out_p.t3214 7.173
R32540 out_p.n1290 out_p.t1222 7.173
R32541 out_p.n1289 out_p.t769 7.173
R32542 out_p.n1289 out_p.t447 7.173
R32543 out_p.n1288 out_p.t2550 7.173
R32544 out_p.n1288 out_p.t1690 7.173
R32545 out_p.n1287 out_p.t1834 7.173
R32546 out_p.n1287 out_p.t2785 7.173
R32547 out_p.n1286 out_p.t2205 7.173
R32548 out_p.n1286 out_p.t2531 7.173
R32549 out_p.n1285 out_p.t1426 7.173
R32550 out_p.n1285 out_p.t819 7.173
R32551 out_p.n1284 out_p.t2632 7.173
R32552 out_p.n1284 out_p.t1820 7.173
R32553 out_p.n1283 out_p.t1067 7.173
R32554 out_p.n1283 out_p.t1388 7.173
R32555 out_p.n1282 out_p.t2830 7.173
R32556 out_p.n1282 out_p.t574 7.173
R32557 out_p.n1281 out_p.t2580 7.173
R32558 out_p.n1281 out_p.t1276 7.173
R32559 out_p.n1324 out_p.t690 7.173
R32560 out_p.n1324 out_p.t3032 7.173
R32561 out_p.n1323 out_p.t1088 7.173
R32562 out_p.n1323 out_p.t1480 7.173
R32563 out_p.n1322 out_p.t2666 7.173
R32564 out_p.n1322 out_p.t2310 7.173
R32565 out_p.n1321 out_p.t1487 7.173
R32566 out_p.n1321 out_p.t533 7.173
R32567 out_p.n1320 out_p.t3324 7.173
R32568 out_p.n1320 out_p.t1546 7.173
R32569 out_p.n1319 out_p.t1953 7.173
R32570 out_p.n1319 out_p.t1162 7.173
R32571 out_p.n1318 out_p.t2586 7.173
R32572 out_p.n1318 out_p.t1965 7.173
R32573 out_p.n1317 out_p.t2289 7.173
R32574 out_p.n1317 out_p.t3337 7.173
R32575 out_p.n1316 out_p.t1219 7.173
R32576 out_p.n1316 out_p.t613 7.173
R32577 out_p.n1315 out_p.t1014 7.173
R32578 out_p.n1315 out_p.t1871 7.173
R32579 out_p.n1314 out_p.t591 7.173
R32580 out_p.n1314 out_p.t1887 7.173
R32581 out_p.n1313 out_p.t1429 7.173
R32582 out_p.n1313 out_p.t2877 7.173
R32583 out_p.n1312 out_p.t2339 7.173
R32584 out_p.n1312 out_p.t3355 7.173
R32585 out_p.n1311 out_p.t3108 7.173
R32586 out_p.n1311 out_p.t906 7.173
R32587 out_p.n1310 out_p.t2852 7.173
R32588 out_p.n1310 out_p.t672 7.173
R32589 out_p.n1309 out_p.t1121 7.173
R32590 out_p.n1309 out_p.t451 7.173
R32591 out_p.n1308 out_p.t1364 7.173
R32592 out_p.n1308 out_p.t3423 7.173
R32593 out_p.n1307 out_p.t1972 7.173
R32594 out_p.n1307 out_p.t3180 7.173
R32595 out_p.n1306 out_p.t1886 7.173
R32596 out_p.n1306 out_p.t741 7.173
R32597 out_p.n1305 out_p.t1452 7.173
R32598 out_p.n1305 out_p.t512 7.173
R32599 out_p.n1348 out_p.t3184 7.173
R32600 out_p.n1348 out_p.t3266 7.173
R32601 out_p.n1347 out_p.t1755 7.173
R32602 out_p.n1347 out_p.t2185 7.173
R32603 out_p.n1346 out_p.t1566 7.173
R32604 out_p.n1346 out_p.t1688 7.173
R32605 out_p.n1345 out_p.t676 7.173
R32606 out_p.n1345 out_p.t742 7.173
R32607 out_p.n1344 out_p.t2116 7.173
R32608 out_p.n1344 out_p.t1228 7.173
R32609 out_p.n1343 out_p.t2648 7.173
R32610 out_p.n1343 out_p.t2710 7.173
R32611 out_p.n1342 out_p.t1463 7.173
R32612 out_p.n1342 out_p.t1577 7.173
R32613 out_p.n1341 out_p.t2899 7.173
R32614 out_p.n1341 out_p.t1643 7.173
R32615 out_p.n1340 out_p.t642 7.173
R32616 out_p.n1340 out_p.t1954 7.173
R32617 out_p.n1339 out_p.t1852 7.173
R32618 out_p.n1339 out_p.t695 7.173
R32619 out_p.n1338 out_p.t1670 7.173
R32620 out_p.n1338 out_p.t2400 7.173
R32621 out_p.n1337 out_p.t1125 7.173
R32622 out_p.n1337 out_p.t1372 7.173
R32623 out_p.n1336 out_p.t2933 7.173
R32624 out_p.n1336 out_p.t1710 7.173
R32625 out_p.n1335 out_p.t490 7.173
R32626 out_p.n1335 out_p.t2792 7.173
R32627 out_p.n1334 out_p.t2223 7.173
R32628 out_p.n1334 out_p.t2537 7.173
R32629 out_p.n1333 out_p.t2134 7.173
R32630 out_p.n1333 out_p.t829 7.173
R32631 out_p.n1332 out_p.t2990 7.173
R32632 out_p.n1332 out_p.t1839 7.173
R32633 out_p.n1331 out_p.t2747 7.173
R32634 out_p.n1331 out_p.t1411 7.173
R32635 out_p.n1330 out_p.t889 7.173
R32636 out_p.n1330 out_p.t977 7.173
R32637 out_p.n1329 out_p.t658 7.173
R32638 out_p.n1329 out_p.t718 7.173
R32639 out_p.n1372 out_p.t1314 7.173
R32640 out_p.n1372 out_p.t489 7.173
R32641 out_p.n1371 out_p.t740 7.173
R32642 out_p.n1371 out_p.t887 7.173
R32643 out_p.n1370 out_p.t996 7.173
R32644 out_p.n1370 out_p.t1122 7.173
R32645 out_p.n1369 out_p.t441 7.173
R32646 out_p.n1369 out_p.t1647 7.173
R32647 out_p.n1368 out_p.t2962 7.173
R32648 out_p.n1368 out_p.t3109 7.173
R32649 out_p.n1367 out_p.t2040 7.173
R32650 out_p.n1367 out_p.t2340 7.173
R32651 out_p.n1366 out_p.t922 7.173
R32652 out_p.n1366 out_p.t1064 7.173
R32653 out_p.n1365 out_p.t693 7.173
R32654 out_p.n1365 out_p.t1357 7.173
R32655 out_p.n1364 out_p.t1646 7.173
R32656 out_p.n1364 out_p.t1825 7.173
R32657 out_p.n1363 out_p.t3100 7.173
R32658 out_p.n1363 out_p.t2672 7.173
R32659 out_p.n1362 out_p.t2684 7.173
R32660 out_p.n1362 out_p.t949 7.173
R32661 out_p.n1361 out_p.t2224 7.173
R32662 out_p.n1361 out_p.t2098 7.173
R32663 out_p.n1360 out_p.t711 7.173
R32664 out_p.n1360 out_p.t2439 7.173
R32665 out_p.n1359 out_p.t1628 7.173
R32666 out_p.n1359 out_p.t1193 7.173
R32667 out_p.n1358 out_p.t2034 7.173
R32668 out_p.n1358 out_p.t3209 7.173
R32669 out_p.n1357 out_p.t3225 7.173
R32670 out_p.n1357 out_p.t2800 7.173
R32671 out_p.n1356 out_p.t781 7.173
R32672 out_p.n1356 out_p.t2476 7.173
R32673 out_p.n1355 out_p.t542 7.173
R32674 out_p.n1355 out_p.t1811 7.173
R32675 out_p.n1354 out_p.t2079 7.173
R32676 out_p.n1354 out_p.t1507 7.173
R32677 out_p.n1353 out_p.t3409 7.173
R32678 out_p.n1353 out_p.t1484 7.173
R32679 out_p.n1396 out_p.t2829 7.173
R32680 out_p.n1396 out_p.t656 7.173
R32681 out_p.n1395 out_p.t3243 7.173
R32682 out_p.n1395 out_p.t1061 7.173
R32683 out_p.n1394 out_p.t1821 7.173
R32684 out_p.n1394 out_p.t2624 7.173
R32685 out_p.n1393 out_p.t1321 7.173
R32686 out_p.n1393 out_p.t1420 7.173
R32687 out_p.n1392 out_p.t2166 7.173
R32688 out_p.n1392 out_p.t3282 7.173
R32689 out_p.n1391 out_p.t982 7.173
R32690 out_p.n1391 out_p.t1790 7.173
R32691 out_p.n1390 out_p.t3415 7.173
R32692 out_p.n1390 out_p.t2542 7.173
R32693 out_p.n1389 out_p.t2234 7.173
R32694 out_p.n1389 out_p.t1856 7.173
R32695 out_p.n1388 out_p.t682 7.173
R32696 out_p.n1388 out_p.t2322 7.173
R32697 out_p.n1387 out_p.t484 7.173
R32698 out_p.n1387 out_p.t796 7.173
R32699 out_p.n1386 out_p.t1573 7.173
R32700 out_p.n1386 out_p.t1243 7.173
R32701 out_p.n1385 out_p.t3229 7.173
R32702 out_p.n1385 out_p.t1391 7.173
R32703 out_p.n1384 out_p.t2390 7.173
R32704 out_p.n1384 out_p.t1910 7.173
R32705 out_p.n1383 out_p.t2567 7.173
R32706 out_p.n1383 out_p.t2892 7.173
R32707 out_p.n1382 out_p.t1031 7.173
R32708 out_p.n1382 out_p.t2660 7.173
R32709 out_p.n1381 out_p.t604 7.173
R32710 out_p.n1381 out_p.t927 7.173
R32711 out_p.n1380 out_p.t1461 7.173
R32712 out_p.n1380 out_p.t2051 7.173
R32713 out_p.n1379 out_p.t2369 7.173
R32714 out_p.n1379 out_p.t1578 7.173
R32715 out_p.n1378 out_p.t539 7.173
R32716 out_p.n1378 out_p.t1803 7.173
R32717 out_p.n1377 out_p.t2451 7.173
R32718 out_p.n1377 out_p.t1371 7.173
R32719 out_p.n1420 out_p.t465 7.173
R32720 out_p.n1420 out_p.t3151 7.173
R32721 out_p.n1419 out_p.t870 7.173
R32722 out_p.n1419 out_p.t1483 7.173
R32723 out_p.n1418 out_p.t1103 7.173
R32724 out_p.n1418 out_p.t1515 7.173
R32725 out_p.n1417 out_p.t1498 7.173
R32726 out_p.n1417 out_p.t643 7.173
R32727 out_p.n1416 out_p.t3084 7.173
R32728 out_p.n1416 out_p.t1997 7.173
R32729 out_p.n1415 out_p.t2303 7.173
R32730 out_p.n1415 out_p.t2602 7.173
R32731 out_p.n1414 out_p.t1048 7.173
R32732 out_p.n1414 out_p.t1381 7.173
R32733 out_p.n1413 out_p.t2436 7.173
R32734 out_p.n1413 out_p.t2687 7.173
R32735 out_p.n1412 out_p.t2054 7.173
R32736 out_p.n1412 out_p.t2642 7.173
R32737 out_p.n1411 out_p.t2691 7.173
R32738 out_p.n1411 out_p.t1479 7.173
R32739 out_p.n1410 out_p.t974 7.173
R32740 out_p.n1410 out_p.t3368 7.173
R32741 out_p.n1409 out_p.t2155 7.173
R32742 out_p.n1409 out_p.t931 7.173
R32743 out_p.n1408 out_p.t2492 7.173
R32744 out_p.n1408 out_p.t2708 7.173
R32745 out_p.n1407 out_p.t1751 7.173
R32746 out_p.n1407 out_p.t1231 7.173
R32747 out_p.n1406 out_p.t3234 7.173
R32748 out_p.n1406 out_p.t1472 7.173
R32749 out_p.n1405 out_p.t2821 7.173
R32750 out_p.n1405 out_p.t1679 7.173
R32751 out_p.n1404 out_p.t1323 7.173
R32752 out_p.n1404 out_p.t2780 7.173
R32753 out_p.n1403 out_p.t1916 7.173
R32754 out_p.n1403 out_p.t2526 7.173
R32755 out_p.n1402 out_p.t1478 7.173
R32756 out_p.n1402 out_p.t856 7.173
R32757 out_p.n1401 out_p.t1218 7.173
R32758 out_p.n1401 out_p.t619 7.173
R32759 out_p.n1444 out_p.t638 7.173
R32760 out_p.n1444 out_p.t1473 7.173
R32761 out_p.n1443 out_p.t1046 7.173
R32762 out_p.n1443 out_p.t1342 7.173
R32763 out_p.n1442 out_p.t2595 7.173
R32764 out_p.n1442 out_p.t688 7.173
R32765 out_p.n1441 out_p.t1377 7.173
R32766 out_p.n1441 out_p.t3136 7.173
R32767 out_p.n1440 out_p.t3262 7.173
R32768 out_p.n1440 out_p.t2661 7.173
R32769 out_p.n1439 out_p.t1708 7.173
R32770 out_p.n1439 out_p.t1485 7.173
R32771 out_p.n1438 out_p.t2523 7.173
R32772 out_p.n1438 out_p.t625 7.173
R32773 out_p.n1437 out_p.t1901 7.173
R32774 out_p.n1437 out_p.t1595 7.173
R32775 out_p.n1436 out_p.t2132 7.173
R32776 out_p.n1436 out_p.t1920 7.173
R32777 out_p.n1435 out_p.t825 7.173
R32778 out_p.n1435 out_p.t1143 7.173
R32779 out_p.n1434 out_p.t1339 7.173
R32780 out_p.n1434 out_p.t743 7.173
R32781 out_p.n1433 out_p.t1581 7.173
R32782 out_p.n1433 out_p.t1689 7.173
R32783 out_p.n1432 out_p.t1947 7.173
R32784 out_p.n1432 out_p.t1728 7.173
R32785 out_p.n1431 out_p.t2920 7.173
R32786 out_p.n1431 out_p.t3267 7.173
R32787 out_p.n1430 out_p.t2674 7.173
R32788 out_p.n1430 out_p.t3016 7.173
R32789 out_p.n1429 out_p.t956 7.173
R32790 out_p.n1429 out_p.t2603 7.173
R32791 out_p.n1428 out_p.t2118 7.173
R32792 out_p.n1428 out_p.t1998 7.173
R32793 out_p.n1427 out_p.t1612 7.173
R32794 out_p.n1427 out_p.t2300 7.173
R32795 out_p.n1426 out_p.t1761 7.173
R32796 out_p.n1426 out_p.t3352 7.173
R32797 out_p.n1425 out_p.t2418 7.173
R32798 out_p.n1425 out_p.t3113 7.173
R32799 out_p.n1468 out_p.t1580 7.173
R32800 out_p.n1468 out_p.t957 7.173
R32801 out_p.n1467 out_p.t1620 7.173
R32802 out_p.n1467 out_p.t2677 7.173
R32803 out_p.n1466 out_p.t2130 7.173
R32804 out_p.n1466 out_p.t2923 7.173
R32805 out_p.n1465 out_p.t961 7.173
R32806 out_p.n1465 out_p.t1957 7.173
R32807 out_p.n1464 out_p.t485 7.173
R32808 out_p.n1464 out_p.t1604 7.173
R32809 out_p.n1463 out_p.t2927 7.173
R32810 out_p.n1463 out_p.t1252 7.173
R32811 out_p.n1462 out_p.t1961 7.173
R32812 out_p.n1462 out_p.t2842 7.173
R32813 out_p.n1461 out_p.t1234 7.173
R32814 out_p.n1461 out_p.t3026 7.173
R32815 out_p.n1460 out_p.t3286 7.173
R32816 out_p.n1460 out_p.t473 7.173
R32817 out_p.n1459 out_p.t2797 7.173
R32818 out_p.n1459 out_p.t2144 7.173
R32819 out_p.n1458 out_p.t1065 7.173
R32820 out_p.n1458 out_p.t2466 7.173
R32821 out_p.n1457 out_p.t2341 7.173
R32822 out_p.n1457 out_p.t2575 7.173
R32823 out_p.n1456 out_p.t2479 7.173
R32824 out_p.n1456 out_p.t3057 7.173
R32825 out_p.n1455 out_p.t1626 7.173
R32826 out_p.n1455 out_p.t620 7.173
R32827 out_p.n1454 out_p.t3341 7.173
R32828 out_p.n1454 out_p.t1288 7.173
R32829 out_p.n1453 out_p.t2929 7.173
R32830 out_p.n1453 out_p.t2378 7.173
R32831 out_p.n1452 out_p.t487 7.173
R32832 out_p.n1452 out_p.t3133 7.173
R32833 out_p.n1451 out_p.t2220 7.173
R32834 out_p.n1451 out_p.t2875 7.173
R32835 out_p.n1450 out_p.t1154 7.173
R32836 out_p.n1450 out_p.t2410 7.173
R32837 out_p.n1449 out_p.t937 7.173
R32838 out_p.n1449 out_p.t1921 7.173
R32839 out_p.n1492 out_p.t1239 7.173
R32840 out_p.n1492 out_p.t446 7.173
R32841 out_p.n1491 out_p.t759 7.173
R32842 out_p.n1491 out_p.t1597 7.173
R32843 out_p.n1490 out_p.t1009 7.173
R32844 out_p.n1490 out_p.t2071 7.173
R32845 out_p.n1489 out_p.t1390 7.173
R32846 out_p.n1489 out_p.t938 7.173
R32847 out_p.n1488 out_p.t2969 7.173
R32848 out_p.n1488 out_p.t461 7.173
R32849 out_p.n1487 out_p.t2073 7.173
R32850 out_p.n1487 out_p.t2900 7.173
R32851 out_p.n1486 out_p.t941 7.173
R32852 out_p.n1486 out_p.t1925 7.173
R32853 out_p.n1485 out_p.t3374 7.173
R32854 out_p.n1485 out_p.t2517 7.173
R32855 out_p.n1484 out_p.t1327 7.173
R32856 out_p.n1484 out_p.t3174 7.173
R32857 out_p.n1483 out_p.t2042 7.173
R32858 out_p.n1483 out_p.t2818 7.173
R32859 out_p.n1482 out_p.t1969 7.173
R32860 out_p.n1482 out_p.t1079 7.173
R32861 out_p.n1481 out_p.t2930 7.173
R32862 out_p.n1481 out_p.t2384 7.173
R32863 out_p.n1480 out_p.t3396 7.173
R32864 out_p.n1480 out_p.t2494 7.173
R32865 out_p.n1479 out_p.t965 7.173
R32866 out_p.n1479 out_p.t1778 7.173
R32867 out_p.n1478 out_p.t709 7.173
R32868 out_p.n1478 out_p.t3358 7.173
R32869 out_p.n1477 out_p.t2404 7.173
R32870 out_p.n1477 out_p.t2951 7.173
R32871 out_p.n1476 out_p.t1209 7.173
R32872 out_p.n1476 out_p.t507 7.173
R32873 out_p.n1475 out_p.t3224 7.173
R32874 out_p.n1475 out_p.t453 7.173
R32875 out_p.n1474 out_p.t2150 7.173
R32876 out_p.n1474 out_p.t1137 7.173
R32877 out_p.n1473 out_p.t433 7.173
R32878 out_p.n1473 out_p.t907 7.173
R32879 out_p.n1516 out_p.t2835 7.173
R32880 out_p.n1516 out_p.t1261 7.173
R32881 out_p.n1515 out_p.t3260 7.173
R32882 out_p.n1515 out_p.t735 7.173
R32883 out_p.n1514 out_p.t1949 7.173
R32884 out_p.n1514 out_p.t992 7.173
R32885 out_p.n1513 out_p.t2512 7.173
R32886 out_p.n1513 out_p.t432 7.173
R32887 out_p.n1512 out_p.t2189 7.173
R32888 out_p.n1512 out_p.t2957 7.173
R32889 out_p.n1511 out_p.t994 7.173
R32890 out_p.n1511 out_p.t2027 7.173
R32891 out_p.n1510 out_p.t436 7.173
R32892 out_p.n1510 out_p.t914 7.173
R32893 out_p.n1509 out_p.t751 7.173
R32894 out_p.n1509 out_p.t3393 7.173
R32895 out_p.n1508 out_p.t3079 7.173
R32896 out_p.n1508 out_p.t1233 7.173
R32897 out_p.n1507 out_p.t3162 7.173
R32898 out_p.n1507 out_p.t2091 7.173
R32899 out_p.n1506 out_p.t2745 7.173
R32900 out_p.n1506 out_p.t2015 7.173
R32901 out_p.n1505 out_p.t2445 7.173
R32902 out_p.n1505 out_p.t2954 7.173
R32903 out_p.n1504 out_p.t777 7.173
R32904 out_p.n1504 out_p.t3424 7.173
R32905 out_p.n1503 out_p.t1757 7.173
R32906 out_p.n1503 out_p.t990 7.173
R32907 out_p.n1502 out_p.t2373 7.173
R32908 out_p.n1502 out_p.t730 7.173
R32909 out_p.n1501 out_p.t3298 7.173
R32910 out_p.n1501 out_p.t1332 7.173
R32911 out_p.n1500 out_p.t848 7.173
R32912 out_p.n1500 out_p.t1213 7.173
R32913 out_p.n1499 out_p.t603 7.173
R32914 out_p.n1499 out_p.t3249 7.173
R32915 out_p.n1498 out_p.t550 7.173
R32916 out_p.n1498 out_p.t2058 7.173
R32917 out_p.n1497 out_p.t1294 7.173
R32918 out_p.n1497 out_p.t3402 7.173
R32919 out_p.n1540 out_p.t1427 7.173
R32920 out_p.n1540 out_p.t2822 7.173
R32921 out_p.n1539 out_p.t2215 7.173
R32922 out_p.n1539 out_p.t3236 7.173
R32923 out_p.n1538 out_p.t1846 7.173
R32924 out_p.n1538 out_p.t1210 7.173
R32925 out_p.n1537 out_p.t2552 7.173
R32926 out_p.n1537 out_p.t1290 7.173
R32927 out_p.n1536 out_p.t770 7.173
R32928 out_p.n1536 out_p.t2156 7.173
R32929 out_p.n1535 out_p.t3216 7.173
R32930 out_p.n1535 out_p.t975 7.173
R32931 out_p.n1534 out_p.t1547 7.173
R32932 out_p.n1534 out_p.t3408 7.173
R32933 out_p.n1533 out_p.t1433 7.173
R32934 out_p.n1533 out_p.t772 7.173
R32935 out_p.n1532 out_p.t1533 7.173
R32936 out_p.n1532 out_p.t2977 7.173
R32937 out_p.n1531 out_p.t523 7.173
R32938 out_p.n1531 out_p.t3185 7.173
R32939 out_p.n1530 out_p.t1744 7.173
R32940 out_p.n1530 out_p.t2770 7.173
R32941 out_p.n1529 out_p.t3272 7.173
R32942 out_p.n1529 out_p.t1254 7.173
R32943 out_p.n1528 out_p.t1395 7.173
R32944 out_p.n1528 out_p.t806 7.173
R32945 out_p.n1527 out_p.t2612 7.173
R32946 out_p.n1527 out_p.t1794 7.173
R32947 out_p.n1526 out_p.t1052 7.173
R32948 out_p.n1526 out_p.t2503 7.173
R32949 out_p.n1525 out_p.t648 7.173
R32950 out_p.n1525 out_p.t3320 7.173
R32951 out_p.n1524 out_p.t1528 7.173
R32952 out_p.n1524 out_p.t862 7.173
R32953 out_p.n1523 out_p.t1536 7.173
R32954 out_p.n1523 out_p.t630 7.173
R32955 out_p.n1522 out_p.t2784 7.173
R32956 out_p.n1522 out_p.t537 7.173
R32957 out_p.n1521 out_p.t2530 7.173
R32958 out_p.n1521 out_p.t2428 7.173
R32959 out_p.n1564 out_p.t650 7.173
R32960 out_p.n1564 out_p.t3336 7.173
R32961 out_p.n1563 out_p.t1054 7.173
R32962 out_p.n1563 out_p.t1396 7.173
R32963 out_p.n1562 out_p.t2618 7.173
R32964 out_p.n1562 out_p.t1826 7.173
R32965 out_p.n1561 out_p.t1400 7.173
R32966 out_p.n1561 out_p.t822 7.173
R32967 out_p.n1560 out_p.t3275 7.173
R32968 out_p.n1560 out_p.t1258 7.173
R32969 out_p.n1559 out_p.t1764 7.173
R32970 out_p.n1559 out_p.t2788 7.173
R32971 out_p.n1558 out_p.t2535 7.173
R32972 out_p.n1558 out_p.t1699 7.173
R32973 out_p.n1557 out_p.t1083 7.173
R32974 out_p.n1557 out_p.t1216 7.173
R32975 out_p.n1556 out_p.t915 7.173
R32976 out_p.n1556 out_p.t1527 7.173
R32977 out_p.n1555 out_p.t2077 7.173
R32978 out_p.n1555 out_p.t2433 7.173
R32979 out_p.n1554 out_p.t3089 7.173
R32980 out_p.n1554 out_p.t2237 7.173
R32981 out_p.n1553 out_p.t651 7.173
R32982 out_p.n1553 out_p.t3047 7.173
R32983 out_p.n1552 out_p.t1107 7.173
R32984 out_p.n1552 out_p.t1223 7.173
R32985 out_p.n1551 out_p.t2460 7.173
R32986 out_p.n1551 out_p.t1074 7.173
R32987 out_p.n1550 out_p.t1945 7.173
R32988 out_p.n1550 out_p.t845 7.173
R32989 out_p.n1549 out_p.t1988 7.173
R32990 out_p.n1549 out_p.t1256 7.173
R32991 out_p.n1548 out_p.t1167 7.173
R32992 out_p.n1548 out_p.t1752 7.173
R32993 out_p.n1547 out_p.t950 7.173
R32994 out_p.n1547 out_p.t3353 7.173
R32995 out_p.n1546 out_p.t1793 7.173
R32996 out_p.n1546 out_p.t1042 7.173
R32997 out_p.n1545 out_p.t2508 7.173
R32998 out_p.n1545 out_p.t797 7.173
R32999 out_p.n1588 out_p.t3143 7.173
R33000 out_p.n1588 out_p.t969 7.173
R33001 out_p.n1587 out_p.t1416 7.173
R33002 out_p.n1587 out_p.t2685 7.173
R33003 out_p.n1586 out_p.t1495 7.173
R33004 out_p.n1586 out_p.t2937 7.173
R33005 out_p.n1585 out_p.t634 7.173
R33006 out_p.n1585 out_p.t1979 7.173
R33007 out_p.n1584 out_p.t1977 7.173
R33008 out_p.n1584 out_p.t1694 7.173
R33009 out_p.n1583 out_p.t2593 7.173
R33010 out_p.n1583 out_p.t1312 7.173
R33011 out_p.n1582 out_p.t1369 7.173
R33012 out_p.n1582 out_p.t2853 7.173
R33013 out_p.n1581 out_p.t2028 7.173
R33014 out_p.n1581 out_p.t1786 7.173
R33015 out_p.n1580 out_p.t1930 7.173
R33016 out_p.n1580 out_p.t2871 7.173
R33017 out_p.n1579 out_p.t873 7.173
R33018 out_p.n1579 out_p.t1179 7.173
R33019 out_p.n1578 out_p.t470 7.173
R33020 out_p.n1578 out_p.t787 7.173
R33021 out_p.n1577 out_p.t1989 7.173
R33022 out_p.n1577 out_p.t1768 7.173
R33023 out_p.n1576 out_p.t2084 7.173
R33024 out_p.n1576 out_p.t1894 7.173
R33025 out_p.n1575 out_p.t2974 7.173
R33026 out_p.n1575 out_p.t3308 7.173
R33027 out_p.n1574 out_p.t2730 7.173
R33028 out_p.n1574 out_p.t3050 7.173
R33029 out_p.n1573 out_p.t1015 7.173
R33030 out_p.n1573 out_p.t2646 7.173
R33031 out_p.n1572 out_p.t2216 7.173
R33032 out_p.n1572 out_p.t2093 7.173
R33033 out_p.n1571 out_p.t1723 7.173
R33034 out_p.n1571 out_p.t2375 7.173
R33035 out_p.n1570 out_p.t853 7.173
R33036 out_p.n1570 out_p.t2424 7.173
R33037 out_p.n1569 out_p.t609 7.173
R33038 out_p.n1569 out_p.t1932 7.173
R33039 out_p.n1612 out_p.t3318 7.173
R33040 out_p.n1612 out_p.t1497 7.173
R33041 out_p.n1611 out_p.t2509 7.173
R33042 out_p.n1611 out_p.t1611 7.173
R33043 out_p.n1610 out_p.t1792 7.173
R33044 out_p.n1610 out_p.t2108 7.173
R33045 out_p.n1609 out_p.t802 7.173
R33046 out_p.n1609 out_p.t953 7.173
R33047 out_p.n1608 out_p.t1271 7.173
R33048 out_p.n1608 out_p.t477 7.173
R33049 out_p.n1607 out_p.t2768 7.173
R33050 out_p.n1607 out_p.t2917 7.173
R33051 out_p.n1606 out_p.t1653 7.173
R33052 out_p.n1606 out_p.t1946 7.173
R33053 out_p.n1605 out_p.t2269 7.173
R33054 out_p.n1605 out_p.t3094 7.173
R33055 out_p.n1604 out_p.t2361 7.173
R33056 out_p.n1604 out_p.t2396 7.173
R33057 out_p.n1603 out_p.t1326 7.173
R33058 out_p.n1603 out_p.t2251 7.173
R33059 out_p.n1602 out_p.t2279 7.173
R33060 out_p.n1602 out_p.t1464 7.173
R33061 out_p.n1601 out_p.t3072 7.173
R33062 out_p.n1601 out_p.t2651 7.173
R33063 out_p.n1600 out_p.t2345 7.173
R33064 out_p.n1600 out_p.t3125 7.173
R33065 out_p.n1599 out_p.t1093 7.173
R33066 out_p.n1599 out_p.t679 7.173
R33067 out_p.n1598 out_p.t859 7.173
R33068 out_p.n1598 out_p.t2491 7.173
R33069 out_p.n1597 out_p.t1345 7.173
R33070 out_p.n1597 out_p.t1448 7.173
R33071 out_p.n1596 out_p.t1881 7.173
R33072 out_p.n1596 out_p.t3189 7.173
R33073 out_p.n1595 out_p.t3371 7.173
R33074 out_p.n1595 out_p.t2950 7.173
R33075 out_p.n1594 out_p.t1032 7.173
R33076 out_p.n1594 out_p.t1147 7.173
R33077 out_p.n1593 out_p.t775 7.173
R33078 out_p.n1593 out_p.t928 7.173
R33079 out_p.n1636 out_p.t2782 7.173
R33080 out_p.n1636 out_p.t605 7.173
R33081 out_p.n1635 out_p.t3198 7.173
R33082 out_p.n1635 out_p.t1028 7.173
R33083 out_p.n1634 out_p.t443 7.173
R33084 out_p.n1634 out_p.t2568 7.173
R33085 out_p.n1633 out_p.t1238 7.173
R33086 out_p.n1633 out_p.t2391 7.173
R33087 out_p.n1632 out_p.t2059 7.173
R33088 out_p.n1632 out_p.t3230 7.173
R33089 out_p.n1631 out_p.t932 7.173
R33090 out_p.n1631 out_p.t1591 7.173
R33091 out_p.n1630 out_p.t3369 7.173
R33092 out_p.n1630 out_p.t1171 7.173
R33093 out_p.n1629 out_p.t564 7.173
R33094 out_p.n1629 out_p.t877 7.173
R33095 out_p.n1628 out_p.t2127 7.173
R33096 out_p.n1628 out_p.t2921 7.173
R33097 out_p.n1627 out_p.t2970 7.173
R33098 out_p.n1627 out_p.t3299 7.173
R33099 out_p.n1626 out_p.t2547 7.173
R33100 out_p.n1626 out_p.t2874 7.173
R33101 out_p.n1625 out_p.t1813 7.173
R33102 out_p.n1625 out_p.t2495 7.173
R33103 out_p.n1624 out_p.t588 7.173
R33104 out_p.n1624 out_p.t904 7.173
R33105 out_p.n1623 out_p.t1422 7.173
R33106 out_p.n1623 out_p.t2007 7.173
R33107 out_p.n1622 out_p.t2183 7.173
R33108 out_p.n1622 out_p.t1556 7.173
R33109 out_p.n1621 out_p.t3101 7.173
R33110 out_p.n1621 out_p.t3419 7.173
R33111 out_p.n1620 out_p.t662 7.173
R33112 out_p.n1620 out_p.t984 7.173
R33113 out_p.n1619 out_p.t2481 7.173
R33114 out_p.n1619 out_p.t723 7.173
R33115 out_p.n1618 out_p.t501 7.173
R33116 out_p.n1618 out_p.t1720 7.173
R33117 out_p.n1617 out_p.t2281 7.173
R33118 out_p.n1617 out_p.t2271 7.173
R33119 out_p.n1660 out_p.t748 7.173
R33120 out_p.n1660 out_p.t3102 7.173
R33121 out_p.n1659 out_p.t1148 7.173
R33122 out_p.n1659 out_p.t2206 7.173
R33123 out_p.n1658 out_p.t2715 7.173
R33124 out_p.n1658 out_p.t1423 7.173
R33125 out_p.n1657 out_p.t1587 7.173
R33126 out_p.n1657 out_p.t586 7.173
R33127 out_p.n1656 out_p.t3377 7.173
R33128 out_p.n1656 out_p.t1814 7.173
R33129 out_p.n1655 out_p.t2163 7.173
R33130 out_p.n1655 out_p.t2548 7.173
R33131 out_p.n1654 out_p.t2662 7.173
R33132 out_p.n1654 out_p.t2295 7.173
R33133 out_p.n1653 out_p.t2500 7.173
R33134 out_p.n1653 out_p.t1613 7.173
R33135 out_p.n1652 out_p.t2946 7.173
R33136 out_p.n1652 out_p.t1406 7.173
R33137 out_p.n1651 out_p.t2848 7.173
R33138 out_p.n1651 out_p.t673 7.173
R33139 out_p.n1650 out_p.t1120 7.173
R33140 out_p.n1650 out_p.t449 7.173
R33141 out_p.n1649 out_p.t1361 7.173
R33142 out_p.n1649 out_p.t3425 7.173
R33143 out_p.n1648 out_p.t488 7.173
R33144 out_p.n1648 out_p.t1644 7.173
R33145 out_p.n1647 out_p.t2057 7.173
R33146 out_p.n1647 out_p.t2766 7.173
R33147 out_p.n1646 out_p.t3399 7.173
R33148 out_p.n1646 out_p.t1189 7.173
R33149 out_p.n1645 out_p.t2988 7.173
R33150 out_p.n1645 out_p.t798 7.173
R33151 out_p.n1644 out_p.t546 7.173
R33152 out_p.n1644 out_p.t1782 7.173
R33153 out_p.n1643 out_p.t2408 7.173
R33154 out_p.n1643 out_p.t2507 7.173
R33155 out_p.n1642 out_p.t2005 7.173
R33156 out_p.n1642 out_p.t816 7.173
R33157 out_p.n1641 out_p.t1554 7.173
R33158 out_p.n1641 out_p.t565 7.173
R33159 out_p.n1684 out_p.t923 7.173
R33160 out_p.n1684 out_p.t2423 7.173
R33161 out_p.n1683 out_p.t2656 7.173
R33162 out_p.n1683 out_p.t1356 7.173
R33163 out_p.n1682 out_p.t2887 7.173
R33164 out_p.n1682 out_p.t646 7.173
R33165 out_p.n1681 out_p.t1902 7.173
R33166 out_p.n1681 out_p.t3082 7.173
R33167 out_p.n1680 out_p.t1373 7.173
R33168 out_p.n1680 out_p.t2611 7.173
R33169 out_p.n1679 out_p.t1268 7.173
R33170 out_p.n1679 out_p.t1389 7.173
R33171 out_p.n1678 out_p.t2826 7.173
R33172 out_p.n1678 out_p.t570 7.173
R33173 out_p.n1677 out_p.t2253 7.173
R33174 out_p.n1677 out_p.t2553 7.173
R33175 out_p.n1676 out_p.t1499 7.173
R33176 out_p.n1676 out_p.t2711 7.173
R33177 out_p.n1675 out_p.t997 7.173
R33178 out_p.n1675 out_p.t2102 7.173
R33179 out_p.n1674 out_p.t572 7.173
R33180 out_p.n1674 out_p.t3244 7.173
R33181 out_p.n1673 out_p.t1397 7.173
R33182 out_p.n1673 out_p.t804 7.173
R33183 out_p.n1672 out_p.t2304 7.173
R33184 out_p.n1672 out_p.t2581 7.173
R33185 out_p.n1671 out_p.t3085 7.173
R33186 out_p.n1671 out_p.t1950 7.173
R33187 out_p.n1670 out_p.t2837 7.173
R33188 out_p.n1670 out_p.t2275 7.173
R33189 out_p.n1669 out_p.t1101 7.173
R33190 out_p.n1669 out_p.t1486 7.173
R33191 out_p.n1668 out_p.t2425 7.173
R33192 out_p.n1668 out_p.t2663 7.173
R33193 out_p.n1667 out_p.t1933 7.173
R33194 out_p.n1667 out_p.t1086 7.173
R33195 out_p.n1666 out_p.t2362 7.173
R33196 out_p.n1666 out_p.t3314 7.173
R33197 out_p.n1665 out_p.t1863 7.173
R33198 out_p.n1665 out_p.t3064 7.173
R33199 out_p.n1708 out_p.t3416 7.173
R33200 out_p.n1708 out_p.t898 7.173
R33201 out_p.n1707 out_p.t1553 7.173
R33202 out_p.n1707 out_p.t2637 7.173
R33203 out_p.n1706 out_p.t2003 7.173
R33204 out_p.n1706 out_p.t2867 7.173
R33205 out_p.n1705 out_p.t900 7.173
R33206 out_p.n1705 out_p.t1864 7.173
R33207 out_p.n1704 out_p.t2489 7.173
R33208 out_p.n1704 out_p.t2325 7.173
R33209 out_p.n1703 out_p.t2872 7.173
R33210 out_p.n1703 out_p.t1319 7.173
R33211 out_p.n1702 out_p.t1875 7.173
R33212 out_p.n1702 out_p.t2810 7.173
R33213 out_p.n1701 out_p.t2878 7.173
R33214 out_p.n1701 out_p.t2298 7.173
R33215 out_p.n1700 out_p.t664 7.173
R33216 out_p.n1700 out_p.t1521 7.173
R33217 out_p.n1699 out_p.t1807 7.173
R33218 out_p.n1699 out_p.t1017 7.173
R33219 out_p.n1698 out_p.t1500 7.173
R33220 out_p.n1698 out_p.t595 7.173
R33221 out_p.n1697 out_p.t1108 7.173
R33222 out_p.n1697 out_p.t1440 7.173
R33223 out_p.n1696 out_p.t2904 7.173
R33224 out_p.n1696 out_p.t2357 7.173
R33225 out_p.n1695 out_p.t466 7.173
R33226 out_p.n1695 out_p.t3114 7.173
R33227 out_p.n1694 out_p.t2176 7.173
R33228 out_p.n1694 out_p.t2854 7.173
R33229 out_p.n1693 out_p.t2082 7.173
R33230 out_p.n1693 out_p.t1124 7.173
R33231 out_p.n1692 out_p.t2971 7.173
R33232 out_p.n1692 out_p.t1365 7.173
R33233 out_p.n1691 out_p.t2724 7.173
R33234 out_p.n1691 out_p.t1980 7.173
R33235 out_p.n1690 out_p.t1114 7.173
R33236 out_p.n1690 out_p.t2323 7.173
R33237 out_p.n1689 out_p.t880 7.173
R33238 out_p.n1689 out_p.t1816 7.173
R33239 out_p.n1732 out_p.t2438 7.173
R33240 out_p.n1732 out_p.t1382 7.173
R33241 out_p.n1731 out_p.t710 7.173
R33242 out_p.n1731 out_p.t2181 7.173
R33243 out_p.n1730 out_p.t966 7.173
R33244 out_p.n1730 out_p.t1729 7.173
R33245 out_p.n1729 out_p.t3397 7.173
R33246 out_p.n1729 out_p.t2525 7.173
R33247 out_p.n1728 out_p.t2931 7.173
R33248 out_p.n1728 out_p.t744 7.173
R33249 out_p.n1727 out_p.t1970 7.173
R33250 out_p.n1727 out_p.t3196 7.173
R33251 out_p.n1726 out_p.t885 7.173
R33252 out_p.n1726 out_p.t1469 7.173
R33253 out_p.n1725 out_p.t456 7.173
R33254 out_p.n1725 out_p.t576 7.173
R33255 out_p.n1724 out_p.t3362 7.173
R33256 out_p.n1724 out_p.t2620 7.173
R33257 out_p.n1723 out_p.t2670 7.173
R33258 out_p.n1723 out_p.t2986 7.173
R33259 out_p.n1722 out_p.t947 7.173
R33260 out_p.n1722 out_p.t2564 7.173
R33261 out_p.n1721 out_p.t2085 7.173
R33262 out_p.n1721 out_p.t1872 7.173
R33263 out_p.n1720 out_p.t2456 7.173
R33264 out_p.n1720 out_p.t606 7.173
R33265 out_p.n1719 out_p.t1194 7.173
R33266 out_p.n1719 out_p.t1453 7.173
R33267 out_p.n1718 out_p.t3208 7.173
R33268 out_p.n1718 out_p.t1224 7.173
R33269 out_p.n1717 out_p.t2798 7.173
R33270 out_p.n1717 out_p.t3121 7.173
R33271 out_p.n1716 out_p.t1226 7.173
R33272 out_p.n1716 out_p.t674 7.173
R33273 out_p.n1715 out_p.t1791 7.173
R33274 out_p.n1715 out_p.t2453 7.173
R33275 out_p.n1714 out_p.t1927 7.173
R33276 out_p.n1714 out_p.t2758 7.173
R33277 out_p.n1713 out_p.t3380 7.173
R33278 out_p.n1713 out_p.t1181 7.173
R33279 out_p.n1756 out_p.t478 7.173
R33280 out_p.n1756 out_p.t622 7.173
R33281 out_p.n1755 out_p.t878 7.173
R33282 out_p.n1755 out_p.t1036 7.173
R33283 out_p.n1754 out_p.t1115 7.173
R33284 out_p.n1754 out_p.t2582 7.173
R33285 out_p.n1753 out_p.t1582 7.173
R33286 out_p.n1753 out_p.t1436 7.173
R33287 out_p.n1752 out_p.t3096 7.173
R33288 out_p.n1752 out_p.t3245 7.173
R33289 out_p.n1751 out_p.t2324 7.173
R33290 out_p.n1751 out_p.t1661 7.173
R33291 out_p.n1750 out_p.t1056 7.173
R33292 out_p.n1750 out_p.t1186 7.173
R33293 out_p.n1749 out_p.t1853 7.173
R33294 out_p.n1749 out_p.t1538 7.173
R33295 out_p.n1748 out_p.t1827 7.173
R33296 out_p.n1748 out_p.t1885 7.173
R33297 out_p.n1747 out_p.t795 7.173
R33298 out_p.n1747 out_p.t1257 7.173
R33299 out_p.n1746 out_p.t1269 7.173
R33300 out_p.n1746 out_p.t2374 7.173
R33301 out_p.n1745 out_p.t1374 7.173
R33302 out_p.n1745 out_p.t3126 7.173
R33303 out_p.n1744 out_p.t1908 7.173
R33304 out_p.n1744 out_p.t1753 7.173
R33305 out_p.n1743 out_p.t2888 7.173
R33306 out_p.n1743 out_p.t1135 7.173
R33307 out_p.n1742 out_p.t2657 7.173
R33308 out_p.n1742 out_p.t901 7.173
R33309 out_p.n1741 out_p.t924 7.173
R33310 out_p.n1741 out_p.t500 7.173
R33311 out_p.n1740 out_p.t2041 7.173
R33312 out_p.n1740 out_p.t2103 7.173
R33313 out_p.n1739 out_p.t1575 7.173
R33314 out_p.n1739 out_p.t3417 7.173
R33315 out_p.n1738 out_p.t1491 7.173
R33316 out_p.n1738 out_p.t1737 7.173
R33317 out_p.n1737 out_p.t1394 7.173
R33318 out_p.n1737 out_p.t2354 7.173
R33319 out_p.n1780 out_p.t2467 7.173
R33320 out_p.n1780 out_p.t789 7.173
R33321 out_p.n1779 out_p.t2146 7.173
R33322 out_p.n1779 out_p.t1180 7.173
R33323 out_p.n1778 out_p.t1658 7.173
R33324 out_p.n1778 out_p.t2754 7.173
R33325 out_p.n1777 out_p.t1182 7.173
R33326 out_p.n1777 out_p.t1630 7.173
R33327 out_p.n1776 out_p.t719 7.173
R33328 out_p.n1776 out_p.t3412 7.173
R33329 out_p.n1775 out_p.t3171 7.173
R33330 out_p.n1775 out_p.t2260 7.173
R33331 out_p.n1774 out_p.t1402 7.173
R33332 out_p.n1774 out_p.t2688 7.173
R33333 out_p.n1773 out_p.t599 7.173
R33334 out_p.n1773 out_p.t3003 7.173
R33335 out_p.n1772 out_p.t1177 7.173
R33336 out_p.n1772 out_p.t1287 7.173
R33337 out_p.n1771 out_p.t3006 7.173
R33338 out_p.n1771 out_p.t2076 7.173
R33339 out_p.n1770 out_p.t2589 7.173
R33340 out_p.n1770 out_p.t2292 7.173
R33341 out_p.n1769 out_p.t1955 7.173
R33342 out_p.n1769 out_p.t2549 7.173
R33343 out_p.n1768 out_p.t632 7.173
R33344 out_p.n1768 out_p.t3027 7.173
R33345 out_p.n1767 out_p.t1492 7.173
R33346 out_p.n1767 out_p.t587 7.173
R33347 out_p.n1766 out_p.t1415 7.173
R33348 out_p.n1766 out_p.t1230 7.173
R33349 out_p.n1765 out_p.t3141 7.173
R33350 out_p.n1765 out_p.t2334 7.173
R33351 out_p.n1764 out_p.t696 7.173
R33352 out_p.n1764 out_p.t3103 7.173
R33353 out_p.n1763 out_p.t2496 7.173
R33354 out_p.n1763 out_p.t2846 7.173
R33355 out_p.n1762 out_p.t2737 7.173
R33356 out_p.n1762 out_p.t2094 7.173
R33357 out_p.n1761 out_p.t1163 7.173
R33358 out_p.n1761 out_p.t1608 7.173
R33359 out_p.n1804 out_p.t596 7.173
R33360 out_p.n1804 out_p.t3290 7.173
R33361 out_p.n1803 out_p.t1019 7.173
R33362 out_p.n1803 out_p.t2329 7.173
R33363 out_p.n1802 out_p.t2560 7.173
R33364 out_p.n1802 out_p.t1733 7.173
R33365 out_p.n1801 out_p.t2355 7.173
R33366 out_p.n1801 out_p.t765 7.173
R33367 out_p.n1800 out_p.t3222 7.173
R33368 out_p.n1800 out_p.t2435 7.173
R33369 out_p.n1799 out_p.t1568 7.173
R33370 out_p.n1799 out_p.t2739 7.173
R33371 out_p.n1798 out_p.t1168 7.173
R33372 out_p.n1798 out_p.t1616 7.173
R33373 out_p.n1797 out_p.t1716 7.173
R33374 out_p.n1797 out_p.t1245 7.173
R33375 out_p.n1796 out_p.t1674 7.173
R33376 out_p.n1796 out_p.t3033 7.173
R33377 out_p.n1795 out_p.t1235 7.173
R33378 out_p.n1795 out_p.t2794 7.173
R33379 out_p.n1794 out_p.t2412 7.173
R33380 out_p.n1794 out_p.t1063 7.173
R33381 out_p.n1793 out_p.t3146 7.173
R33382 out_p.n1793 out_p.t2336 7.173
R33383 out_p.n1792 out_p.t1882 7.173
R33384 out_p.n1792 out_p.t2478 7.173
R33385 out_p.n1791 out_p.t1152 7.173
R33386 out_p.n1791 out_p.t1625 7.173
R33387 out_p.n1790 out_p.t933 7.173
R33388 out_p.n1790 out_p.t3340 7.173
R33389 out_p.n1789 out_p.t520 7.173
R33390 out_p.n1789 out_p.t2928 7.173
R33391 out_p.n1788 out_p.t2235 7.173
R33392 out_p.n1788 out_p.t486 7.173
R33393 out_p.n1787 out_p.t450 7.173
R33394 out_p.n1787 out_p.t2212 7.173
R33395 out_p.n1786 out_p.t1702 7.173
R33396 out_p.n1786 out_p.t1001 7.173
R33397 out_p.n1785 out_p.t2187 7.173
R33398 out_p.n1785 out_p.t749 7.173
R33399 out_p.n1828 out_p.t1094 7.173
R33400 out_p.n1828 out_p.t916 7.173
R33401 out_p.n1827 out_p.t2831 7.173
R33402 out_p.n1827 out_p.t2649 7.173
R33403 out_p.n1826 out_p.t3073 7.173
R33404 out_p.n1826 out_p.t2881 7.173
R33405 out_p.n1825 out_p.t2285 7.173
R33406 out_p.n1825 out_p.t1897 7.173
R33407 out_p.n1824 out_p.t1378 7.173
R33408 out_p.n1824 out_p.t2256 7.173
R33409 out_p.n1823 out_p.t562 7.173
R33410 out_p.n1823 out_p.t1322 7.173
R33411 out_p.n1822 out_p.t3004 7.173
R33412 out_p.n1822 out_p.t2819 7.173
R33413 out_p.n1821 out_p.t703 7.173
R33414 out_p.n1821 out_p.t2596 7.173
R33415 out_p.n1820 out_p.t985 7.173
R33416 out_p.n1820 out_p.t2282 7.173
R33417 out_p.n1819 out_p.t3117 7.173
R33418 out_p.n1819 out_p.t2327 7.173
R33419 out_p.n1818 out_p.t2695 7.173
R33420 out_p.n1818 out_p.t3289 7.173
R33421 out_p.n1817 out_p.t2284 7.173
R33422 out_p.n1817 out_p.t842 7.173
R33423 out_p.n1816 out_p.t720 7.173
R33424 out_p.n1816 out_p.t2626 7.173
R33425 out_p.n1815 out_p.t1650 7.173
R33426 out_p.n1815 out_p.t2045 7.173
R33427 out_p.n1814 out_p.t2080 7.173
R33428 out_p.n1814 out_p.t2346 7.173
R33429 out_p.n1813 out_p.t3241 7.173
R33430 out_p.n1813 out_p.t1539 7.173
R33431 out_p.n1812 out_p.t799 7.173
R33432 out_p.n1812 out_p.t2689 7.173
R33433 out_p.n1811 out_p.t552 7.173
R33434 out_p.n1811 out_p.t1123 7.173
R33435 out_p.n1810 out_p.t1873 7.173
R33436 out_p.n1810 out_p.t2348 7.173
R33437 out_p.n1809 out_p.t2242 7.173
R33438 out_p.n1809 out_p.t1843 7.173
R33439 out_p.n740 out_p.t357 4.355
R33440 out_p.n740 out_p.t387 4.355
R33441 out_p.n741 out_p.t245 4.355
R33442 out_p.n741 out_p.t31 4.355
R33443 out_p.n742 out_p.t3493 4.355
R33444 out_p.n742 out_p.t3497 4.355
R33445 out_p.n743 out_p.t4 4.355
R33446 out_p.n743 out_p.t89 4.355
R33447 out_p.n716 out_p.t126 4.355
R33448 out_p.n716 out_p.t254 4.355
R33449 out_p.n717 out_p.t11 4.355
R33450 out_p.n717 out_p.t355 4.355
R33451 out_p.n718 out_p.t167 4.355
R33452 out_p.n718 out_p.t58 4.355
R33453 out_p.n719 out_p.t3515 4.355
R33454 out_p.n719 out_p.t282 4.355
R33455 out_p.n692 out_p.t10 4.355
R33456 out_p.n692 out_p.t26 4.355
R33457 out_p.n693 out_p.t3556 4.355
R33458 out_p.n693 out_p.t185 4.355
R33459 out_p.n694 out_p.t159 4.355
R33460 out_p.n694 out_p.t221 4.355
R33461 out_p.n695 out_p.t3529 4.355
R33462 out_p.n695 out_p.t3506 4.355
R33463 out_p.n668 out_p.t19 4.355
R33464 out_p.n668 out_p.t339 4.355
R33465 out_p.n669 out_p.t3463 4.355
R33466 out_p.n669 out_p.t374 4.355
R33467 out_p.n670 out_p.t291 4.355
R33468 out_p.n670 out_p.t14 4.355
R33469 out_p.n671 out_p.t109 4.355
R33470 out_p.n671 out_p.t395 4.355
R33471 out_p.n644 out_p.t77 4.355
R33472 out_p.n644 out_p.t313 4.355
R33473 out_p.n645 out_p.t251 4.355
R33474 out_p.n645 out_p.t46 4.355
R33475 out_p.n646 out_p.t3555 4.355
R33476 out_p.n646 out_p.t3577 4.355
R33477 out_p.n647 out_p.t3456 4.355
R33478 out_p.n647 out_p.t222 4.355
R33479 out_p.n620 out_p.t294 4.355
R33480 out_p.n620 out_p.t3523 4.355
R33481 out_p.n621 out_p.t287 4.355
R33482 out_p.n621 out_p.t246 4.355
R33483 out_p.n622 out_p.t143 4.355
R33484 out_p.n622 out_p.t203 4.355
R33485 out_p.n623 out_p.t3581 4.355
R33486 out_p.n623 out_p.t186 4.355
R33487 out_p.n596 out_p.t52 4.355
R33488 out_p.n596 out_p.t3537 4.355
R33489 out_p.n597 out_p.t3501 4.355
R33490 out_p.n597 out_p.t3589 4.355
R33491 out_p.n598 out_p.t270 4.355
R33492 out_p.n598 out_p.t99 4.355
R33493 out_p.n599 out_p.t3433 4.355
R33494 out_p.n599 out_p.t370 4.355
R33495 out_p.n572 out_p.t3520 4.355
R33496 out_p.n572 out_p.t284 4.355
R33497 out_p.n573 out_p.t191 4.355
R33498 out_p.n573 out_p.t3551 4.355
R33499 out_p.n574 out_p.t342 4.355
R33500 out_p.n574 out_p.t178 4.355
R33501 out_p.n575 out_p.t67 4.355
R33502 out_p.n575 out_p.t135 4.355
R33503 out_p.n548 out_p.t278 4.355
R33504 out_p.n548 out_p.t273 4.355
R33505 out_p.n549 out_p.t328 4.355
R33506 out_p.n549 out_p.t283 4.355
R33507 out_p.n550 out_p.t368 4.355
R33508 out_p.n550 out_p.t3579 4.355
R33509 out_p.n551 out_p.t3484 4.355
R33510 out_p.n551 out_p.t297 4.355
R33511 out_p.n524 out_p.t318 4.355
R33512 out_p.n524 out_p.t3509 4.355
R33513 out_p.n525 out_p.t290 4.355
R33514 out_p.n525 out_p.t362 4.355
R33515 out_p.n526 out_p.t3436 4.355
R33516 out_p.n526 out_p.t3502 4.355
R33517 out_p.n527 out_p.t3568 4.355
R33518 out_p.n527 out_p.t219 4.355
R33519 out_p.n500 out_p.t234 4.355
R33520 out_p.n500 out_p.t3595 4.355
R33521 out_p.n501 out_p.t3488 4.355
R33522 out_p.n501 out_p.t3583 4.355
R33523 out_p.n502 out_p.t277 4.355
R33524 out_p.n502 out_p.t3532 4.355
R33525 out_p.n503 out_p.t340 4.355
R33526 out_p.n503 out_p.t371 4.355
R33527 out_p.n476 out_p.t322 4.355
R33528 out_p.n476 out_p.t3527 4.355
R33529 out_p.n477 out_p.t304 4.355
R33530 out_p.n477 out_p.t56 4.355
R33531 out_p.n478 out_p.t3557 4.355
R33532 out_p.n478 out_p.t248 4.355
R33533 out_p.n479 out_p.t349 4.355
R33534 out_p.n479 out_p.t3437 4.355
R33535 out_p.n452 out_p.t187 4.355
R33536 out_p.n452 out_p.t3486 4.355
R33537 out_p.n453 out_p.t386 4.355
R33538 out_p.n453 out_p.t389 4.355
R33539 out_p.n454 out_p.t133 4.355
R33540 out_p.n454 out_p.t32 4.355
R33541 out_p.n455 out_p.t417 4.355
R33542 out_p.n455 out_p.t412 4.355
R33543 out_p.n428 out_p.t272 4.355
R33544 out_p.n428 out_p.t38 4.355
R33545 out_p.n429 out_p.t259 4.355
R33546 out_p.n429 out_p.t12 4.355
R33547 out_p.n430 out_p.t154 4.355
R33548 out_p.n430 out_p.t3535 4.355
R33549 out_p.n431 out_p.t3507 4.355
R33550 out_p.n431 out_p.t116 4.355
R33551 out_p.n404 out_p.t377 4.355
R33552 out_p.n404 out_p.t286 4.355
R33553 out_p.n405 out_p.t25 4.355
R33554 out_p.n405 out_p.t424 4.355
R33555 out_p.n406 out_p.t3550 4.355
R33556 out_p.n406 out_p.t3461 4.355
R33557 out_p.n407 out_p.t111 4.355
R33558 out_p.n407 out_p.t150 4.355
R33559 out_p.n380 out_p.t43 4.355
R33560 out_p.n380 out_p.t68 4.355
R33561 out_p.n381 out_p.t18 4.355
R33562 out_p.n381 out_p.t80 4.355
R33563 out_p.n382 out_p.t3599 4.355
R33564 out_p.n382 out_p.t247 4.355
R33565 out_p.n383 out_p.t122 4.355
R33566 out_p.n383 out_p.t61 4.355
R33567 out_p.n356 out_p.t3470 4.355
R33568 out_p.n356 out_p.t3511 4.355
R33569 out_p.n357 out_p.t327 4.355
R33570 out_p.n357 out_p.t310 4.355
R33571 out_p.n358 out_p.t217 4.355
R33572 out_p.n358 out_p.t44 4.355
R33573 out_p.n359 out_p.t3539 4.355
R33574 out_p.n359 out_p.t3 4.355
R33575 out_p.n332 out_p.t100 4.355
R33576 out_p.n332 out_p.t3513 4.355
R33577 out_p.n333 out_p.t3505 4.355
R33578 out_p.n333 out_p.t285 4.355
R33579 out_p.n334 out_p.t3571 4.355
R33580 out_p.n334 out_p.t49 4.355
R33581 out_p.n335 out_p.t231 4.355
R33582 out_p.n335 out_p.t3530 4.355
R33583 out_p.n308 out_p.t194 4.355
R33584 out_p.n308 out_p.t88 4.355
R33585 out_p.n309 out_p.t48 4.355
R33586 out_p.n309 out_p.t3566 4.355
R33587 out_p.n310 out_p.t343 4.355
R33588 out_p.n310 out_p.t197 4.355
R33589 out_p.n311 out_p.t237 4.355
R33590 out_p.n311 out_p.t385 4.355
R33591 out_p.n284 out_p.t279 4.355
R33592 out_p.n284 out_p.t363 4.355
R33593 out_p.n285 out_p.t366 4.355
R33594 out_p.n285 out_p.t3469 4.355
R33595 out_p.n286 out_p.t425 4.355
R33596 out_p.n286 out_p.t333 4.355
R33597 out_p.n287 out_p.t220 4.355
R33598 out_p.n287 out_p.t27 4.355
R33599 out_p.n260 out_p.t47 4.355
R33600 out_p.n260 out_p.t53 4.355
R33601 out_p.n261 out_p.t3465 4.355
R33602 out_p.n261 out_p.t317 4.355
R33603 out_p.n262 out_p.t311 4.355
R33604 out_p.n262 out_p.t3526 4.355
R33605 out_p.n263 out_p.t136 4.355
R33606 out_p.n263 out_p.t3573 4.355
R33607 out_p.n236 out_p.t225 4.355
R33608 out_p.n236 out_p.t6 4.355
R33609 out_p.n237 out_p.t3510 4.355
R33610 out_p.n237 out_p.t3435 4.355
R33611 out_p.n238 out_p.t215 4.355
R33612 out_p.n238 out_p.t51 4.355
R33613 out_p.n239 out_p.t3503 4.355
R33614 out_p.n239 out_p.t3591 4.355
R33615 out_p.n212 out_p.t252 4.355
R33616 out_p.n212 out_p.t392 4.355
R33617 out_p.n213 out_p.t189 4.355
R33618 out_p.n213 out_p.t123 4.355
R33619 out_p.n214 out_p.t274 4.355
R33620 out_p.n214 out_p.t98 4.355
R33621 out_p.n215 out_p.t180 4.355
R33622 out_p.n215 out_p.t82 4.355
R33623 out_p.n188 out_p.t132 4.355
R33624 out_p.n188 out_p.t9 4.355
R33625 out_p.n189 out_p.t3490 4.355
R33626 out_p.n189 out_p.t419 4.355
R33627 out_p.n190 out_p.t223 4.355
R33628 out_p.n190 out_p.t296 4.355
R33629 out_p.n191 out_p.t330 4.355
R33630 out_p.n191 out_p.t158 4.355
R33631 out_p.n164 out_p.t148 4.355
R33632 out_p.n164 out_p.t3548 4.355
R33633 out_p.n165 out_p.t3541 4.355
R33634 out_p.n165 out_p.t384 4.355
R33635 out_p.n166 out_p.t300 4.355
R33636 out_p.n166 out_p.t3562 4.355
R33637 out_p.n167 out_p.t3561 4.355
R33638 out_p.n167 out_p.t3517 4.355
R33639 out_p.n140 out_p.t23 4.355
R33640 out_p.n140 out_p.t3597 4.355
R33641 out_p.n141 out_p.t3474 4.355
R33642 out_p.n141 out_p.t3477 4.355
R33643 out_p.n142 out_p.t380 4.355
R33644 out_p.n142 out_p.t3445 4.355
R33645 out_p.n143 out_p.t83 4.355
R33646 out_p.n143 out_p.t308 4.355
R33647 out_p.n116 out_p.t268 4.355
R33648 out_p.n116 out_p.t352 4.355
R33649 out_p.n117 out_p.t3553 4.355
R33650 out_p.n117 out_p.t218 4.355
R33651 out_p.n118 out_p.t72 4.355
R33652 out_p.n118 out_p.t21 4.355
R33653 out_p.n119 out_p.t367 4.355
R33654 out_p.n119 out_p.t170 4.355
R33655 out_p.n92 out_p.t332 4.355
R33656 out_p.n92 out_p.t3500 4.355
R33657 out_p.n93 out_p.t266 4.355
R33658 out_p.n93 out_p.t3496 4.355
R33659 out_p.n94 out_p.t3481 4.355
R33660 out_p.n94 out_p.t3448 4.355
R33661 out_p.n95 out_p.t3543 4.355
R33662 out_p.n95 out_p.t364 4.355
R33663 out_p.n68 out_p.t365 4.355
R33664 out_p.n68 out_p.t3514 4.355
R33665 out_p.n69 out_p.t305 4.355
R33666 out_p.n69 out_p.t102 4.355
R33667 out_p.n70 out_p.t312 4.355
R33668 out_p.n70 out_p.t350 4.355
R33669 out_p.n71 out_p.t3432 4.355
R33670 out_p.n71 out_p.t210 4.355
R33671 out_p.n44 out_p.t176 4.355
R33672 out_p.n44 out_p.t306 4.355
R33673 out_p.n45 out_p.t97 4.355
R33674 out_p.n45 out_p.t118 4.355
R33675 out_p.n46 out_p.t326 4.355
R33676 out_p.n46 out_p.t96 4.355
R33677 out_p.n47 out_p.t65 4.355
R33678 out_p.n47 out_p.t207 4.355
R33679 out_p.n20 out_p.t3590 4.355
R33680 out_p.n20 out_p.t3586 4.355
R33681 out_p.n21 out_p.t3575 4.355
R33682 out_p.n21 out_p.t334 4.355
R33683 out_p.n22 out_p.t3567 4.355
R33684 out_p.n22 out_p.t3462 4.355
R33685 out_p.n23 out_p.t208 4.355
R33686 out_p.n23 out_p.t230 4.355
R33687 out_p.n801 out_p.t3522 4.355
R33688 out_p.n801 out_p.t288 4.355
R33689 out_p.n802 out_p.t50 4.355
R33690 out_p.n802 out_p.t216 4.355
R33691 out_p.n803 out_p.t3466 4.355
R33692 out_p.n803 out_p.t3450 4.355
R33693 out_p.n804 out_p.t378 4.355
R33694 out_p.n804 out_p.t33 4.355
R33695 out_p.n845 out_p.t39 4.355
R33696 out_p.n845 out_p.t3491 4.355
R33697 out_p.n846 out_p.t3504 4.355
R33698 out_p.n846 out_p.t276 4.355
R33699 out_p.n847 out_p.t104 4.355
R33700 out_p.n847 out_p.t319 4.355
R33701 out_p.n848 out_p.t3549 4.355
R33702 out_p.n848 out_p.t40 4.355
R33703 out_p.n869 out_p.t144 4.355
R33704 out_p.n869 out_p.t303 4.355
R33705 out_p.n870 out_p.t3588 4.355
R33706 out_p.n870 out_p.t193 4.355
R33707 out_p.n871 out_p.t127 4.355
R33708 out_p.n871 out_p.t63 4.355
R33709 out_p.n872 out_p.t3457 4.355
R33710 out_p.n872 out_p.t3482 4.355
R33711 out_p.n893 out_p.t164 4.355
R33712 out_p.n893 out_p.t160 4.355
R33713 out_p.n894 out_p.t302 4.355
R33714 out_p.n894 out_p.t3563 4.355
R33715 out_p.n895 out_p.t141 4.355
R33716 out_p.n895 out_p.t3455 4.355
R33717 out_p.n896 out_p.t3569 4.355
R33718 out_p.n896 out_p.t3593 4.355
R33719 out_p.n917 out_p.t3533 4.355
R33720 out_p.n917 out_p.t292 4.355
R33721 out_p.n918 out_p.t295 4.355
R33722 out_p.n918 out_p.t182 4.355
R33723 out_p.n919 out_p.t3430 4.355
R33724 out_p.n919 out_p.t3544 4.355
R33725 out_p.n920 out_p.t3519 4.355
R33726 out_p.n920 out_p.t108 4.355
R33727 out_p.n941 out_p.t24 4.355
R33728 out_p.n941 out_p.t289 4.355
R33729 out_p.n942 out_p.t3554 4.355
R33730 out_p.n942 out_p.t22 4.355
R33731 out_p.n943 out_p.t383 4.355
R33732 out_p.n943 out_p.t3458 4.355
R33733 out_p.n944 out_p.t57 4.355
R33734 out_p.n944 out_p.t129 4.355
R33735 out_p.n965 out_p.t20 4.355
R33736 out_p.n965 out_p.t400 4.355
R33737 out_p.n966 out_p.t257 4.355
R33738 out_p.n966 out_p.t74 4.355
R33739 out_p.n967 out_p.t375 4.355
R33740 out_p.n967 out_p.t244 4.355
R33741 out_p.n968 out_p.t101 4.355
R33742 out_p.n968 out_p.t354 4.355
R33743 out_p.n989 out_p.t423 4.355
R33744 out_p.n989 out_p.t3585 4.355
R33745 out_p.n990 out_p.t177 4.355
R33746 out_p.n990 out_p.t325 4.355
R33747 out_p.n991 out_p.t3438 4.355
R33748 out_p.n991 out_p.t262 4.355
R33749 out_p.n992 out_p.t8 4.355
R33750 out_p.n992 out_p.t229 4.355
R33751 out_p.n1013 out_p.t202 4.355
R33752 out_p.n1013 out_p.t3525 4.355
R33753 out_p.n1014 out_p.t3578 4.355
R33754 out_p.n1014 out_p.t280 4.355
R33755 out_p.n1015 out_p.t406 4.355
R33756 out_p.n1015 out_p.t316 4.355
R33757 out_p.n1016 out_p.t236 4.355
R33758 out_p.n1016 out_p.t34 4.355
R33759 out_p.n1037 out_p.t190 4.355
R33760 out_p.n1037 out_p.t60 4.355
R33761 out_p.n1038 out_p.t3524 4.355
R33762 out_p.n1038 out_p.t329 4.355
R33763 out_p.n1039 out_p.t181 4.355
R33764 out_p.n1039 out_p.t199 4.355
R33765 out_p.n1040 out_p.t242 4.355
R33766 out_p.n1040 out_p.t3538 4.355
R33767 out_p.n1061 out_p.t131 4.355
R33768 out_p.n1061 out_p.t107 4.355
R33769 out_p.n1062 out_p.t169 4.355
R33770 out_p.n1062 out_p.t399 4.355
R33771 out_p.n1063 out_p.t3558 4.355
R33772 out_p.n1063 out_p.t115 4.355
R33773 out_p.n1064 out_p.t394 4.355
R33774 out_p.n1064 out_p.t3473 4.355
R33775 out_p.n1085 out_p.t3453 4.355
R33776 out_p.n1085 out_p.t3584 4.355
R33777 out_p.n1086 out_p.t200 4.355
R33778 out_p.n1086 out_p.t3518 4.355
R33779 out_p.n1087 out_p.t337 4.355
R33780 out_p.n1087 out_p.t275 4.355
R33781 out_p.n1088 out_p.t66 4.355
R33782 out_p.n1088 out_p.t3574 4.355
R33783 out_p.n1109 out_p.t3489 4.355
R33784 out_p.n1109 out_p.t119 4.355
R33785 out_p.n1110 out_p.t3528 4.355
R33786 out_p.n1110 out_p.t91 4.355
R33787 out_p.n1111 out_p.t281 4.355
R33788 out_p.n1111 out_p.t3512 4.355
R33789 out_p.n1112 out_p.t353 4.355
R33790 out_p.n1112 out_p.t255 4.355
R33791 out_p.n1133 out_p.t241 4.355
R33792 out_p.n1133 out_p.t138 4.355
R33793 out_p.n1134 out_p.t3495 4.355
R33794 out_p.n1134 out_p.t137 4.355
R33795 out_p.n1135 out_p.t360 4.355
R33796 out_p.n1135 out_p.t173 4.355
R33797 out_p.n1136 out_p.t348 4.355
R33798 out_p.n1136 out_p.t345 4.355
R33799 out_p.n1157 out_p.t3560 4.355
R33800 out_p.n1157 out_p.t28 4.355
R33801 out_p.n1158 out_p.t103 4.355
R33802 out_p.n1158 out_p.t3487 4.355
R33803 out_p.n1159 out_p.t309 4.355
R33804 out_p.n1159 out_p.t161 4.355
R33805 out_p.n1160 out_p.t264 4.355
R33806 out_p.n1160 out_p.t351 4.355
R33807 out_p.n1181 out_p.t153 4.355
R33808 out_p.n1181 out_p.t3492 4.355
R33809 out_p.n1182 out_p.t3447 4.355
R33810 out_p.n1182 out_p.t3580 4.355
R33811 out_p.n1183 out_p.t125 4.355
R33812 out_p.n1183 out_p.t3428 4.355
R33813 out_p.n1184 out_p.t179 4.355
R33814 out_p.n1184 out_p.t411 4.355
R33815 out_p.n1205 out_p.t175 4.355
R33816 out_p.n1205 out_p.t3476 4.355
R33817 out_p.n1206 out_p.t37 4.355
R33818 out_p.n1206 out_p.t293 4.355
R33819 out_p.n1207 out_p.t7 4.355
R33820 out_p.n1207 out_p.t146 4.355
R33821 out_p.n1208 out_p.t3565 4.355
R33822 out_p.n1208 out_p.t188 4.355
R33823 out_p.n1229 out_p.t3444 4.355
R33824 out_p.n1229 out_p.t369 4.355
R33825 out_p.n1230 out_p.t388 4.355
R33826 out_p.n1230 out_p.t3471 4.355
R33827 out_p.n1231 out_p.t3440 4.355
R33828 out_p.n1231 out_p.t3570 4.355
R33829 out_p.n1232 out_p.t3485 4.355
R33830 out_p.n1232 out_p.t192 4.355
R33831 out_p.n1253 out_p.t267 4.355
R33832 out_p.n1253 out_p.t405 4.355
R33833 out_p.n1254 out_p.t418 4.355
R33834 out_p.n1254 out_p.t204 4.355
R33835 out_p.n1255 out_p.t76 4.355
R33836 out_p.n1255 out_p.t260 4.355
R33837 out_p.n1256 out_p.t3545 4.355
R33838 out_p.n1256 out_p.t212 4.355
R33839 out_p.n1277 out_p.t341 4.355
R33840 out_p.n1277 out_p.t347 4.355
R33841 out_p.n1278 out_p.t3598 4.355
R33842 out_p.n1278 out_p.t94 4.355
R33843 out_p.n1279 out_p.t86 4.355
R33844 out_p.n1279 out_p.t331 4.355
R33845 out_p.n1280 out_p.t379 4.355
R33846 out_p.n1280 out_p.t3441 4.355
R33847 out_p.n1301 out_p.t198 4.355
R33848 out_p.n1301 out_p.t402 4.355
R33849 out_p.n1302 out_p.t3499 4.355
R33850 out_p.n1302 out_p.t196 4.355
R33851 out_p.n1303 out_p.t408 4.355
R33852 out_p.n1303 out_p.t3508 4.355
R33853 out_p.n1304 out_p.t228 4.355
R33854 out_p.n1304 out_p.t70 4.355
R33855 out_p.n1325 out_p.t117 4.355
R33856 out_p.n1325 out_p.t0 4.355
R33857 out_p.n1326 out_p.t45 4.355
R33858 out_p.n1326 out_p.t3480 4.355
R33859 out_p.n1327 out_p.t338 4.355
R33860 out_p.n1327 out_p.t422 4.355
R33861 out_p.n1328 out_p.t235 4.355
R33862 out_p.n1328 out_p.t356 4.355
R33863 out_p.n1349 out_p.t3559 4.355
R33864 out_p.n1349 out_p.t54 4.355
R33865 out_p.n1350 out_p.t183 4.355
R33866 out_p.n1350 out_p.t335 4.355
R33867 out_p.n1351 out_p.t398 4.355
R33868 out_p.n1351 out_p.t3452 4.355
R33869 out_p.n1352 out_p.t263 4.355
R33870 out_p.n1352 out_p.t391 4.355
R33871 out_p.n1373 out_p.t36 4.355
R33872 out_p.n1373 out_p.t55 4.355
R33873 out_p.n1374 out_p.t416 4.355
R33874 out_p.n1374 out_p.t314 4.355
R33875 out_p.n1375 out_p.t201 4.355
R33876 out_p.n1375 out_p.t3521 4.355
R33877 out_p.n1376 out_p.t3531 4.355
R33878 out_p.n1376 out_p.t16 4.355
R33879 out_p.n1397 out_p.t149 4.355
R33880 out_p.n1397 out_p.t172 4.355
R33881 out_p.n1398 out_p.t5 4.355
R33882 out_p.n1398 out_p.t427 4.355
R33883 out_p.n1399 out_p.t3576 4.355
R33884 out_p.n1399 out_p.t42 4.355
R33885 out_p.n1400 out_p.t382 4.355
R33886 out_p.n1400 out_p.t73 4.355
R33887 out_p.n1421 out_p.t299 4.355
R33888 out_p.n1421 out_p.t301 4.355
R33889 out_p.n1422 out_p.t139 4.355
R33890 out_p.n1422 out_p.t151 4.355
R33891 out_p.n1423 out_p.t140 4.355
R33892 out_p.n1423 out_p.t147 4.355
R33893 out_p.n1424 out_p.t87 4.355
R33894 out_p.n1424 out_p.t84 4.355
R33895 out_p.n1445 out_p.t358 4.355
R33896 out_p.n1445 out_p.t3446 4.355
R33897 out_p.n1446 out_p.t3479 4.355
R33898 out_p.n1446 out_p.t29 4.355
R33899 out_p.n1447 out_p.t3472 4.355
R33900 out_p.n1447 out_p.t165 4.355
R33901 out_p.n1448 out_p.t213 4.355
R33902 out_p.n1448 out_p.t3451 4.355
R33903 out_p.n1469 out_p.t3431 4.355
R33904 out_p.n1469 out_p.t209 4.355
R33905 out_p.n1470 out_p.t3546 4.355
R33906 out_p.n1470 out_p.t233 4.355
R33907 out_p.n1471 out_p.t162 4.355
R33908 out_p.n1471 out_p.t3534 4.355
R33909 out_p.n1472 out_p.t258 4.355
R33910 out_p.n1472 out_p.t3468 4.355
R33911 out_p.n1493 out_p.t15 4.355
R33912 out_p.n1493 out_p.t206 4.355
R33913 out_p.n1494 out_p.t3459 4.355
R33914 out_p.n1494 out_p.t253 4.355
R33915 out_p.n1495 out_p.t3478 4.355
R33916 out_p.n1495 out_p.t3547 4.355
R33917 out_p.n1496 out_p.t69 4.355
R33918 out_p.n1496 out_p.t3467 4.355
R33919 out_p.n1517 out_p.t3536 4.355
R33920 out_p.n1517 out_p.t3442 4.355
R33921 out_p.n1518 out_p.t344 4.355
R33922 out_p.n1518 out_p.t250 4.355
R33923 out_p.n1519 out_p.t3439 4.355
R33924 out_p.n1519 out_p.t407 4.355
R33925 out_p.n1520 out_p.t3494 4.355
R33926 out_p.n1520 out_p.t227 4.355
R33927 out_p.n1541 out_p.t320 4.355
R33928 out_p.n1541 out_p.t105 4.355
R33929 out_p.n1542 out_p.t409 4.355
R33930 out_p.n1542 out_p.t324 4.355
R33931 out_p.n1543 out_p.t81 4.355
R33932 out_p.n1543 out_p.t3596 4.355
R33933 out_p.n1544 out_p.t361 4.355
R33934 out_p.n1544 out_p.t243 4.355
R33935 out_p.n1565 out_p.t166 4.355
R33936 out_p.n1565 out_p.t3564 4.355
R33937 out_p.n1566 out_p.t415 4.355
R33938 out_p.n1566 out_p.t3464 4.355
R33939 out_p.n1567 out_p.t95 4.355
R33940 out_p.n1567 out_p.t90 4.355
R33941 out_p.n1568 out_p.t373 4.355
R33942 out_p.n1568 out_p.t376 4.355
R33943 out_p.n1589 out_p.t121 4.355
R33944 out_p.n1589 out_p.t307 4.355
R33945 out_p.n1590 out_p.t401 4.355
R33946 out_p.n1590 out_p.t426 4.355
R33947 out_p.n1591 out_p.t112 4.355
R33948 out_p.n1591 out_p.t93 4.355
R33949 out_p.n1592 out_p.t403 4.355
R33950 out_p.n1592 out_p.t3449 4.355
R33951 out_p.n1613 out_p.t3460 4.355
R33952 out_p.n1613 out_p.t390 4.355
R33953 out_p.n1614 out_p.t3483 4.355
R33954 out_p.n1614 out_p.t3429 4.355
R33955 out_p.n1615 out_p.t271 4.355
R33956 out_p.n1615 out_p.t134 4.355
R33957 out_p.n1616 out_p.t152 4.355
R33958 out_p.n1616 out_p.t3443 4.355
R33959 out_p.n1637 out_p.t404 4.355
R33960 out_p.n1637 out_p.t195 4.355
R33961 out_p.n1638 out_p.t106 4.355
R33962 out_p.n1638 out_p.t171 4.355
R33963 out_p.n1639 out_p.t3552 4.355
R33964 out_p.n1639 out_p.t414 4.355
R33965 out_p.n1640 out_p.t3592 4.355
R33966 out_p.n1640 out_p.t239 4.355
R33967 out_p.n1661 out_p.t3454 4.355
R33968 out_p.n1661 out_p.t78 4.355
R33969 out_p.n1662 out_p.t214 4.355
R33970 out_p.n1662 out_p.t114 4.355
R33971 out_p.n1663 out_p.t298 4.355
R33972 out_p.n1663 out_p.t224 4.355
R33973 out_p.n1664 out_p.t372 4.355
R33974 out_p.n1664 out_p.t265 4.355
R33975 out_p.n1685 out_p.t124 4.355
R33976 out_p.n1685 out_p.t30 4.355
R33977 out_p.n1686 out_p.t396 4.355
R33978 out_p.n1686 out_p.t13 4.355
R33979 out_p.n1687 out_p.t128 4.355
R33980 out_p.n1687 out_p.t393 4.355
R33981 out_p.n1688 out_p.t397 4.355
R33982 out_p.n1688 out_p.t323 4.355
R33983 out_p.n1709 out_p.t1 4.355
R33984 out_p.n1709 out_p.t226 4.355
R33985 out_p.n1710 out_p.t168 4.355
R33986 out_p.n1710 out_p.t184 4.355
R33987 out_p.n1711 out_p.t142 4.355
R33988 out_p.n1711 out_p.t269 4.355
R33989 out_p.n1712 out_p.t174 4.355
R33990 out_p.n1712 out_p.t163 4.355
R33991 out_p.n1733 out_p.t321 4.355
R33992 out_p.n1733 out_p.t35 4.355
R33993 out_p.n1734 out_p.t381 4.355
R33994 out_p.n1734 out_p.t3434 4.355
R33995 out_p.n1735 out_p.t145 4.355
R33996 out_p.n1735 out_p.t156 4.355
R33997 out_p.n1736 out_p.t3498 4.355
R33998 out_p.n1736 out_p.t110 4.355
R33999 out_p.n1757 out_p.t240 4.355
R34000 out_p.n1757 out_p.t41 4.355
R34001 out_p.n1758 out_p.t3540 4.355
R34002 out_p.n1758 out_p.t17 4.355
R34003 out_p.n1759 out_p.t64 4.355
R34004 out_p.n1759 out_p.t421 4.355
R34005 out_p.n1760 out_p.t2 4.355
R34006 out_p.n1760 out_p.t130 4.355
R34007 out_p.n1781 out_p.t346 4.355
R34008 out_p.n1781 out_p.t420 4.355
R34009 out_p.n1782 out_p.t205 4.355
R34010 out_p.n1782 out_p.t75 4.355
R34011 out_p.n1783 out_p.t249 4.355
R34012 out_p.n1783 out_p.t256 4.355
R34013 out_p.n1784 out_p.t59 4.355
R34014 out_p.n1784 out_p.t155 4.355
R34015 out_p.n1805 out_p.t410 4.355
R34016 out_p.n1805 out_p.t413 4.355
R34017 out_p.n1806 out_p.t3594 4.355
R34018 out_p.n1806 out_p.t85 4.355
R34019 out_p.n1807 out_p.t157 4.355
R34020 out_p.n1807 out_p.t261 4.355
R34021 out_p.n1808 out_p.t211 4.355
R34022 out_p.n1808 out_p.t62 4.355
R34023 out_p.n1829 out_p.t92 4.355
R34024 out_p.n1829 out_p.t113 4.355
R34025 out_p.n1830 out_p.t3572 4.355
R34026 out_p.n1830 out_p.t3542 4.355
R34027 out_p.n1831 out_p.t3475 4.355
R34028 out_p.n1831 out_p.t336 4.355
R34029 out_p.n1832 out_p.t232 4.355
R34030 out_p.n1832 out_p.t238 4.355
R34031 out_p.n744 out_p.t359 4.355
R34032 out_p.n744 out_p.t3582 4.355
R34033 out_p.n745 out_p.t315 4.355
R34034 out_p.n745 out_p.t120 4.355
R34035 out_p.n747 out_p.t3516 4.355
R34036 out_p.n747 out_p.t71 4.355
R34037 out_p.n748 out_p.t3587 4.355
R34038 out_p.n748 out_p.t79 4.355
R34039 out_p.n750 out_p.n749 0.151
R34040 out_p.n751 out_p.n750 0.151
R34041 out_p.n752 out_p.n751 0.151
R34042 out_p.n753 out_p.n752 0.151
R34043 out_p.n754 out_p.n753 0.151
R34044 out_p.n755 out_p.n754 0.151
R34045 out_p.n756 out_p.n755 0.151
R34046 out_p.n757 out_p.n756 0.151
R34047 out_p.n758 out_p.n757 0.151
R34048 out_p.n759 out_p.n758 0.151
R34049 out_p.n760 out_p.n759 0.151
R34050 out_p.n761 out_p.n760 0.151
R34051 out_p.n762 out_p.n761 0.151
R34052 out_p.n763 out_p.n762 0.151
R34053 out_p.n764 out_p.n763 0.151
R34054 out_p.n765 out_p.n764 0.151
R34055 out_p.n766 out_p.n765 0.151
R34056 out_p.n767 out_p.n766 0.151
R34057 out_p.n768 out_p.n767 0.151
R34058 out_p.n721 out_p.n720 0.151
R34059 out_p.n722 out_p.n721 0.151
R34060 out_p.n723 out_p.n722 0.151
R34061 out_p.n724 out_p.n723 0.151
R34062 out_p.n725 out_p.n724 0.151
R34063 out_p.n726 out_p.n725 0.151
R34064 out_p.n727 out_p.n726 0.151
R34065 out_p.n728 out_p.n727 0.151
R34066 out_p.n729 out_p.n728 0.151
R34067 out_p.n730 out_p.n729 0.151
R34068 out_p.n731 out_p.n730 0.151
R34069 out_p.n732 out_p.n731 0.151
R34070 out_p.n733 out_p.n732 0.151
R34071 out_p.n734 out_p.n733 0.151
R34072 out_p.n735 out_p.n734 0.151
R34073 out_p.n736 out_p.n735 0.151
R34074 out_p.n737 out_p.n736 0.151
R34075 out_p.n738 out_p.n737 0.151
R34076 out_p.n739 out_p.n738 0.151
R34077 out_p.n697 out_p.n696 0.151
R34078 out_p.n698 out_p.n697 0.151
R34079 out_p.n699 out_p.n698 0.151
R34080 out_p.n700 out_p.n699 0.151
R34081 out_p.n701 out_p.n700 0.151
R34082 out_p.n702 out_p.n701 0.151
R34083 out_p.n703 out_p.n702 0.151
R34084 out_p.n704 out_p.n703 0.151
R34085 out_p.n705 out_p.n704 0.151
R34086 out_p.n706 out_p.n705 0.151
R34087 out_p.n707 out_p.n706 0.151
R34088 out_p.n708 out_p.n707 0.151
R34089 out_p.n709 out_p.n708 0.151
R34090 out_p.n710 out_p.n709 0.151
R34091 out_p.n711 out_p.n710 0.151
R34092 out_p.n712 out_p.n711 0.151
R34093 out_p.n713 out_p.n712 0.151
R34094 out_p.n714 out_p.n713 0.151
R34095 out_p.n715 out_p.n714 0.151
R34096 out_p.n673 out_p.n672 0.151
R34097 out_p.n674 out_p.n673 0.151
R34098 out_p.n675 out_p.n674 0.151
R34099 out_p.n676 out_p.n675 0.151
R34100 out_p.n677 out_p.n676 0.151
R34101 out_p.n678 out_p.n677 0.151
R34102 out_p.n679 out_p.n678 0.151
R34103 out_p.n680 out_p.n679 0.151
R34104 out_p.n681 out_p.n680 0.151
R34105 out_p.n682 out_p.n681 0.151
R34106 out_p.n683 out_p.n682 0.151
R34107 out_p.n684 out_p.n683 0.151
R34108 out_p.n685 out_p.n684 0.151
R34109 out_p.n686 out_p.n685 0.151
R34110 out_p.n687 out_p.n686 0.151
R34111 out_p.n688 out_p.n687 0.151
R34112 out_p.n689 out_p.n688 0.151
R34113 out_p.n690 out_p.n689 0.151
R34114 out_p.n691 out_p.n690 0.151
R34115 out_p.n649 out_p.n648 0.151
R34116 out_p.n650 out_p.n649 0.151
R34117 out_p.n651 out_p.n650 0.151
R34118 out_p.n652 out_p.n651 0.151
R34119 out_p.n653 out_p.n652 0.151
R34120 out_p.n654 out_p.n653 0.151
R34121 out_p.n655 out_p.n654 0.151
R34122 out_p.n656 out_p.n655 0.151
R34123 out_p.n657 out_p.n656 0.151
R34124 out_p.n658 out_p.n657 0.151
R34125 out_p.n659 out_p.n658 0.151
R34126 out_p.n660 out_p.n659 0.151
R34127 out_p.n661 out_p.n660 0.151
R34128 out_p.n662 out_p.n661 0.151
R34129 out_p.n663 out_p.n662 0.151
R34130 out_p.n664 out_p.n663 0.151
R34131 out_p.n665 out_p.n664 0.151
R34132 out_p.n666 out_p.n665 0.151
R34133 out_p.n667 out_p.n666 0.151
R34134 out_p.n625 out_p.n624 0.151
R34135 out_p.n626 out_p.n625 0.151
R34136 out_p.n627 out_p.n626 0.151
R34137 out_p.n628 out_p.n627 0.151
R34138 out_p.n629 out_p.n628 0.151
R34139 out_p.n630 out_p.n629 0.151
R34140 out_p.n631 out_p.n630 0.151
R34141 out_p.n632 out_p.n631 0.151
R34142 out_p.n633 out_p.n632 0.151
R34143 out_p.n634 out_p.n633 0.151
R34144 out_p.n635 out_p.n634 0.151
R34145 out_p.n636 out_p.n635 0.151
R34146 out_p.n637 out_p.n636 0.151
R34147 out_p.n638 out_p.n637 0.151
R34148 out_p.n639 out_p.n638 0.151
R34149 out_p.n640 out_p.n639 0.151
R34150 out_p.n641 out_p.n640 0.151
R34151 out_p.n642 out_p.n641 0.151
R34152 out_p.n643 out_p.n642 0.151
R34153 out_p.n601 out_p.n600 0.151
R34154 out_p.n602 out_p.n601 0.151
R34155 out_p.n603 out_p.n602 0.151
R34156 out_p.n604 out_p.n603 0.151
R34157 out_p.n605 out_p.n604 0.151
R34158 out_p.n606 out_p.n605 0.151
R34159 out_p.n607 out_p.n606 0.151
R34160 out_p.n608 out_p.n607 0.151
R34161 out_p.n609 out_p.n608 0.151
R34162 out_p.n610 out_p.n609 0.151
R34163 out_p.n611 out_p.n610 0.151
R34164 out_p.n612 out_p.n611 0.151
R34165 out_p.n613 out_p.n612 0.151
R34166 out_p.n614 out_p.n613 0.151
R34167 out_p.n615 out_p.n614 0.151
R34168 out_p.n616 out_p.n615 0.151
R34169 out_p.n617 out_p.n616 0.151
R34170 out_p.n618 out_p.n617 0.151
R34171 out_p.n619 out_p.n618 0.151
R34172 out_p.n577 out_p.n576 0.151
R34173 out_p.n578 out_p.n577 0.151
R34174 out_p.n579 out_p.n578 0.151
R34175 out_p.n580 out_p.n579 0.151
R34176 out_p.n581 out_p.n580 0.151
R34177 out_p.n582 out_p.n581 0.151
R34178 out_p.n583 out_p.n582 0.151
R34179 out_p.n584 out_p.n583 0.151
R34180 out_p.n585 out_p.n584 0.151
R34181 out_p.n586 out_p.n585 0.151
R34182 out_p.n587 out_p.n586 0.151
R34183 out_p.n588 out_p.n587 0.151
R34184 out_p.n589 out_p.n588 0.151
R34185 out_p.n590 out_p.n589 0.151
R34186 out_p.n591 out_p.n590 0.151
R34187 out_p.n592 out_p.n591 0.151
R34188 out_p.n593 out_p.n592 0.151
R34189 out_p.n594 out_p.n593 0.151
R34190 out_p.n595 out_p.n594 0.151
R34191 out_p.n553 out_p.n552 0.151
R34192 out_p.n554 out_p.n553 0.151
R34193 out_p.n555 out_p.n554 0.151
R34194 out_p.n556 out_p.n555 0.151
R34195 out_p.n557 out_p.n556 0.151
R34196 out_p.n558 out_p.n557 0.151
R34197 out_p.n559 out_p.n558 0.151
R34198 out_p.n560 out_p.n559 0.151
R34199 out_p.n561 out_p.n560 0.151
R34200 out_p.n562 out_p.n561 0.151
R34201 out_p.n563 out_p.n562 0.151
R34202 out_p.n564 out_p.n563 0.151
R34203 out_p.n565 out_p.n564 0.151
R34204 out_p.n566 out_p.n565 0.151
R34205 out_p.n567 out_p.n566 0.151
R34206 out_p.n568 out_p.n567 0.151
R34207 out_p.n569 out_p.n568 0.151
R34208 out_p.n570 out_p.n569 0.151
R34209 out_p.n571 out_p.n570 0.151
R34210 out_p.n529 out_p.n528 0.151
R34211 out_p.n530 out_p.n529 0.151
R34212 out_p.n531 out_p.n530 0.151
R34213 out_p.n532 out_p.n531 0.151
R34214 out_p.n533 out_p.n532 0.151
R34215 out_p.n534 out_p.n533 0.151
R34216 out_p.n535 out_p.n534 0.151
R34217 out_p.n536 out_p.n535 0.151
R34218 out_p.n537 out_p.n536 0.151
R34219 out_p.n538 out_p.n537 0.151
R34220 out_p.n539 out_p.n538 0.151
R34221 out_p.n540 out_p.n539 0.151
R34222 out_p.n541 out_p.n540 0.151
R34223 out_p.n542 out_p.n541 0.151
R34224 out_p.n543 out_p.n542 0.151
R34225 out_p.n544 out_p.n543 0.151
R34226 out_p.n545 out_p.n544 0.151
R34227 out_p.n546 out_p.n545 0.151
R34228 out_p.n547 out_p.n546 0.151
R34229 out_p.n505 out_p.n504 0.151
R34230 out_p.n506 out_p.n505 0.151
R34231 out_p.n507 out_p.n506 0.151
R34232 out_p.n508 out_p.n507 0.151
R34233 out_p.n509 out_p.n508 0.151
R34234 out_p.n510 out_p.n509 0.151
R34235 out_p.n511 out_p.n510 0.151
R34236 out_p.n512 out_p.n511 0.151
R34237 out_p.n513 out_p.n512 0.151
R34238 out_p.n514 out_p.n513 0.151
R34239 out_p.n515 out_p.n514 0.151
R34240 out_p.n516 out_p.n515 0.151
R34241 out_p.n517 out_p.n516 0.151
R34242 out_p.n518 out_p.n517 0.151
R34243 out_p.n519 out_p.n518 0.151
R34244 out_p.n520 out_p.n519 0.151
R34245 out_p.n521 out_p.n520 0.151
R34246 out_p.n522 out_p.n521 0.151
R34247 out_p.n523 out_p.n522 0.151
R34248 out_p.n481 out_p.n480 0.151
R34249 out_p.n482 out_p.n481 0.151
R34250 out_p.n483 out_p.n482 0.151
R34251 out_p.n484 out_p.n483 0.151
R34252 out_p.n485 out_p.n484 0.151
R34253 out_p.n486 out_p.n485 0.151
R34254 out_p.n487 out_p.n486 0.151
R34255 out_p.n488 out_p.n487 0.151
R34256 out_p.n489 out_p.n488 0.151
R34257 out_p.n490 out_p.n489 0.151
R34258 out_p.n491 out_p.n490 0.151
R34259 out_p.n492 out_p.n491 0.151
R34260 out_p.n493 out_p.n492 0.151
R34261 out_p.n494 out_p.n493 0.151
R34262 out_p.n495 out_p.n494 0.151
R34263 out_p.n496 out_p.n495 0.151
R34264 out_p.n497 out_p.n496 0.151
R34265 out_p.n498 out_p.n497 0.151
R34266 out_p.n499 out_p.n498 0.151
R34267 out_p.n457 out_p.n456 0.151
R34268 out_p.n458 out_p.n457 0.151
R34269 out_p.n459 out_p.n458 0.151
R34270 out_p.n460 out_p.n459 0.151
R34271 out_p.n461 out_p.n460 0.151
R34272 out_p.n462 out_p.n461 0.151
R34273 out_p.n463 out_p.n462 0.151
R34274 out_p.n464 out_p.n463 0.151
R34275 out_p.n465 out_p.n464 0.151
R34276 out_p.n466 out_p.n465 0.151
R34277 out_p.n467 out_p.n466 0.151
R34278 out_p.n468 out_p.n467 0.151
R34279 out_p.n469 out_p.n468 0.151
R34280 out_p.n470 out_p.n469 0.151
R34281 out_p.n471 out_p.n470 0.151
R34282 out_p.n472 out_p.n471 0.151
R34283 out_p.n473 out_p.n472 0.151
R34284 out_p.n474 out_p.n473 0.151
R34285 out_p.n475 out_p.n474 0.151
R34286 out_p.n433 out_p.n432 0.151
R34287 out_p.n434 out_p.n433 0.151
R34288 out_p.n435 out_p.n434 0.151
R34289 out_p.n436 out_p.n435 0.151
R34290 out_p.n437 out_p.n436 0.151
R34291 out_p.n438 out_p.n437 0.151
R34292 out_p.n439 out_p.n438 0.151
R34293 out_p.n440 out_p.n439 0.151
R34294 out_p.n441 out_p.n440 0.151
R34295 out_p.n442 out_p.n441 0.151
R34296 out_p.n443 out_p.n442 0.151
R34297 out_p.n444 out_p.n443 0.151
R34298 out_p.n445 out_p.n444 0.151
R34299 out_p.n446 out_p.n445 0.151
R34300 out_p.n447 out_p.n446 0.151
R34301 out_p.n448 out_p.n447 0.151
R34302 out_p.n449 out_p.n448 0.151
R34303 out_p.n450 out_p.n449 0.151
R34304 out_p.n451 out_p.n450 0.151
R34305 out_p.n409 out_p.n408 0.151
R34306 out_p.n410 out_p.n409 0.151
R34307 out_p.n411 out_p.n410 0.151
R34308 out_p.n412 out_p.n411 0.151
R34309 out_p.n413 out_p.n412 0.151
R34310 out_p.n414 out_p.n413 0.151
R34311 out_p.n415 out_p.n414 0.151
R34312 out_p.n416 out_p.n415 0.151
R34313 out_p.n417 out_p.n416 0.151
R34314 out_p.n418 out_p.n417 0.151
R34315 out_p.n419 out_p.n418 0.151
R34316 out_p.n420 out_p.n419 0.151
R34317 out_p.n421 out_p.n420 0.151
R34318 out_p.n422 out_p.n421 0.151
R34319 out_p.n423 out_p.n422 0.151
R34320 out_p.n424 out_p.n423 0.151
R34321 out_p.n425 out_p.n424 0.151
R34322 out_p.n426 out_p.n425 0.151
R34323 out_p.n427 out_p.n426 0.151
R34324 out_p.n385 out_p.n384 0.151
R34325 out_p.n386 out_p.n385 0.151
R34326 out_p.n387 out_p.n386 0.151
R34327 out_p.n388 out_p.n387 0.151
R34328 out_p.n389 out_p.n388 0.151
R34329 out_p.n390 out_p.n389 0.151
R34330 out_p.n391 out_p.n390 0.151
R34331 out_p.n392 out_p.n391 0.151
R34332 out_p.n393 out_p.n392 0.151
R34333 out_p.n394 out_p.n393 0.151
R34334 out_p.n395 out_p.n394 0.151
R34335 out_p.n396 out_p.n395 0.151
R34336 out_p.n397 out_p.n396 0.151
R34337 out_p.n398 out_p.n397 0.151
R34338 out_p.n399 out_p.n398 0.151
R34339 out_p.n400 out_p.n399 0.151
R34340 out_p.n401 out_p.n400 0.151
R34341 out_p.n402 out_p.n401 0.151
R34342 out_p.n403 out_p.n402 0.151
R34343 out_p.n361 out_p.n360 0.151
R34344 out_p.n362 out_p.n361 0.151
R34345 out_p.n363 out_p.n362 0.151
R34346 out_p.n364 out_p.n363 0.151
R34347 out_p.n365 out_p.n364 0.151
R34348 out_p.n366 out_p.n365 0.151
R34349 out_p.n367 out_p.n366 0.151
R34350 out_p.n368 out_p.n367 0.151
R34351 out_p.n369 out_p.n368 0.151
R34352 out_p.n370 out_p.n369 0.151
R34353 out_p.n371 out_p.n370 0.151
R34354 out_p.n372 out_p.n371 0.151
R34355 out_p.n373 out_p.n372 0.151
R34356 out_p.n374 out_p.n373 0.151
R34357 out_p.n375 out_p.n374 0.151
R34358 out_p.n376 out_p.n375 0.151
R34359 out_p.n377 out_p.n376 0.151
R34360 out_p.n378 out_p.n377 0.151
R34361 out_p.n379 out_p.n378 0.151
R34362 out_p.n337 out_p.n336 0.151
R34363 out_p.n338 out_p.n337 0.151
R34364 out_p.n339 out_p.n338 0.151
R34365 out_p.n340 out_p.n339 0.151
R34366 out_p.n341 out_p.n340 0.151
R34367 out_p.n342 out_p.n341 0.151
R34368 out_p.n343 out_p.n342 0.151
R34369 out_p.n344 out_p.n343 0.151
R34370 out_p.n345 out_p.n344 0.151
R34371 out_p.n346 out_p.n345 0.151
R34372 out_p.n347 out_p.n346 0.151
R34373 out_p.n348 out_p.n347 0.151
R34374 out_p.n349 out_p.n348 0.151
R34375 out_p.n350 out_p.n349 0.151
R34376 out_p.n351 out_p.n350 0.151
R34377 out_p.n352 out_p.n351 0.151
R34378 out_p.n353 out_p.n352 0.151
R34379 out_p.n354 out_p.n353 0.151
R34380 out_p.n355 out_p.n354 0.151
R34381 out_p.n313 out_p.n312 0.151
R34382 out_p.n314 out_p.n313 0.151
R34383 out_p.n315 out_p.n314 0.151
R34384 out_p.n316 out_p.n315 0.151
R34385 out_p.n317 out_p.n316 0.151
R34386 out_p.n318 out_p.n317 0.151
R34387 out_p.n319 out_p.n318 0.151
R34388 out_p.n320 out_p.n319 0.151
R34389 out_p.n321 out_p.n320 0.151
R34390 out_p.n322 out_p.n321 0.151
R34391 out_p.n323 out_p.n322 0.151
R34392 out_p.n324 out_p.n323 0.151
R34393 out_p.n325 out_p.n324 0.151
R34394 out_p.n326 out_p.n325 0.151
R34395 out_p.n327 out_p.n326 0.151
R34396 out_p.n328 out_p.n327 0.151
R34397 out_p.n329 out_p.n328 0.151
R34398 out_p.n330 out_p.n329 0.151
R34399 out_p.n331 out_p.n330 0.151
R34400 out_p.n289 out_p.n288 0.151
R34401 out_p.n290 out_p.n289 0.151
R34402 out_p.n291 out_p.n290 0.151
R34403 out_p.n292 out_p.n291 0.151
R34404 out_p.n293 out_p.n292 0.151
R34405 out_p.n294 out_p.n293 0.151
R34406 out_p.n295 out_p.n294 0.151
R34407 out_p.n296 out_p.n295 0.151
R34408 out_p.n297 out_p.n296 0.151
R34409 out_p.n298 out_p.n297 0.151
R34410 out_p.n299 out_p.n298 0.151
R34411 out_p.n300 out_p.n299 0.151
R34412 out_p.n301 out_p.n300 0.151
R34413 out_p.n302 out_p.n301 0.151
R34414 out_p.n303 out_p.n302 0.151
R34415 out_p.n304 out_p.n303 0.151
R34416 out_p.n305 out_p.n304 0.151
R34417 out_p.n306 out_p.n305 0.151
R34418 out_p.n307 out_p.n306 0.151
R34419 out_p.n265 out_p.n264 0.151
R34420 out_p.n266 out_p.n265 0.151
R34421 out_p.n267 out_p.n266 0.151
R34422 out_p.n268 out_p.n267 0.151
R34423 out_p.n269 out_p.n268 0.151
R34424 out_p.n270 out_p.n269 0.151
R34425 out_p.n271 out_p.n270 0.151
R34426 out_p.n272 out_p.n271 0.151
R34427 out_p.n273 out_p.n272 0.151
R34428 out_p.n274 out_p.n273 0.151
R34429 out_p.n275 out_p.n274 0.151
R34430 out_p.n276 out_p.n275 0.151
R34431 out_p.n277 out_p.n276 0.151
R34432 out_p.n278 out_p.n277 0.151
R34433 out_p.n279 out_p.n278 0.151
R34434 out_p.n280 out_p.n279 0.151
R34435 out_p.n281 out_p.n280 0.151
R34436 out_p.n282 out_p.n281 0.151
R34437 out_p.n283 out_p.n282 0.151
R34438 out_p.n241 out_p.n240 0.151
R34439 out_p.n242 out_p.n241 0.151
R34440 out_p.n243 out_p.n242 0.151
R34441 out_p.n244 out_p.n243 0.151
R34442 out_p.n245 out_p.n244 0.151
R34443 out_p.n246 out_p.n245 0.151
R34444 out_p.n247 out_p.n246 0.151
R34445 out_p.n248 out_p.n247 0.151
R34446 out_p.n249 out_p.n248 0.151
R34447 out_p.n250 out_p.n249 0.151
R34448 out_p.n251 out_p.n250 0.151
R34449 out_p.n252 out_p.n251 0.151
R34450 out_p.n253 out_p.n252 0.151
R34451 out_p.n254 out_p.n253 0.151
R34452 out_p.n255 out_p.n254 0.151
R34453 out_p.n256 out_p.n255 0.151
R34454 out_p.n257 out_p.n256 0.151
R34455 out_p.n258 out_p.n257 0.151
R34456 out_p.n259 out_p.n258 0.151
R34457 out_p.n217 out_p.n216 0.151
R34458 out_p.n218 out_p.n217 0.151
R34459 out_p.n219 out_p.n218 0.151
R34460 out_p.n220 out_p.n219 0.151
R34461 out_p.n221 out_p.n220 0.151
R34462 out_p.n222 out_p.n221 0.151
R34463 out_p.n223 out_p.n222 0.151
R34464 out_p.n224 out_p.n223 0.151
R34465 out_p.n225 out_p.n224 0.151
R34466 out_p.n226 out_p.n225 0.151
R34467 out_p.n227 out_p.n226 0.151
R34468 out_p.n228 out_p.n227 0.151
R34469 out_p.n229 out_p.n228 0.151
R34470 out_p.n230 out_p.n229 0.151
R34471 out_p.n231 out_p.n230 0.151
R34472 out_p.n232 out_p.n231 0.151
R34473 out_p.n233 out_p.n232 0.151
R34474 out_p.n234 out_p.n233 0.151
R34475 out_p.n235 out_p.n234 0.151
R34476 out_p.n193 out_p.n192 0.151
R34477 out_p.n194 out_p.n193 0.151
R34478 out_p.n195 out_p.n194 0.151
R34479 out_p.n196 out_p.n195 0.151
R34480 out_p.n197 out_p.n196 0.151
R34481 out_p.n198 out_p.n197 0.151
R34482 out_p.n199 out_p.n198 0.151
R34483 out_p.n200 out_p.n199 0.151
R34484 out_p.n201 out_p.n200 0.151
R34485 out_p.n202 out_p.n201 0.151
R34486 out_p.n203 out_p.n202 0.151
R34487 out_p.n204 out_p.n203 0.151
R34488 out_p.n205 out_p.n204 0.151
R34489 out_p.n206 out_p.n205 0.151
R34490 out_p.n207 out_p.n206 0.151
R34491 out_p.n208 out_p.n207 0.151
R34492 out_p.n209 out_p.n208 0.151
R34493 out_p.n210 out_p.n209 0.151
R34494 out_p.n211 out_p.n210 0.151
R34495 out_p.n169 out_p.n168 0.151
R34496 out_p.n170 out_p.n169 0.151
R34497 out_p.n171 out_p.n170 0.151
R34498 out_p.n172 out_p.n171 0.151
R34499 out_p.n173 out_p.n172 0.151
R34500 out_p.n174 out_p.n173 0.151
R34501 out_p.n175 out_p.n174 0.151
R34502 out_p.n176 out_p.n175 0.151
R34503 out_p.n177 out_p.n176 0.151
R34504 out_p.n178 out_p.n177 0.151
R34505 out_p.n179 out_p.n178 0.151
R34506 out_p.n180 out_p.n179 0.151
R34507 out_p.n181 out_p.n180 0.151
R34508 out_p.n182 out_p.n181 0.151
R34509 out_p.n183 out_p.n182 0.151
R34510 out_p.n184 out_p.n183 0.151
R34511 out_p.n185 out_p.n184 0.151
R34512 out_p.n186 out_p.n185 0.151
R34513 out_p.n187 out_p.n186 0.151
R34514 out_p.n145 out_p.n144 0.151
R34515 out_p.n146 out_p.n145 0.151
R34516 out_p.n147 out_p.n146 0.151
R34517 out_p.n148 out_p.n147 0.151
R34518 out_p.n149 out_p.n148 0.151
R34519 out_p.n150 out_p.n149 0.151
R34520 out_p.n151 out_p.n150 0.151
R34521 out_p.n152 out_p.n151 0.151
R34522 out_p.n153 out_p.n152 0.151
R34523 out_p.n154 out_p.n153 0.151
R34524 out_p.n155 out_p.n154 0.151
R34525 out_p.n156 out_p.n155 0.151
R34526 out_p.n157 out_p.n156 0.151
R34527 out_p.n158 out_p.n157 0.151
R34528 out_p.n159 out_p.n158 0.151
R34529 out_p.n160 out_p.n159 0.151
R34530 out_p.n161 out_p.n160 0.151
R34531 out_p.n162 out_p.n161 0.151
R34532 out_p.n163 out_p.n162 0.151
R34533 out_p.n121 out_p.n120 0.151
R34534 out_p.n122 out_p.n121 0.151
R34535 out_p.n123 out_p.n122 0.151
R34536 out_p.n124 out_p.n123 0.151
R34537 out_p.n125 out_p.n124 0.151
R34538 out_p.n126 out_p.n125 0.151
R34539 out_p.n127 out_p.n126 0.151
R34540 out_p.n128 out_p.n127 0.151
R34541 out_p.n129 out_p.n128 0.151
R34542 out_p.n130 out_p.n129 0.151
R34543 out_p.n131 out_p.n130 0.151
R34544 out_p.n132 out_p.n131 0.151
R34545 out_p.n133 out_p.n132 0.151
R34546 out_p.n134 out_p.n133 0.151
R34547 out_p.n135 out_p.n134 0.151
R34548 out_p.n136 out_p.n135 0.151
R34549 out_p.n137 out_p.n136 0.151
R34550 out_p.n138 out_p.n137 0.151
R34551 out_p.n139 out_p.n138 0.151
R34552 out_p.n97 out_p.n96 0.151
R34553 out_p.n98 out_p.n97 0.151
R34554 out_p.n99 out_p.n98 0.151
R34555 out_p.n100 out_p.n99 0.151
R34556 out_p.n101 out_p.n100 0.151
R34557 out_p.n102 out_p.n101 0.151
R34558 out_p.n103 out_p.n102 0.151
R34559 out_p.n104 out_p.n103 0.151
R34560 out_p.n105 out_p.n104 0.151
R34561 out_p.n106 out_p.n105 0.151
R34562 out_p.n107 out_p.n106 0.151
R34563 out_p.n108 out_p.n107 0.151
R34564 out_p.n109 out_p.n108 0.151
R34565 out_p.n110 out_p.n109 0.151
R34566 out_p.n111 out_p.n110 0.151
R34567 out_p.n112 out_p.n111 0.151
R34568 out_p.n113 out_p.n112 0.151
R34569 out_p.n114 out_p.n113 0.151
R34570 out_p.n115 out_p.n114 0.151
R34571 out_p.n73 out_p.n72 0.151
R34572 out_p.n74 out_p.n73 0.151
R34573 out_p.n75 out_p.n74 0.151
R34574 out_p.n76 out_p.n75 0.151
R34575 out_p.n77 out_p.n76 0.151
R34576 out_p.n78 out_p.n77 0.151
R34577 out_p.n79 out_p.n78 0.151
R34578 out_p.n80 out_p.n79 0.151
R34579 out_p.n81 out_p.n80 0.151
R34580 out_p.n82 out_p.n81 0.151
R34581 out_p.n83 out_p.n82 0.151
R34582 out_p.n84 out_p.n83 0.151
R34583 out_p.n85 out_p.n84 0.151
R34584 out_p.n86 out_p.n85 0.151
R34585 out_p.n87 out_p.n86 0.151
R34586 out_p.n88 out_p.n87 0.151
R34587 out_p.n89 out_p.n88 0.151
R34588 out_p.n90 out_p.n89 0.151
R34589 out_p.n91 out_p.n90 0.151
R34590 out_p.n49 out_p.n48 0.151
R34591 out_p.n50 out_p.n49 0.151
R34592 out_p.n51 out_p.n50 0.151
R34593 out_p.n52 out_p.n51 0.151
R34594 out_p.n53 out_p.n52 0.151
R34595 out_p.n54 out_p.n53 0.151
R34596 out_p.n55 out_p.n54 0.151
R34597 out_p.n56 out_p.n55 0.151
R34598 out_p.n57 out_p.n56 0.151
R34599 out_p.n58 out_p.n57 0.151
R34600 out_p.n59 out_p.n58 0.151
R34601 out_p.n60 out_p.n59 0.151
R34602 out_p.n61 out_p.n60 0.151
R34603 out_p.n62 out_p.n61 0.151
R34604 out_p.n63 out_p.n62 0.151
R34605 out_p.n64 out_p.n63 0.151
R34606 out_p.n65 out_p.n64 0.151
R34607 out_p.n66 out_p.n65 0.151
R34608 out_p.n67 out_p.n66 0.151
R34609 out_p.n25 out_p.n24 0.151
R34610 out_p.n26 out_p.n25 0.151
R34611 out_p.n27 out_p.n26 0.151
R34612 out_p.n28 out_p.n27 0.151
R34613 out_p.n29 out_p.n28 0.151
R34614 out_p.n30 out_p.n29 0.151
R34615 out_p.n31 out_p.n30 0.151
R34616 out_p.n32 out_p.n31 0.151
R34617 out_p.n33 out_p.n32 0.151
R34618 out_p.n34 out_p.n33 0.151
R34619 out_p.n35 out_p.n34 0.151
R34620 out_p.n36 out_p.n35 0.151
R34621 out_p.n37 out_p.n36 0.151
R34622 out_p.n38 out_p.n37 0.151
R34623 out_p.n39 out_p.n38 0.151
R34624 out_p.n40 out_p.n39 0.151
R34625 out_p.n41 out_p.n40 0.151
R34626 out_p.n42 out_p.n41 0.151
R34627 out_p.n43 out_p.n42 0.151
R34628 out_p.n1 out_p.n0 0.151
R34629 out_p.n2 out_p.n1 0.151
R34630 out_p.n3 out_p.n2 0.151
R34631 out_p.n4 out_p.n3 0.151
R34632 out_p.n5 out_p.n4 0.151
R34633 out_p.n6 out_p.n5 0.151
R34634 out_p.n7 out_p.n6 0.151
R34635 out_p.n8 out_p.n7 0.151
R34636 out_p.n9 out_p.n8 0.151
R34637 out_p.n10 out_p.n9 0.151
R34638 out_p.n11 out_p.n10 0.151
R34639 out_p.n12 out_p.n11 0.151
R34640 out_p.n13 out_p.n12 0.151
R34641 out_p.n14 out_p.n13 0.151
R34642 out_p.n15 out_p.n14 0.151
R34643 out_p.n16 out_p.n15 0.151
R34644 out_p.n17 out_p.n16 0.151
R34645 out_p.n18 out_p.n17 0.151
R34646 out_p.n19 out_p.n18 0.151
R34647 out_p.n806 out_p.n805 0.151
R34648 out_p.n807 out_p.n806 0.151
R34649 out_p.n808 out_p.n807 0.151
R34650 out_p.n809 out_p.n808 0.151
R34651 out_p.n810 out_p.n809 0.151
R34652 out_p.n811 out_p.n810 0.151
R34653 out_p.n812 out_p.n811 0.151
R34654 out_p.n813 out_p.n812 0.151
R34655 out_p.n814 out_p.n813 0.151
R34656 out_p.n815 out_p.n814 0.151
R34657 out_p.n816 out_p.n815 0.151
R34658 out_p.n817 out_p.n816 0.151
R34659 out_p.n818 out_p.n817 0.151
R34660 out_p.n819 out_p.n818 0.151
R34661 out_p.n820 out_p.n819 0.151
R34662 out_p.n821 out_p.n820 0.151
R34663 out_p.n822 out_p.n821 0.151
R34664 out_p.n823 out_p.n822 0.151
R34665 out_p.n824 out_p.n823 0.151
R34666 out_p.n826 out_p.n825 0.151
R34667 out_p.n827 out_p.n826 0.151
R34668 out_p.n828 out_p.n827 0.151
R34669 out_p.n829 out_p.n828 0.151
R34670 out_p.n830 out_p.n829 0.151
R34671 out_p.n831 out_p.n830 0.151
R34672 out_p.n832 out_p.n831 0.151
R34673 out_p.n833 out_p.n832 0.151
R34674 out_p.n834 out_p.n833 0.151
R34675 out_p.n835 out_p.n834 0.151
R34676 out_p.n836 out_p.n835 0.151
R34677 out_p.n837 out_p.n836 0.151
R34678 out_p.n838 out_p.n837 0.151
R34679 out_p.n839 out_p.n838 0.151
R34680 out_p.n840 out_p.n839 0.151
R34681 out_p.n841 out_p.n840 0.151
R34682 out_p.n842 out_p.n841 0.151
R34683 out_p.n843 out_p.n842 0.151
R34684 out_p.n844 out_p.n843 0.151
R34685 out_p.n850 out_p.n849 0.151
R34686 out_p.n851 out_p.n850 0.151
R34687 out_p.n852 out_p.n851 0.151
R34688 out_p.n853 out_p.n852 0.151
R34689 out_p.n854 out_p.n853 0.151
R34690 out_p.n855 out_p.n854 0.151
R34691 out_p.n856 out_p.n855 0.151
R34692 out_p.n857 out_p.n856 0.151
R34693 out_p.n858 out_p.n857 0.151
R34694 out_p.n859 out_p.n858 0.151
R34695 out_p.n860 out_p.n859 0.151
R34696 out_p.n861 out_p.n860 0.151
R34697 out_p.n862 out_p.n861 0.151
R34698 out_p.n863 out_p.n862 0.151
R34699 out_p.n864 out_p.n863 0.151
R34700 out_p.n865 out_p.n864 0.151
R34701 out_p.n866 out_p.n865 0.151
R34702 out_p.n867 out_p.n866 0.151
R34703 out_p.n868 out_p.n867 0.151
R34704 out_p.n874 out_p.n873 0.151
R34705 out_p.n875 out_p.n874 0.151
R34706 out_p.n876 out_p.n875 0.151
R34707 out_p.n877 out_p.n876 0.151
R34708 out_p.n878 out_p.n877 0.151
R34709 out_p.n879 out_p.n878 0.151
R34710 out_p.n880 out_p.n879 0.151
R34711 out_p.n881 out_p.n880 0.151
R34712 out_p.n882 out_p.n881 0.151
R34713 out_p.n883 out_p.n882 0.151
R34714 out_p.n884 out_p.n883 0.151
R34715 out_p.n885 out_p.n884 0.151
R34716 out_p.n886 out_p.n885 0.151
R34717 out_p.n887 out_p.n886 0.151
R34718 out_p.n888 out_p.n887 0.151
R34719 out_p.n889 out_p.n888 0.151
R34720 out_p.n890 out_p.n889 0.151
R34721 out_p.n891 out_p.n890 0.151
R34722 out_p.n892 out_p.n891 0.151
R34723 out_p.n898 out_p.n897 0.151
R34724 out_p.n899 out_p.n898 0.151
R34725 out_p.n900 out_p.n899 0.151
R34726 out_p.n901 out_p.n900 0.151
R34727 out_p.n902 out_p.n901 0.151
R34728 out_p.n903 out_p.n902 0.151
R34729 out_p.n904 out_p.n903 0.151
R34730 out_p.n905 out_p.n904 0.151
R34731 out_p.n906 out_p.n905 0.151
R34732 out_p.n907 out_p.n906 0.151
R34733 out_p.n908 out_p.n907 0.151
R34734 out_p.n909 out_p.n908 0.151
R34735 out_p.n910 out_p.n909 0.151
R34736 out_p.n911 out_p.n910 0.151
R34737 out_p.n912 out_p.n911 0.151
R34738 out_p.n913 out_p.n912 0.151
R34739 out_p.n914 out_p.n913 0.151
R34740 out_p.n915 out_p.n914 0.151
R34741 out_p.n916 out_p.n915 0.151
R34742 out_p.n922 out_p.n921 0.151
R34743 out_p.n923 out_p.n922 0.151
R34744 out_p.n924 out_p.n923 0.151
R34745 out_p.n925 out_p.n924 0.151
R34746 out_p.n926 out_p.n925 0.151
R34747 out_p.n927 out_p.n926 0.151
R34748 out_p.n928 out_p.n927 0.151
R34749 out_p.n929 out_p.n928 0.151
R34750 out_p.n930 out_p.n929 0.151
R34751 out_p.n931 out_p.n930 0.151
R34752 out_p.n932 out_p.n931 0.151
R34753 out_p.n933 out_p.n932 0.151
R34754 out_p.n934 out_p.n933 0.151
R34755 out_p.n935 out_p.n934 0.151
R34756 out_p.n936 out_p.n935 0.151
R34757 out_p.n937 out_p.n936 0.151
R34758 out_p.n938 out_p.n937 0.151
R34759 out_p.n939 out_p.n938 0.151
R34760 out_p.n940 out_p.n939 0.151
R34761 out_p.n946 out_p.n945 0.151
R34762 out_p.n947 out_p.n946 0.151
R34763 out_p.n948 out_p.n947 0.151
R34764 out_p.n949 out_p.n948 0.151
R34765 out_p.n950 out_p.n949 0.151
R34766 out_p.n951 out_p.n950 0.151
R34767 out_p.n952 out_p.n951 0.151
R34768 out_p.n953 out_p.n952 0.151
R34769 out_p.n954 out_p.n953 0.151
R34770 out_p.n955 out_p.n954 0.151
R34771 out_p.n956 out_p.n955 0.151
R34772 out_p.n957 out_p.n956 0.151
R34773 out_p.n958 out_p.n957 0.151
R34774 out_p.n959 out_p.n958 0.151
R34775 out_p.n960 out_p.n959 0.151
R34776 out_p.n961 out_p.n960 0.151
R34777 out_p.n962 out_p.n961 0.151
R34778 out_p.n963 out_p.n962 0.151
R34779 out_p.n964 out_p.n963 0.151
R34780 out_p.n970 out_p.n969 0.151
R34781 out_p.n971 out_p.n970 0.151
R34782 out_p.n972 out_p.n971 0.151
R34783 out_p.n973 out_p.n972 0.151
R34784 out_p.n974 out_p.n973 0.151
R34785 out_p.n975 out_p.n974 0.151
R34786 out_p.n976 out_p.n975 0.151
R34787 out_p.n977 out_p.n976 0.151
R34788 out_p.n978 out_p.n977 0.151
R34789 out_p.n979 out_p.n978 0.151
R34790 out_p.n980 out_p.n979 0.151
R34791 out_p.n981 out_p.n980 0.151
R34792 out_p.n982 out_p.n981 0.151
R34793 out_p.n983 out_p.n982 0.151
R34794 out_p.n984 out_p.n983 0.151
R34795 out_p.n985 out_p.n984 0.151
R34796 out_p.n986 out_p.n985 0.151
R34797 out_p.n987 out_p.n986 0.151
R34798 out_p.n988 out_p.n987 0.151
R34799 out_p.n994 out_p.n993 0.151
R34800 out_p.n995 out_p.n994 0.151
R34801 out_p.n996 out_p.n995 0.151
R34802 out_p.n997 out_p.n996 0.151
R34803 out_p.n998 out_p.n997 0.151
R34804 out_p.n999 out_p.n998 0.151
R34805 out_p.n1000 out_p.n999 0.151
R34806 out_p.n1001 out_p.n1000 0.151
R34807 out_p.n1002 out_p.n1001 0.151
R34808 out_p.n1003 out_p.n1002 0.151
R34809 out_p.n1004 out_p.n1003 0.151
R34810 out_p.n1005 out_p.n1004 0.151
R34811 out_p.n1006 out_p.n1005 0.151
R34812 out_p.n1007 out_p.n1006 0.151
R34813 out_p.n1008 out_p.n1007 0.151
R34814 out_p.n1009 out_p.n1008 0.151
R34815 out_p.n1010 out_p.n1009 0.151
R34816 out_p.n1011 out_p.n1010 0.151
R34817 out_p.n1012 out_p.n1011 0.151
R34818 out_p.n1018 out_p.n1017 0.151
R34819 out_p.n1019 out_p.n1018 0.151
R34820 out_p.n1020 out_p.n1019 0.151
R34821 out_p.n1021 out_p.n1020 0.151
R34822 out_p.n1022 out_p.n1021 0.151
R34823 out_p.n1023 out_p.n1022 0.151
R34824 out_p.n1024 out_p.n1023 0.151
R34825 out_p.n1025 out_p.n1024 0.151
R34826 out_p.n1026 out_p.n1025 0.151
R34827 out_p.n1027 out_p.n1026 0.151
R34828 out_p.n1028 out_p.n1027 0.151
R34829 out_p.n1029 out_p.n1028 0.151
R34830 out_p.n1030 out_p.n1029 0.151
R34831 out_p.n1031 out_p.n1030 0.151
R34832 out_p.n1032 out_p.n1031 0.151
R34833 out_p.n1033 out_p.n1032 0.151
R34834 out_p.n1034 out_p.n1033 0.151
R34835 out_p.n1035 out_p.n1034 0.151
R34836 out_p.n1036 out_p.n1035 0.151
R34837 out_p.n1042 out_p.n1041 0.151
R34838 out_p.n1043 out_p.n1042 0.151
R34839 out_p.n1044 out_p.n1043 0.151
R34840 out_p.n1045 out_p.n1044 0.151
R34841 out_p.n1046 out_p.n1045 0.151
R34842 out_p.n1047 out_p.n1046 0.151
R34843 out_p.n1048 out_p.n1047 0.151
R34844 out_p.n1049 out_p.n1048 0.151
R34845 out_p.n1050 out_p.n1049 0.151
R34846 out_p.n1051 out_p.n1050 0.151
R34847 out_p.n1052 out_p.n1051 0.151
R34848 out_p.n1053 out_p.n1052 0.151
R34849 out_p.n1054 out_p.n1053 0.151
R34850 out_p.n1055 out_p.n1054 0.151
R34851 out_p.n1056 out_p.n1055 0.151
R34852 out_p.n1057 out_p.n1056 0.151
R34853 out_p.n1058 out_p.n1057 0.151
R34854 out_p.n1059 out_p.n1058 0.151
R34855 out_p.n1060 out_p.n1059 0.151
R34856 out_p.n1066 out_p.n1065 0.151
R34857 out_p.n1067 out_p.n1066 0.151
R34858 out_p.n1068 out_p.n1067 0.151
R34859 out_p.n1069 out_p.n1068 0.151
R34860 out_p.n1070 out_p.n1069 0.151
R34861 out_p.n1071 out_p.n1070 0.151
R34862 out_p.n1072 out_p.n1071 0.151
R34863 out_p.n1073 out_p.n1072 0.151
R34864 out_p.n1074 out_p.n1073 0.151
R34865 out_p.n1075 out_p.n1074 0.151
R34866 out_p.n1076 out_p.n1075 0.151
R34867 out_p.n1077 out_p.n1076 0.151
R34868 out_p.n1078 out_p.n1077 0.151
R34869 out_p.n1079 out_p.n1078 0.151
R34870 out_p.n1080 out_p.n1079 0.151
R34871 out_p.n1081 out_p.n1080 0.151
R34872 out_p.n1082 out_p.n1081 0.151
R34873 out_p.n1083 out_p.n1082 0.151
R34874 out_p.n1084 out_p.n1083 0.151
R34875 out_p.n1090 out_p.n1089 0.151
R34876 out_p.n1091 out_p.n1090 0.151
R34877 out_p.n1092 out_p.n1091 0.151
R34878 out_p.n1093 out_p.n1092 0.151
R34879 out_p.n1094 out_p.n1093 0.151
R34880 out_p.n1095 out_p.n1094 0.151
R34881 out_p.n1096 out_p.n1095 0.151
R34882 out_p.n1097 out_p.n1096 0.151
R34883 out_p.n1098 out_p.n1097 0.151
R34884 out_p.n1099 out_p.n1098 0.151
R34885 out_p.n1100 out_p.n1099 0.151
R34886 out_p.n1101 out_p.n1100 0.151
R34887 out_p.n1102 out_p.n1101 0.151
R34888 out_p.n1103 out_p.n1102 0.151
R34889 out_p.n1104 out_p.n1103 0.151
R34890 out_p.n1105 out_p.n1104 0.151
R34891 out_p.n1106 out_p.n1105 0.151
R34892 out_p.n1107 out_p.n1106 0.151
R34893 out_p.n1108 out_p.n1107 0.151
R34894 out_p.n1114 out_p.n1113 0.151
R34895 out_p.n1115 out_p.n1114 0.151
R34896 out_p.n1116 out_p.n1115 0.151
R34897 out_p.n1117 out_p.n1116 0.151
R34898 out_p.n1118 out_p.n1117 0.151
R34899 out_p.n1119 out_p.n1118 0.151
R34900 out_p.n1120 out_p.n1119 0.151
R34901 out_p.n1121 out_p.n1120 0.151
R34902 out_p.n1122 out_p.n1121 0.151
R34903 out_p.n1123 out_p.n1122 0.151
R34904 out_p.n1124 out_p.n1123 0.151
R34905 out_p.n1125 out_p.n1124 0.151
R34906 out_p.n1126 out_p.n1125 0.151
R34907 out_p.n1127 out_p.n1126 0.151
R34908 out_p.n1128 out_p.n1127 0.151
R34909 out_p.n1129 out_p.n1128 0.151
R34910 out_p.n1130 out_p.n1129 0.151
R34911 out_p.n1131 out_p.n1130 0.151
R34912 out_p.n1132 out_p.n1131 0.151
R34913 out_p.n1138 out_p.n1137 0.151
R34914 out_p.n1139 out_p.n1138 0.151
R34915 out_p.n1140 out_p.n1139 0.151
R34916 out_p.n1141 out_p.n1140 0.151
R34917 out_p.n1142 out_p.n1141 0.151
R34918 out_p.n1143 out_p.n1142 0.151
R34919 out_p.n1144 out_p.n1143 0.151
R34920 out_p.n1145 out_p.n1144 0.151
R34921 out_p.n1146 out_p.n1145 0.151
R34922 out_p.n1147 out_p.n1146 0.151
R34923 out_p.n1148 out_p.n1147 0.151
R34924 out_p.n1149 out_p.n1148 0.151
R34925 out_p.n1150 out_p.n1149 0.151
R34926 out_p.n1151 out_p.n1150 0.151
R34927 out_p.n1152 out_p.n1151 0.151
R34928 out_p.n1153 out_p.n1152 0.151
R34929 out_p.n1154 out_p.n1153 0.151
R34930 out_p.n1155 out_p.n1154 0.151
R34931 out_p.n1156 out_p.n1155 0.151
R34932 out_p.n1162 out_p.n1161 0.151
R34933 out_p.n1163 out_p.n1162 0.151
R34934 out_p.n1164 out_p.n1163 0.151
R34935 out_p.n1165 out_p.n1164 0.151
R34936 out_p.n1166 out_p.n1165 0.151
R34937 out_p.n1167 out_p.n1166 0.151
R34938 out_p.n1168 out_p.n1167 0.151
R34939 out_p.n1169 out_p.n1168 0.151
R34940 out_p.n1170 out_p.n1169 0.151
R34941 out_p.n1171 out_p.n1170 0.151
R34942 out_p.n1172 out_p.n1171 0.151
R34943 out_p.n1173 out_p.n1172 0.151
R34944 out_p.n1174 out_p.n1173 0.151
R34945 out_p.n1175 out_p.n1174 0.151
R34946 out_p.n1176 out_p.n1175 0.151
R34947 out_p.n1177 out_p.n1176 0.151
R34948 out_p.n1178 out_p.n1177 0.151
R34949 out_p.n1179 out_p.n1178 0.151
R34950 out_p.n1180 out_p.n1179 0.151
R34951 out_p.n1186 out_p.n1185 0.151
R34952 out_p.n1187 out_p.n1186 0.151
R34953 out_p.n1188 out_p.n1187 0.151
R34954 out_p.n1189 out_p.n1188 0.151
R34955 out_p.n1190 out_p.n1189 0.151
R34956 out_p.n1191 out_p.n1190 0.151
R34957 out_p.n1192 out_p.n1191 0.151
R34958 out_p.n1193 out_p.n1192 0.151
R34959 out_p.n1194 out_p.n1193 0.151
R34960 out_p.n1195 out_p.n1194 0.151
R34961 out_p.n1196 out_p.n1195 0.151
R34962 out_p.n1197 out_p.n1196 0.151
R34963 out_p.n1198 out_p.n1197 0.151
R34964 out_p.n1199 out_p.n1198 0.151
R34965 out_p.n1200 out_p.n1199 0.151
R34966 out_p.n1201 out_p.n1200 0.151
R34967 out_p.n1202 out_p.n1201 0.151
R34968 out_p.n1203 out_p.n1202 0.151
R34969 out_p.n1204 out_p.n1203 0.151
R34970 out_p.n1210 out_p.n1209 0.151
R34971 out_p.n1211 out_p.n1210 0.151
R34972 out_p.n1212 out_p.n1211 0.151
R34973 out_p.n1213 out_p.n1212 0.151
R34974 out_p.n1214 out_p.n1213 0.151
R34975 out_p.n1215 out_p.n1214 0.151
R34976 out_p.n1216 out_p.n1215 0.151
R34977 out_p.n1217 out_p.n1216 0.151
R34978 out_p.n1218 out_p.n1217 0.151
R34979 out_p.n1219 out_p.n1218 0.151
R34980 out_p.n1220 out_p.n1219 0.151
R34981 out_p.n1221 out_p.n1220 0.151
R34982 out_p.n1222 out_p.n1221 0.151
R34983 out_p.n1223 out_p.n1222 0.151
R34984 out_p.n1224 out_p.n1223 0.151
R34985 out_p.n1225 out_p.n1224 0.151
R34986 out_p.n1226 out_p.n1225 0.151
R34987 out_p.n1227 out_p.n1226 0.151
R34988 out_p.n1228 out_p.n1227 0.151
R34989 out_p.n1234 out_p.n1233 0.151
R34990 out_p.n1235 out_p.n1234 0.151
R34991 out_p.n1236 out_p.n1235 0.151
R34992 out_p.n1237 out_p.n1236 0.151
R34993 out_p.n1238 out_p.n1237 0.151
R34994 out_p.n1239 out_p.n1238 0.151
R34995 out_p.n1240 out_p.n1239 0.151
R34996 out_p.n1241 out_p.n1240 0.151
R34997 out_p.n1242 out_p.n1241 0.151
R34998 out_p.n1243 out_p.n1242 0.151
R34999 out_p.n1244 out_p.n1243 0.151
R35000 out_p.n1245 out_p.n1244 0.151
R35001 out_p.n1246 out_p.n1245 0.151
R35002 out_p.n1247 out_p.n1246 0.151
R35003 out_p.n1248 out_p.n1247 0.151
R35004 out_p.n1249 out_p.n1248 0.151
R35005 out_p.n1250 out_p.n1249 0.151
R35006 out_p.n1251 out_p.n1250 0.151
R35007 out_p.n1252 out_p.n1251 0.151
R35008 out_p.n1258 out_p.n1257 0.151
R35009 out_p.n1259 out_p.n1258 0.151
R35010 out_p.n1260 out_p.n1259 0.151
R35011 out_p.n1261 out_p.n1260 0.151
R35012 out_p.n1262 out_p.n1261 0.151
R35013 out_p.n1263 out_p.n1262 0.151
R35014 out_p.n1264 out_p.n1263 0.151
R35015 out_p.n1265 out_p.n1264 0.151
R35016 out_p.n1266 out_p.n1265 0.151
R35017 out_p.n1267 out_p.n1266 0.151
R35018 out_p.n1268 out_p.n1267 0.151
R35019 out_p.n1269 out_p.n1268 0.151
R35020 out_p.n1270 out_p.n1269 0.151
R35021 out_p.n1271 out_p.n1270 0.151
R35022 out_p.n1272 out_p.n1271 0.151
R35023 out_p.n1273 out_p.n1272 0.151
R35024 out_p.n1274 out_p.n1273 0.151
R35025 out_p.n1275 out_p.n1274 0.151
R35026 out_p.n1276 out_p.n1275 0.151
R35027 out_p.n1282 out_p.n1281 0.151
R35028 out_p.n1283 out_p.n1282 0.151
R35029 out_p.n1284 out_p.n1283 0.151
R35030 out_p.n1285 out_p.n1284 0.151
R35031 out_p.n1286 out_p.n1285 0.151
R35032 out_p.n1287 out_p.n1286 0.151
R35033 out_p.n1288 out_p.n1287 0.151
R35034 out_p.n1289 out_p.n1288 0.151
R35035 out_p.n1290 out_p.n1289 0.151
R35036 out_p.n1291 out_p.n1290 0.151
R35037 out_p.n1292 out_p.n1291 0.151
R35038 out_p.n1293 out_p.n1292 0.151
R35039 out_p.n1294 out_p.n1293 0.151
R35040 out_p.n1295 out_p.n1294 0.151
R35041 out_p.n1296 out_p.n1295 0.151
R35042 out_p.n1297 out_p.n1296 0.151
R35043 out_p.n1298 out_p.n1297 0.151
R35044 out_p.n1299 out_p.n1298 0.151
R35045 out_p.n1300 out_p.n1299 0.151
R35046 out_p.n1306 out_p.n1305 0.151
R35047 out_p.n1307 out_p.n1306 0.151
R35048 out_p.n1308 out_p.n1307 0.151
R35049 out_p.n1309 out_p.n1308 0.151
R35050 out_p.n1310 out_p.n1309 0.151
R35051 out_p.n1311 out_p.n1310 0.151
R35052 out_p.n1312 out_p.n1311 0.151
R35053 out_p.n1313 out_p.n1312 0.151
R35054 out_p.n1314 out_p.n1313 0.151
R35055 out_p.n1315 out_p.n1314 0.151
R35056 out_p.n1316 out_p.n1315 0.151
R35057 out_p.n1317 out_p.n1316 0.151
R35058 out_p.n1318 out_p.n1317 0.151
R35059 out_p.n1319 out_p.n1318 0.151
R35060 out_p.n1320 out_p.n1319 0.151
R35061 out_p.n1321 out_p.n1320 0.151
R35062 out_p.n1322 out_p.n1321 0.151
R35063 out_p.n1323 out_p.n1322 0.151
R35064 out_p.n1324 out_p.n1323 0.151
R35065 out_p.n1330 out_p.n1329 0.151
R35066 out_p.n1331 out_p.n1330 0.151
R35067 out_p.n1332 out_p.n1331 0.151
R35068 out_p.n1333 out_p.n1332 0.151
R35069 out_p.n1334 out_p.n1333 0.151
R35070 out_p.n1335 out_p.n1334 0.151
R35071 out_p.n1336 out_p.n1335 0.151
R35072 out_p.n1337 out_p.n1336 0.151
R35073 out_p.n1338 out_p.n1337 0.151
R35074 out_p.n1339 out_p.n1338 0.151
R35075 out_p.n1340 out_p.n1339 0.151
R35076 out_p.n1341 out_p.n1340 0.151
R35077 out_p.n1342 out_p.n1341 0.151
R35078 out_p.n1343 out_p.n1342 0.151
R35079 out_p.n1344 out_p.n1343 0.151
R35080 out_p.n1345 out_p.n1344 0.151
R35081 out_p.n1346 out_p.n1345 0.151
R35082 out_p.n1347 out_p.n1346 0.151
R35083 out_p.n1348 out_p.n1347 0.151
R35084 out_p.n1354 out_p.n1353 0.151
R35085 out_p.n1355 out_p.n1354 0.151
R35086 out_p.n1356 out_p.n1355 0.151
R35087 out_p.n1357 out_p.n1356 0.151
R35088 out_p.n1358 out_p.n1357 0.151
R35089 out_p.n1359 out_p.n1358 0.151
R35090 out_p.n1360 out_p.n1359 0.151
R35091 out_p.n1361 out_p.n1360 0.151
R35092 out_p.n1362 out_p.n1361 0.151
R35093 out_p.n1363 out_p.n1362 0.151
R35094 out_p.n1364 out_p.n1363 0.151
R35095 out_p.n1365 out_p.n1364 0.151
R35096 out_p.n1366 out_p.n1365 0.151
R35097 out_p.n1367 out_p.n1366 0.151
R35098 out_p.n1368 out_p.n1367 0.151
R35099 out_p.n1369 out_p.n1368 0.151
R35100 out_p.n1370 out_p.n1369 0.151
R35101 out_p.n1371 out_p.n1370 0.151
R35102 out_p.n1372 out_p.n1371 0.151
R35103 out_p.n1378 out_p.n1377 0.151
R35104 out_p.n1379 out_p.n1378 0.151
R35105 out_p.n1380 out_p.n1379 0.151
R35106 out_p.n1381 out_p.n1380 0.151
R35107 out_p.n1382 out_p.n1381 0.151
R35108 out_p.n1383 out_p.n1382 0.151
R35109 out_p.n1384 out_p.n1383 0.151
R35110 out_p.n1385 out_p.n1384 0.151
R35111 out_p.n1386 out_p.n1385 0.151
R35112 out_p.n1387 out_p.n1386 0.151
R35113 out_p.n1388 out_p.n1387 0.151
R35114 out_p.n1389 out_p.n1388 0.151
R35115 out_p.n1390 out_p.n1389 0.151
R35116 out_p.n1391 out_p.n1390 0.151
R35117 out_p.n1392 out_p.n1391 0.151
R35118 out_p.n1393 out_p.n1392 0.151
R35119 out_p.n1394 out_p.n1393 0.151
R35120 out_p.n1395 out_p.n1394 0.151
R35121 out_p.n1396 out_p.n1395 0.151
R35122 out_p.n1402 out_p.n1401 0.151
R35123 out_p.n1403 out_p.n1402 0.151
R35124 out_p.n1404 out_p.n1403 0.151
R35125 out_p.n1405 out_p.n1404 0.151
R35126 out_p.n1406 out_p.n1405 0.151
R35127 out_p.n1407 out_p.n1406 0.151
R35128 out_p.n1408 out_p.n1407 0.151
R35129 out_p.n1409 out_p.n1408 0.151
R35130 out_p.n1410 out_p.n1409 0.151
R35131 out_p.n1411 out_p.n1410 0.151
R35132 out_p.n1412 out_p.n1411 0.151
R35133 out_p.n1413 out_p.n1412 0.151
R35134 out_p.n1414 out_p.n1413 0.151
R35135 out_p.n1415 out_p.n1414 0.151
R35136 out_p.n1416 out_p.n1415 0.151
R35137 out_p.n1417 out_p.n1416 0.151
R35138 out_p.n1418 out_p.n1417 0.151
R35139 out_p.n1419 out_p.n1418 0.151
R35140 out_p.n1420 out_p.n1419 0.151
R35141 out_p.n1426 out_p.n1425 0.151
R35142 out_p.n1427 out_p.n1426 0.151
R35143 out_p.n1428 out_p.n1427 0.151
R35144 out_p.n1429 out_p.n1428 0.151
R35145 out_p.n1430 out_p.n1429 0.151
R35146 out_p.n1431 out_p.n1430 0.151
R35147 out_p.n1432 out_p.n1431 0.151
R35148 out_p.n1433 out_p.n1432 0.151
R35149 out_p.n1434 out_p.n1433 0.151
R35150 out_p.n1435 out_p.n1434 0.151
R35151 out_p.n1436 out_p.n1435 0.151
R35152 out_p.n1437 out_p.n1436 0.151
R35153 out_p.n1438 out_p.n1437 0.151
R35154 out_p.n1439 out_p.n1438 0.151
R35155 out_p.n1440 out_p.n1439 0.151
R35156 out_p.n1441 out_p.n1440 0.151
R35157 out_p.n1442 out_p.n1441 0.151
R35158 out_p.n1443 out_p.n1442 0.151
R35159 out_p.n1444 out_p.n1443 0.151
R35160 out_p.n1450 out_p.n1449 0.151
R35161 out_p.n1451 out_p.n1450 0.151
R35162 out_p.n1452 out_p.n1451 0.151
R35163 out_p.n1453 out_p.n1452 0.151
R35164 out_p.n1454 out_p.n1453 0.151
R35165 out_p.n1455 out_p.n1454 0.151
R35166 out_p.n1456 out_p.n1455 0.151
R35167 out_p.n1457 out_p.n1456 0.151
R35168 out_p.n1458 out_p.n1457 0.151
R35169 out_p.n1459 out_p.n1458 0.151
R35170 out_p.n1460 out_p.n1459 0.151
R35171 out_p.n1461 out_p.n1460 0.151
R35172 out_p.n1462 out_p.n1461 0.151
R35173 out_p.n1463 out_p.n1462 0.151
R35174 out_p.n1464 out_p.n1463 0.151
R35175 out_p.n1465 out_p.n1464 0.151
R35176 out_p.n1466 out_p.n1465 0.151
R35177 out_p.n1467 out_p.n1466 0.151
R35178 out_p.n1468 out_p.n1467 0.151
R35179 out_p.n1474 out_p.n1473 0.151
R35180 out_p.n1475 out_p.n1474 0.151
R35181 out_p.n1476 out_p.n1475 0.151
R35182 out_p.n1477 out_p.n1476 0.151
R35183 out_p.n1478 out_p.n1477 0.151
R35184 out_p.n1479 out_p.n1478 0.151
R35185 out_p.n1480 out_p.n1479 0.151
R35186 out_p.n1481 out_p.n1480 0.151
R35187 out_p.n1482 out_p.n1481 0.151
R35188 out_p.n1483 out_p.n1482 0.151
R35189 out_p.n1484 out_p.n1483 0.151
R35190 out_p.n1485 out_p.n1484 0.151
R35191 out_p.n1486 out_p.n1485 0.151
R35192 out_p.n1487 out_p.n1486 0.151
R35193 out_p.n1488 out_p.n1487 0.151
R35194 out_p.n1489 out_p.n1488 0.151
R35195 out_p.n1490 out_p.n1489 0.151
R35196 out_p.n1491 out_p.n1490 0.151
R35197 out_p.n1492 out_p.n1491 0.151
R35198 out_p.n1498 out_p.n1497 0.151
R35199 out_p.n1499 out_p.n1498 0.151
R35200 out_p.n1500 out_p.n1499 0.151
R35201 out_p.n1501 out_p.n1500 0.151
R35202 out_p.n1502 out_p.n1501 0.151
R35203 out_p.n1503 out_p.n1502 0.151
R35204 out_p.n1504 out_p.n1503 0.151
R35205 out_p.n1505 out_p.n1504 0.151
R35206 out_p.n1506 out_p.n1505 0.151
R35207 out_p.n1507 out_p.n1506 0.151
R35208 out_p.n1508 out_p.n1507 0.151
R35209 out_p.n1509 out_p.n1508 0.151
R35210 out_p.n1510 out_p.n1509 0.151
R35211 out_p.n1511 out_p.n1510 0.151
R35212 out_p.n1512 out_p.n1511 0.151
R35213 out_p.n1513 out_p.n1512 0.151
R35214 out_p.n1514 out_p.n1513 0.151
R35215 out_p.n1515 out_p.n1514 0.151
R35216 out_p.n1516 out_p.n1515 0.151
R35217 out_p.n1522 out_p.n1521 0.151
R35218 out_p.n1523 out_p.n1522 0.151
R35219 out_p.n1524 out_p.n1523 0.151
R35220 out_p.n1525 out_p.n1524 0.151
R35221 out_p.n1526 out_p.n1525 0.151
R35222 out_p.n1527 out_p.n1526 0.151
R35223 out_p.n1528 out_p.n1527 0.151
R35224 out_p.n1529 out_p.n1528 0.151
R35225 out_p.n1530 out_p.n1529 0.151
R35226 out_p.n1531 out_p.n1530 0.151
R35227 out_p.n1532 out_p.n1531 0.151
R35228 out_p.n1533 out_p.n1532 0.151
R35229 out_p.n1534 out_p.n1533 0.151
R35230 out_p.n1535 out_p.n1534 0.151
R35231 out_p.n1536 out_p.n1535 0.151
R35232 out_p.n1537 out_p.n1536 0.151
R35233 out_p.n1538 out_p.n1537 0.151
R35234 out_p.n1539 out_p.n1538 0.151
R35235 out_p.n1540 out_p.n1539 0.151
R35236 out_p.n1546 out_p.n1545 0.151
R35237 out_p.n1547 out_p.n1546 0.151
R35238 out_p.n1548 out_p.n1547 0.151
R35239 out_p.n1549 out_p.n1548 0.151
R35240 out_p.n1550 out_p.n1549 0.151
R35241 out_p.n1551 out_p.n1550 0.151
R35242 out_p.n1552 out_p.n1551 0.151
R35243 out_p.n1553 out_p.n1552 0.151
R35244 out_p.n1554 out_p.n1553 0.151
R35245 out_p.n1555 out_p.n1554 0.151
R35246 out_p.n1556 out_p.n1555 0.151
R35247 out_p.n1557 out_p.n1556 0.151
R35248 out_p.n1558 out_p.n1557 0.151
R35249 out_p.n1559 out_p.n1558 0.151
R35250 out_p.n1560 out_p.n1559 0.151
R35251 out_p.n1561 out_p.n1560 0.151
R35252 out_p.n1562 out_p.n1561 0.151
R35253 out_p.n1563 out_p.n1562 0.151
R35254 out_p.n1564 out_p.n1563 0.151
R35255 out_p.n1570 out_p.n1569 0.151
R35256 out_p.n1571 out_p.n1570 0.151
R35257 out_p.n1572 out_p.n1571 0.151
R35258 out_p.n1573 out_p.n1572 0.151
R35259 out_p.n1574 out_p.n1573 0.151
R35260 out_p.n1575 out_p.n1574 0.151
R35261 out_p.n1576 out_p.n1575 0.151
R35262 out_p.n1577 out_p.n1576 0.151
R35263 out_p.n1578 out_p.n1577 0.151
R35264 out_p.n1579 out_p.n1578 0.151
R35265 out_p.n1580 out_p.n1579 0.151
R35266 out_p.n1581 out_p.n1580 0.151
R35267 out_p.n1582 out_p.n1581 0.151
R35268 out_p.n1583 out_p.n1582 0.151
R35269 out_p.n1584 out_p.n1583 0.151
R35270 out_p.n1585 out_p.n1584 0.151
R35271 out_p.n1586 out_p.n1585 0.151
R35272 out_p.n1587 out_p.n1586 0.151
R35273 out_p.n1588 out_p.n1587 0.151
R35274 out_p.n1594 out_p.n1593 0.151
R35275 out_p.n1595 out_p.n1594 0.151
R35276 out_p.n1596 out_p.n1595 0.151
R35277 out_p.n1597 out_p.n1596 0.151
R35278 out_p.n1598 out_p.n1597 0.151
R35279 out_p.n1599 out_p.n1598 0.151
R35280 out_p.n1600 out_p.n1599 0.151
R35281 out_p.n1601 out_p.n1600 0.151
R35282 out_p.n1602 out_p.n1601 0.151
R35283 out_p.n1603 out_p.n1602 0.151
R35284 out_p.n1604 out_p.n1603 0.151
R35285 out_p.n1605 out_p.n1604 0.151
R35286 out_p.n1606 out_p.n1605 0.151
R35287 out_p.n1607 out_p.n1606 0.151
R35288 out_p.n1608 out_p.n1607 0.151
R35289 out_p.n1609 out_p.n1608 0.151
R35290 out_p.n1610 out_p.n1609 0.151
R35291 out_p.n1611 out_p.n1610 0.151
R35292 out_p.n1612 out_p.n1611 0.151
R35293 out_p.n1618 out_p.n1617 0.151
R35294 out_p.n1619 out_p.n1618 0.151
R35295 out_p.n1620 out_p.n1619 0.151
R35296 out_p.n1621 out_p.n1620 0.151
R35297 out_p.n1622 out_p.n1621 0.151
R35298 out_p.n1623 out_p.n1622 0.151
R35299 out_p.n1624 out_p.n1623 0.151
R35300 out_p.n1625 out_p.n1624 0.151
R35301 out_p.n1626 out_p.n1625 0.151
R35302 out_p.n1627 out_p.n1626 0.151
R35303 out_p.n1628 out_p.n1627 0.151
R35304 out_p.n1629 out_p.n1628 0.151
R35305 out_p.n1630 out_p.n1629 0.151
R35306 out_p.n1631 out_p.n1630 0.151
R35307 out_p.n1632 out_p.n1631 0.151
R35308 out_p.n1633 out_p.n1632 0.151
R35309 out_p.n1634 out_p.n1633 0.151
R35310 out_p.n1635 out_p.n1634 0.151
R35311 out_p.n1636 out_p.n1635 0.151
R35312 out_p.n1642 out_p.n1641 0.151
R35313 out_p.n1643 out_p.n1642 0.151
R35314 out_p.n1644 out_p.n1643 0.151
R35315 out_p.n1645 out_p.n1644 0.151
R35316 out_p.n1646 out_p.n1645 0.151
R35317 out_p.n1647 out_p.n1646 0.151
R35318 out_p.n1648 out_p.n1647 0.151
R35319 out_p.n1649 out_p.n1648 0.151
R35320 out_p.n1650 out_p.n1649 0.151
R35321 out_p.n1651 out_p.n1650 0.151
R35322 out_p.n1652 out_p.n1651 0.151
R35323 out_p.n1653 out_p.n1652 0.151
R35324 out_p.n1654 out_p.n1653 0.151
R35325 out_p.n1655 out_p.n1654 0.151
R35326 out_p.n1656 out_p.n1655 0.151
R35327 out_p.n1657 out_p.n1656 0.151
R35328 out_p.n1658 out_p.n1657 0.151
R35329 out_p.n1659 out_p.n1658 0.151
R35330 out_p.n1660 out_p.n1659 0.151
R35331 out_p.n1666 out_p.n1665 0.151
R35332 out_p.n1667 out_p.n1666 0.151
R35333 out_p.n1668 out_p.n1667 0.151
R35334 out_p.n1669 out_p.n1668 0.151
R35335 out_p.n1670 out_p.n1669 0.151
R35336 out_p.n1671 out_p.n1670 0.151
R35337 out_p.n1672 out_p.n1671 0.151
R35338 out_p.n1673 out_p.n1672 0.151
R35339 out_p.n1674 out_p.n1673 0.151
R35340 out_p.n1675 out_p.n1674 0.151
R35341 out_p.n1676 out_p.n1675 0.151
R35342 out_p.n1677 out_p.n1676 0.151
R35343 out_p.n1678 out_p.n1677 0.151
R35344 out_p.n1679 out_p.n1678 0.151
R35345 out_p.n1680 out_p.n1679 0.151
R35346 out_p.n1681 out_p.n1680 0.151
R35347 out_p.n1682 out_p.n1681 0.151
R35348 out_p.n1683 out_p.n1682 0.151
R35349 out_p.n1684 out_p.n1683 0.151
R35350 out_p.n1690 out_p.n1689 0.151
R35351 out_p.n1691 out_p.n1690 0.151
R35352 out_p.n1692 out_p.n1691 0.151
R35353 out_p.n1693 out_p.n1692 0.151
R35354 out_p.n1694 out_p.n1693 0.151
R35355 out_p.n1695 out_p.n1694 0.151
R35356 out_p.n1696 out_p.n1695 0.151
R35357 out_p.n1697 out_p.n1696 0.151
R35358 out_p.n1698 out_p.n1697 0.151
R35359 out_p.n1699 out_p.n1698 0.151
R35360 out_p.n1700 out_p.n1699 0.151
R35361 out_p.n1701 out_p.n1700 0.151
R35362 out_p.n1702 out_p.n1701 0.151
R35363 out_p.n1703 out_p.n1702 0.151
R35364 out_p.n1704 out_p.n1703 0.151
R35365 out_p.n1705 out_p.n1704 0.151
R35366 out_p.n1706 out_p.n1705 0.151
R35367 out_p.n1707 out_p.n1706 0.151
R35368 out_p.n1708 out_p.n1707 0.151
R35369 out_p.n1714 out_p.n1713 0.151
R35370 out_p.n1715 out_p.n1714 0.151
R35371 out_p.n1716 out_p.n1715 0.151
R35372 out_p.n1717 out_p.n1716 0.151
R35373 out_p.n1718 out_p.n1717 0.151
R35374 out_p.n1719 out_p.n1718 0.151
R35375 out_p.n1720 out_p.n1719 0.151
R35376 out_p.n1721 out_p.n1720 0.151
R35377 out_p.n1722 out_p.n1721 0.151
R35378 out_p.n1723 out_p.n1722 0.151
R35379 out_p.n1724 out_p.n1723 0.151
R35380 out_p.n1725 out_p.n1724 0.151
R35381 out_p.n1726 out_p.n1725 0.151
R35382 out_p.n1727 out_p.n1726 0.151
R35383 out_p.n1728 out_p.n1727 0.151
R35384 out_p.n1729 out_p.n1728 0.151
R35385 out_p.n1730 out_p.n1729 0.151
R35386 out_p.n1731 out_p.n1730 0.151
R35387 out_p.n1732 out_p.n1731 0.151
R35388 out_p.n1738 out_p.n1737 0.151
R35389 out_p.n1739 out_p.n1738 0.151
R35390 out_p.n1740 out_p.n1739 0.151
R35391 out_p.n1741 out_p.n1740 0.151
R35392 out_p.n1742 out_p.n1741 0.151
R35393 out_p.n1743 out_p.n1742 0.151
R35394 out_p.n1744 out_p.n1743 0.151
R35395 out_p.n1745 out_p.n1744 0.151
R35396 out_p.n1746 out_p.n1745 0.151
R35397 out_p.n1747 out_p.n1746 0.151
R35398 out_p.n1748 out_p.n1747 0.151
R35399 out_p.n1749 out_p.n1748 0.151
R35400 out_p.n1750 out_p.n1749 0.151
R35401 out_p.n1751 out_p.n1750 0.151
R35402 out_p.n1752 out_p.n1751 0.151
R35403 out_p.n1753 out_p.n1752 0.151
R35404 out_p.n1754 out_p.n1753 0.151
R35405 out_p.n1755 out_p.n1754 0.151
R35406 out_p.n1756 out_p.n1755 0.151
R35407 out_p.n1762 out_p.n1761 0.151
R35408 out_p.n1763 out_p.n1762 0.151
R35409 out_p.n1764 out_p.n1763 0.151
R35410 out_p.n1765 out_p.n1764 0.151
R35411 out_p.n1766 out_p.n1765 0.151
R35412 out_p.n1767 out_p.n1766 0.151
R35413 out_p.n1768 out_p.n1767 0.151
R35414 out_p.n1769 out_p.n1768 0.151
R35415 out_p.n1770 out_p.n1769 0.151
R35416 out_p.n1771 out_p.n1770 0.151
R35417 out_p.n1772 out_p.n1771 0.151
R35418 out_p.n1773 out_p.n1772 0.151
R35419 out_p.n1774 out_p.n1773 0.151
R35420 out_p.n1775 out_p.n1774 0.151
R35421 out_p.n1776 out_p.n1775 0.151
R35422 out_p.n1777 out_p.n1776 0.151
R35423 out_p.n1778 out_p.n1777 0.151
R35424 out_p.n1779 out_p.n1778 0.151
R35425 out_p.n1780 out_p.n1779 0.151
R35426 out_p.n1786 out_p.n1785 0.151
R35427 out_p.n1787 out_p.n1786 0.151
R35428 out_p.n1788 out_p.n1787 0.151
R35429 out_p.n1789 out_p.n1788 0.151
R35430 out_p.n1790 out_p.n1789 0.151
R35431 out_p.n1791 out_p.n1790 0.151
R35432 out_p.n1792 out_p.n1791 0.151
R35433 out_p.n1793 out_p.n1792 0.151
R35434 out_p.n1794 out_p.n1793 0.151
R35435 out_p.n1795 out_p.n1794 0.151
R35436 out_p.n1796 out_p.n1795 0.151
R35437 out_p.n1797 out_p.n1796 0.151
R35438 out_p.n1798 out_p.n1797 0.151
R35439 out_p.n1799 out_p.n1798 0.151
R35440 out_p.n1800 out_p.n1799 0.151
R35441 out_p.n1801 out_p.n1800 0.151
R35442 out_p.n1802 out_p.n1801 0.151
R35443 out_p.n1803 out_p.n1802 0.151
R35444 out_p.n1804 out_p.n1803 0.151
R35445 out_p.n1810 out_p.n1809 0.151
R35446 out_p.n1811 out_p.n1810 0.151
R35447 out_p.n1812 out_p.n1811 0.151
R35448 out_p.n1813 out_p.n1812 0.151
R35449 out_p.n1814 out_p.n1813 0.151
R35450 out_p.n1815 out_p.n1814 0.151
R35451 out_p.n1816 out_p.n1815 0.151
R35452 out_p.n1817 out_p.n1816 0.151
R35453 out_p.n1818 out_p.n1817 0.151
R35454 out_p.n1819 out_p.n1818 0.151
R35455 out_p.n1820 out_p.n1819 0.151
R35456 out_p.n1821 out_p.n1820 0.151
R35457 out_p.n1822 out_p.n1821 0.151
R35458 out_p.n1823 out_p.n1822 0.151
R35459 out_p.n1824 out_p.n1823 0.151
R35460 out_p.n1825 out_p.n1824 0.151
R35461 out_p.n1826 out_p.n1825 0.151
R35462 out_p.n1827 out_p.n1826 0.151
R35463 out_p.n1828 out_p.n1827 0.151
R35464 out_p.n748 out_p.n747 0.148
R35465 out_p.n745 out_p.n744 0.148
R35466 out_p.n743 out_p.n742 0.144
R35467 out_p.n742 out_p.n741 0.144
R35468 out_p.n741 out_p.n740 0.144
R35469 out_p.n719 out_p.n718 0.144
R35470 out_p.n718 out_p.n717 0.144
R35471 out_p.n717 out_p.n716 0.144
R35472 out_p.n695 out_p.n694 0.144
R35473 out_p.n694 out_p.n693 0.144
R35474 out_p.n693 out_p.n692 0.144
R35475 out_p.n671 out_p.n670 0.144
R35476 out_p.n670 out_p.n669 0.144
R35477 out_p.n669 out_p.n668 0.144
R35478 out_p.n647 out_p.n646 0.144
R35479 out_p.n646 out_p.n645 0.144
R35480 out_p.n645 out_p.n644 0.144
R35481 out_p.n623 out_p.n622 0.144
R35482 out_p.n622 out_p.n621 0.144
R35483 out_p.n621 out_p.n620 0.144
R35484 out_p.n599 out_p.n598 0.144
R35485 out_p.n598 out_p.n597 0.144
R35486 out_p.n597 out_p.n596 0.144
R35487 out_p.n575 out_p.n574 0.144
R35488 out_p.n574 out_p.n573 0.144
R35489 out_p.n573 out_p.n572 0.144
R35490 out_p.n551 out_p.n550 0.144
R35491 out_p.n550 out_p.n549 0.144
R35492 out_p.n549 out_p.n548 0.144
R35493 out_p.n527 out_p.n526 0.144
R35494 out_p.n526 out_p.n525 0.144
R35495 out_p.n525 out_p.n524 0.144
R35496 out_p.n503 out_p.n502 0.144
R35497 out_p.n502 out_p.n501 0.144
R35498 out_p.n501 out_p.n500 0.144
R35499 out_p.n479 out_p.n478 0.144
R35500 out_p.n478 out_p.n477 0.144
R35501 out_p.n477 out_p.n476 0.144
R35502 out_p.n455 out_p.n454 0.144
R35503 out_p.n454 out_p.n453 0.144
R35504 out_p.n453 out_p.n452 0.144
R35505 out_p.n431 out_p.n430 0.144
R35506 out_p.n430 out_p.n429 0.144
R35507 out_p.n429 out_p.n428 0.144
R35508 out_p.n407 out_p.n406 0.144
R35509 out_p.n406 out_p.n405 0.144
R35510 out_p.n405 out_p.n404 0.144
R35511 out_p.n383 out_p.n382 0.144
R35512 out_p.n382 out_p.n381 0.144
R35513 out_p.n381 out_p.n380 0.144
R35514 out_p.n359 out_p.n358 0.144
R35515 out_p.n358 out_p.n357 0.144
R35516 out_p.n357 out_p.n356 0.144
R35517 out_p.n335 out_p.n334 0.144
R35518 out_p.n334 out_p.n333 0.144
R35519 out_p.n333 out_p.n332 0.144
R35520 out_p.n311 out_p.n310 0.144
R35521 out_p.n310 out_p.n309 0.144
R35522 out_p.n309 out_p.n308 0.144
R35523 out_p.n287 out_p.n286 0.144
R35524 out_p.n286 out_p.n285 0.144
R35525 out_p.n285 out_p.n284 0.144
R35526 out_p.n263 out_p.n262 0.144
R35527 out_p.n262 out_p.n261 0.144
R35528 out_p.n261 out_p.n260 0.144
R35529 out_p.n239 out_p.n238 0.144
R35530 out_p.n238 out_p.n237 0.144
R35531 out_p.n237 out_p.n236 0.144
R35532 out_p.n215 out_p.n214 0.144
R35533 out_p.n214 out_p.n213 0.144
R35534 out_p.n213 out_p.n212 0.144
R35535 out_p.n191 out_p.n190 0.144
R35536 out_p.n190 out_p.n189 0.144
R35537 out_p.n189 out_p.n188 0.144
R35538 out_p.n167 out_p.n166 0.144
R35539 out_p.n166 out_p.n165 0.144
R35540 out_p.n165 out_p.n164 0.144
R35541 out_p.n143 out_p.n142 0.144
R35542 out_p.n142 out_p.n141 0.144
R35543 out_p.n141 out_p.n140 0.144
R35544 out_p.n119 out_p.n118 0.144
R35545 out_p.n118 out_p.n117 0.144
R35546 out_p.n117 out_p.n116 0.144
R35547 out_p.n95 out_p.n94 0.144
R35548 out_p.n94 out_p.n93 0.144
R35549 out_p.n93 out_p.n92 0.144
R35550 out_p.n71 out_p.n70 0.144
R35551 out_p.n70 out_p.n69 0.144
R35552 out_p.n69 out_p.n68 0.144
R35553 out_p.n47 out_p.n46 0.144
R35554 out_p.n46 out_p.n45 0.144
R35555 out_p.n45 out_p.n44 0.144
R35556 out_p.n23 out_p.n22 0.144
R35557 out_p.n22 out_p.n21 0.144
R35558 out_p.n21 out_p.n20 0.144
R35559 out_p.n804 out_p.n803 0.144
R35560 out_p.n803 out_p.n802 0.144
R35561 out_p.n802 out_p.n801 0.144
R35562 out_p.n848 out_p.n847 0.144
R35563 out_p.n847 out_p.n846 0.144
R35564 out_p.n846 out_p.n845 0.144
R35565 out_p.n872 out_p.n871 0.144
R35566 out_p.n871 out_p.n870 0.144
R35567 out_p.n870 out_p.n869 0.144
R35568 out_p.n896 out_p.n895 0.144
R35569 out_p.n895 out_p.n894 0.144
R35570 out_p.n894 out_p.n893 0.144
R35571 out_p.n920 out_p.n919 0.144
R35572 out_p.n919 out_p.n918 0.144
R35573 out_p.n918 out_p.n917 0.144
R35574 out_p.n944 out_p.n943 0.144
R35575 out_p.n943 out_p.n942 0.144
R35576 out_p.n942 out_p.n941 0.144
R35577 out_p.n968 out_p.n967 0.144
R35578 out_p.n967 out_p.n966 0.144
R35579 out_p.n966 out_p.n965 0.144
R35580 out_p.n992 out_p.n991 0.144
R35581 out_p.n991 out_p.n990 0.144
R35582 out_p.n990 out_p.n989 0.144
R35583 out_p.n1016 out_p.n1015 0.144
R35584 out_p.n1015 out_p.n1014 0.144
R35585 out_p.n1014 out_p.n1013 0.144
R35586 out_p.n1040 out_p.n1039 0.144
R35587 out_p.n1039 out_p.n1038 0.144
R35588 out_p.n1038 out_p.n1037 0.144
R35589 out_p.n1064 out_p.n1063 0.144
R35590 out_p.n1063 out_p.n1062 0.144
R35591 out_p.n1062 out_p.n1061 0.144
R35592 out_p.n1088 out_p.n1087 0.144
R35593 out_p.n1087 out_p.n1086 0.144
R35594 out_p.n1086 out_p.n1085 0.144
R35595 out_p.n1112 out_p.n1111 0.144
R35596 out_p.n1111 out_p.n1110 0.144
R35597 out_p.n1110 out_p.n1109 0.144
R35598 out_p.n1136 out_p.n1135 0.144
R35599 out_p.n1135 out_p.n1134 0.144
R35600 out_p.n1134 out_p.n1133 0.144
R35601 out_p.n1160 out_p.n1159 0.144
R35602 out_p.n1159 out_p.n1158 0.144
R35603 out_p.n1158 out_p.n1157 0.144
R35604 out_p.n1184 out_p.n1183 0.144
R35605 out_p.n1183 out_p.n1182 0.144
R35606 out_p.n1182 out_p.n1181 0.144
R35607 out_p.n1208 out_p.n1207 0.144
R35608 out_p.n1207 out_p.n1206 0.144
R35609 out_p.n1206 out_p.n1205 0.144
R35610 out_p.n1232 out_p.n1231 0.144
R35611 out_p.n1231 out_p.n1230 0.144
R35612 out_p.n1230 out_p.n1229 0.144
R35613 out_p.n1256 out_p.n1255 0.144
R35614 out_p.n1255 out_p.n1254 0.144
R35615 out_p.n1254 out_p.n1253 0.144
R35616 out_p.n1280 out_p.n1279 0.144
R35617 out_p.n1279 out_p.n1278 0.144
R35618 out_p.n1278 out_p.n1277 0.144
R35619 out_p.n1304 out_p.n1303 0.144
R35620 out_p.n1303 out_p.n1302 0.144
R35621 out_p.n1302 out_p.n1301 0.144
R35622 out_p.n1328 out_p.n1327 0.144
R35623 out_p.n1327 out_p.n1326 0.144
R35624 out_p.n1326 out_p.n1325 0.144
R35625 out_p.n1352 out_p.n1351 0.144
R35626 out_p.n1351 out_p.n1350 0.144
R35627 out_p.n1350 out_p.n1349 0.144
R35628 out_p.n1376 out_p.n1375 0.144
R35629 out_p.n1375 out_p.n1374 0.144
R35630 out_p.n1374 out_p.n1373 0.144
R35631 out_p.n1400 out_p.n1399 0.144
R35632 out_p.n1399 out_p.n1398 0.144
R35633 out_p.n1398 out_p.n1397 0.144
R35634 out_p.n1424 out_p.n1423 0.144
R35635 out_p.n1423 out_p.n1422 0.144
R35636 out_p.n1422 out_p.n1421 0.144
R35637 out_p.n1448 out_p.n1447 0.144
R35638 out_p.n1447 out_p.n1446 0.144
R35639 out_p.n1446 out_p.n1445 0.144
R35640 out_p.n1472 out_p.n1471 0.144
R35641 out_p.n1471 out_p.n1470 0.144
R35642 out_p.n1470 out_p.n1469 0.144
R35643 out_p.n1496 out_p.n1495 0.144
R35644 out_p.n1495 out_p.n1494 0.144
R35645 out_p.n1494 out_p.n1493 0.144
R35646 out_p.n1520 out_p.n1519 0.144
R35647 out_p.n1519 out_p.n1518 0.144
R35648 out_p.n1518 out_p.n1517 0.144
R35649 out_p.n1544 out_p.n1543 0.144
R35650 out_p.n1543 out_p.n1542 0.144
R35651 out_p.n1542 out_p.n1541 0.144
R35652 out_p.n1568 out_p.n1567 0.144
R35653 out_p.n1567 out_p.n1566 0.144
R35654 out_p.n1566 out_p.n1565 0.144
R35655 out_p.n1592 out_p.n1591 0.144
R35656 out_p.n1591 out_p.n1590 0.144
R35657 out_p.n1590 out_p.n1589 0.144
R35658 out_p.n1616 out_p.n1615 0.144
R35659 out_p.n1615 out_p.n1614 0.144
R35660 out_p.n1614 out_p.n1613 0.144
R35661 out_p.n1640 out_p.n1639 0.144
R35662 out_p.n1639 out_p.n1638 0.144
R35663 out_p.n1638 out_p.n1637 0.144
R35664 out_p.n1664 out_p.n1663 0.144
R35665 out_p.n1663 out_p.n1662 0.144
R35666 out_p.n1662 out_p.n1661 0.144
R35667 out_p.n1688 out_p.n1687 0.144
R35668 out_p.n1687 out_p.n1686 0.144
R35669 out_p.n1686 out_p.n1685 0.144
R35670 out_p.n1712 out_p.n1711 0.144
R35671 out_p.n1711 out_p.n1710 0.144
R35672 out_p.n1710 out_p.n1709 0.144
R35673 out_p.n1736 out_p.n1735 0.144
R35674 out_p.n1735 out_p.n1734 0.144
R35675 out_p.n1734 out_p.n1733 0.144
R35676 out_p.n1760 out_p.n1759 0.144
R35677 out_p.n1759 out_p.n1758 0.144
R35678 out_p.n1758 out_p.n1757 0.144
R35679 out_p.n1784 out_p.n1783 0.144
R35680 out_p.n1783 out_p.n1782 0.144
R35681 out_p.n1782 out_p.n1781 0.144
R35682 out_p.n1808 out_p.n1807 0.144
R35683 out_p.n1807 out_p.n1806 0.144
R35684 out_p.n1806 out_p.n1805 0.144
R35685 out_p.n1832 out_p.n1831 0.144
R35686 out_p.n1831 out_p.n1830 0.144
R35687 out_p.n1830 out_p.n1829 0.144
R35688 out_p.n769 out_p.n768 0.093
R35689 out_p.n770 out_p.n739 0.093
R35690 out_p.n771 out_p.n715 0.093
R35691 out_p.n772 out_p.n691 0.093
R35692 out_p.n773 out_p.n667 0.093
R35693 out_p.n774 out_p.n643 0.093
R35694 out_p.n775 out_p.n619 0.093
R35695 out_p.n776 out_p.n595 0.093
R35696 out_p.n777 out_p.n571 0.093
R35697 out_p.n778 out_p.n547 0.093
R35698 out_p.n779 out_p.n523 0.093
R35699 out_p.n780 out_p.n499 0.093
R35700 out_p.n781 out_p.n475 0.093
R35701 out_p.n782 out_p.n451 0.093
R35702 out_p.n783 out_p.n427 0.093
R35703 out_p.n784 out_p.n403 0.093
R35704 out_p.n785 out_p.n379 0.093
R35705 out_p.n786 out_p.n355 0.093
R35706 out_p.n787 out_p.n331 0.093
R35707 out_p.n788 out_p.n307 0.093
R35708 out_p.n789 out_p.n283 0.093
R35709 out_p.n790 out_p.n259 0.093
R35710 out_p.n791 out_p.n235 0.093
R35711 out_p.n792 out_p.n211 0.093
R35712 out_p.n793 out_p.n187 0.093
R35713 out_p.n794 out_p.n163 0.093
R35714 out_p.n795 out_p.n139 0.093
R35715 out_p.n796 out_p.n115 0.093
R35716 out_p.n797 out_p.n91 0.093
R35717 out_p.n798 out_p.n67 0.093
R35718 out_p.n799 out_p.n43 0.093
R35719 out_p.n800 out_p.n19 0.093
R35720 out_p out_p.n824 0.093
R35721 out_p.n1874 out_p.n844 0.093
R35722 out_p.n1873 out_p.n868 0.093
R35723 out_p.n1872 out_p.n892 0.093
R35724 out_p.n1871 out_p.n916 0.093
R35725 out_p.n1870 out_p.n940 0.093
R35726 out_p.n1869 out_p.n964 0.093
R35727 out_p.n1868 out_p.n988 0.093
R35728 out_p.n1867 out_p.n1012 0.093
R35729 out_p.n1866 out_p.n1036 0.093
R35730 out_p.n1865 out_p.n1060 0.093
R35731 out_p.n1864 out_p.n1084 0.093
R35732 out_p.n1863 out_p.n1108 0.093
R35733 out_p.n1862 out_p.n1132 0.093
R35734 out_p.n1861 out_p.n1156 0.093
R35735 out_p.n1860 out_p.n1180 0.093
R35736 out_p.n1859 out_p.n1204 0.093
R35737 out_p.n1858 out_p.n1228 0.093
R35738 out_p.n1857 out_p.n1252 0.093
R35739 out_p.n1856 out_p.n1276 0.093
R35740 out_p.n1855 out_p.n1300 0.093
R35741 out_p.n1854 out_p.n1324 0.093
R35742 out_p.n1853 out_p.n1348 0.093
R35743 out_p.n1852 out_p.n1372 0.093
R35744 out_p.n1851 out_p.n1396 0.093
R35745 out_p.n1850 out_p.n1420 0.093
R35746 out_p.n1849 out_p.n1444 0.093
R35747 out_p.n1848 out_p.n1468 0.093
R35748 out_p.n1847 out_p.n1492 0.093
R35749 out_p.n1846 out_p.n1516 0.093
R35750 out_p.n1845 out_p.n1540 0.093
R35751 out_p.n1844 out_p.n1564 0.093
R35752 out_p.n1843 out_p.n1588 0.093
R35753 out_p.n1842 out_p.n1612 0.093
R35754 out_p.n1841 out_p.n1636 0.093
R35755 out_p.n1840 out_p.n1660 0.093
R35756 out_p.n1839 out_p.n1684 0.093
R35757 out_p.n1838 out_p.n1708 0.093
R35758 out_p.n1837 out_p.n1732 0.093
R35759 out_p.n1836 out_p.n1756 0.093
R35760 out_p.n1835 out_p.n1780 0.093
R35761 out_p.n1834 out_p.n1804 0.093
R35762 out_p.n1833 out_p.n1828 0.093
R35763 out_p.n769 out_p.n748 0.093
R35764 out_p.n746 out_p.n745 0.092
R35765 out_p.n770 out_p.n743 0.091
R35766 out_p.n771 out_p.n719 0.091
R35767 out_p.n772 out_p.n695 0.091
R35768 out_p.n773 out_p.n671 0.091
R35769 out_p.n774 out_p.n647 0.091
R35770 out_p.n775 out_p.n623 0.091
R35771 out_p.n776 out_p.n599 0.091
R35772 out_p.n777 out_p.n575 0.091
R35773 out_p.n778 out_p.n551 0.091
R35774 out_p.n779 out_p.n527 0.091
R35775 out_p.n780 out_p.n503 0.091
R35776 out_p.n781 out_p.n479 0.091
R35777 out_p.n782 out_p.n455 0.091
R35778 out_p.n783 out_p.n431 0.091
R35779 out_p.n784 out_p.n407 0.091
R35780 out_p.n785 out_p.n383 0.091
R35781 out_p.n786 out_p.n359 0.091
R35782 out_p.n787 out_p.n335 0.091
R35783 out_p.n788 out_p.n311 0.091
R35784 out_p.n789 out_p.n287 0.091
R35785 out_p.n790 out_p.n263 0.091
R35786 out_p.n791 out_p.n239 0.091
R35787 out_p.n792 out_p.n215 0.091
R35788 out_p.n793 out_p.n191 0.091
R35789 out_p.n794 out_p.n167 0.091
R35790 out_p.n795 out_p.n143 0.091
R35791 out_p.n796 out_p.n119 0.091
R35792 out_p.n797 out_p.n95 0.091
R35793 out_p.n798 out_p.n71 0.091
R35794 out_p.n799 out_p.n47 0.091
R35795 out_p.n800 out_p.n23 0.091
R35796 out_p out_p.n804 0.091
R35797 out_p.n1874 out_p.n848 0.091
R35798 out_p.n1873 out_p.n872 0.091
R35799 out_p.n1872 out_p.n896 0.091
R35800 out_p.n1871 out_p.n920 0.091
R35801 out_p.n1870 out_p.n944 0.091
R35802 out_p.n1869 out_p.n968 0.091
R35803 out_p.n1868 out_p.n992 0.091
R35804 out_p.n1867 out_p.n1016 0.091
R35805 out_p.n1866 out_p.n1040 0.091
R35806 out_p.n1865 out_p.n1064 0.091
R35807 out_p.n1864 out_p.n1088 0.091
R35808 out_p.n1863 out_p.n1112 0.091
R35809 out_p.n1862 out_p.n1136 0.091
R35810 out_p.n1861 out_p.n1160 0.091
R35811 out_p.n1860 out_p.n1184 0.091
R35812 out_p.n1859 out_p.n1208 0.091
R35813 out_p.n1858 out_p.n1232 0.091
R35814 out_p.n1857 out_p.n1256 0.091
R35815 out_p.n1856 out_p.n1280 0.091
R35816 out_p.n1855 out_p.n1304 0.091
R35817 out_p.n1854 out_p.n1328 0.091
R35818 out_p.n1853 out_p.n1352 0.091
R35819 out_p.n1852 out_p.n1376 0.091
R35820 out_p.n1851 out_p.n1400 0.091
R35821 out_p.n1850 out_p.n1424 0.091
R35822 out_p.n1849 out_p.n1448 0.091
R35823 out_p.n1848 out_p.n1472 0.091
R35824 out_p.n1847 out_p.n1496 0.091
R35825 out_p.n1846 out_p.n1520 0.091
R35826 out_p.n1845 out_p.n1544 0.091
R35827 out_p.n1844 out_p.n1568 0.091
R35828 out_p.n1843 out_p.n1592 0.091
R35829 out_p.n1842 out_p.n1616 0.091
R35830 out_p.n1841 out_p.n1640 0.091
R35831 out_p.n1840 out_p.n1664 0.091
R35832 out_p.n1839 out_p.n1688 0.091
R35833 out_p.n1838 out_p.n1712 0.091
R35834 out_p.n1837 out_p.n1736 0.091
R35835 out_p.n1836 out_p.n1760 0.091
R35836 out_p.n1835 out_p.n1784 0.091
R35837 out_p.n1834 out_p.n1808 0.091
R35838 out_p.n1833 out_p.n1832 0.091
R35839 out_p.n747 out_p.n746 0.056
R35840 out_p.n770 out_p.n769 0.001
R35841 out_p.n771 out_p.n770 0.001
R35842 out_p.n772 out_p.n771 0.001
R35843 out_p.n773 out_p.n772 0.001
R35844 out_p.n774 out_p.n773 0.001
R35845 out_p.n775 out_p.n774 0.001
R35846 out_p.n776 out_p.n775 0.001
R35847 out_p.n777 out_p.n776 0.001
R35848 out_p.n778 out_p.n777 0.001
R35849 out_p.n779 out_p.n778 0.001
R35850 out_p.n780 out_p.n779 0.001
R35851 out_p.n781 out_p.n780 0.001
R35852 out_p.n782 out_p.n781 0.001
R35853 out_p.n783 out_p.n782 0.001
R35854 out_p.n784 out_p.n783 0.001
R35855 out_p.n785 out_p.n784 0.001
R35856 out_p.n786 out_p.n785 0.001
R35857 out_p.n787 out_p.n786 0.001
R35858 out_p.n788 out_p.n787 0.001
R35859 out_p.n789 out_p.n788 0.001
R35860 out_p.n790 out_p.n789 0.001
R35861 out_p.n791 out_p.n790 0.001
R35862 out_p.n792 out_p.n791 0.001
R35863 out_p.n793 out_p.n792 0.001
R35864 out_p.n794 out_p.n793 0.001
R35865 out_p.n795 out_p.n794 0.001
R35866 out_p.n796 out_p.n795 0.001
R35867 out_p.n797 out_p.n796 0.001
R35868 out_p.n798 out_p.n797 0.001
R35869 out_p.n799 out_p.n798 0.001
R35870 out_p.n800 out_p.n799 0.001
R35871 out_p out_p.n800 0.001
R35872 out_p out_p.n1874 0.001
R35873 out_p.n1874 out_p.n1873 0.001
R35874 out_p.n1873 out_p.n1872 0.001
R35875 out_p.n1872 out_p.n1871 0.001
R35876 out_p.n1871 out_p.n1870 0.001
R35877 out_p.n1870 out_p.n1869 0.001
R35878 out_p.n1869 out_p.n1868 0.001
R35879 out_p.n1868 out_p.n1867 0.001
R35880 out_p.n1867 out_p.n1866 0.001
R35881 out_p.n1866 out_p.n1865 0.001
R35882 out_p.n1865 out_p.n1864 0.001
R35883 out_p.n1864 out_p.n1863 0.001
R35884 out_p.n1863 out_p.n1862 0.001
R35885 out_p.n1862 out_p.n1861 0.001
R35886 out_p.n1861 out_p.n1860 0.001
R35887 out_p.n1860 out_p.n1859 0.001
R35888 out_p.n1859 out_p.n1858 0.001
R35889 out_p.n1858 out_p.n1857 0.001
R35890 out_p.n1857 out_p.n1856 0.001
R35891 out_p.n1856 out_p.n1855 0.001
R35892 out_p.n1855 out_p.n1854 0.001
R35893 out_p.n1854 out_p.n1853 0.001
R35894 out_p.n1853 out_p.n1852 0.001
R35895 out_p.n1852 out_p.n1851 0.001
R35896 out_p.n1851 out_p.n1850 0.001
R35897 out_p.n1850 out_p.n1849 0.001
R35898 out_p.n1849 out_p.n1848 0.001
R35899 out_p.n1848 out_p.n1847 0.001
R35900 out_p.n1847 out_p.n1846 0.001
R35901 out_p.n1846 out_p.n1845 0.001
R35902 out_p.n1845 out_p.n1844 0.001
R35903 out_p.n1844 out_p.n1843 0.001
R35904 out_p.n1843 out_p.n1842 0.001
R35905 out_p.n1842 out_p.n1841 0.001
R35906 out_p.n1841 out_p.n1840 0.001
R35907 out_p.n1840 out_p.n1839 0.001
R35908 out_p.n1839 out_p.n1838 0.001
R35909 out_p.n1838 out_p.n1837 0.001
R35910 out_p.n1837 out_p.n1836 0.001
R35911 out_p.n1836 out_p.n1835 0.001
R35912 out_p.n1835 out_p.n1834 0.001
R35913 out_p.n1834 out_p.n1833 0.001
R35914 vdd.n13347 vdd.n13345 61.359
R35915 vdd.n13347 vdd.n13346 61.359
R35916 vdd.n13167 vdd.n13165 61.359
R35917 vdd.n13167 vdd.n13166 61.359
R35918 vdd.n12987 vdd.n12985 61.359
R35919 vdd.n12987 vdd.n12986 61.359
R35920 vdd.n12807 vdd.n12805 61.359
R35921 vdd.n12807 vdd.n12806 61.359
R35922 vdd.n12627 vdd.n12625 61.359
R35923 vdd.n12627 vdd.n12626 61.359
R35924 vdd.n12447 vdd.n12445 61.359
R35925 vdd.n12447 vdd.n12446 61.359
R35926 vdd.n12267 vdd.n12265 61.359
R35927 vdd.n12267 vdd.n12266 61.359
R35928 vdd.n12087 vdd.n12085 61.359
R35929 vdd.n12087 vdd.n12086 61.359
R35930 vdd.n11907 vdd.n11905 61.359
R35931 vdd.n11907 vdd.n11906 61.359
R35932 vdd.n11727 vdd.n11725 61.359
R35933 vdd.n11727 vdd.n11726 61.359
R35934 vdd.n11547 vdd.n11545 61.359
R35935 vdd.n11547 vdd.n11546 61.359
R35936 vdd.n68 vdd.n66 61.359
R35937 vdd.n68 vdd.n67 61.359
R35938 vdd.n248 vdd.n246 61.359
R35939 vdd.n248 vdd.n247 61.359
R35940 vdd.n428 vdd.n426 61.359
R35941 vdd.n428 vdd.n427 61.359
R35942 vdd.n608 vdd.n606 61.359
R35943 vdd.n608 vdd.n607 61.359
R35944 vdd.n788 vdd.n786 61.359
R35945 vdd.n788 vdd.n787 61.359
R35946 vdd.n968 vdd.n966 61.359
R35947 vdd.n968 vdd.n967 61.359
R35948 vdd.n1148 vdd.n1146 61.359
R35949 vdd.n1148 vdd.n1147 61.359
R35950 vdd.n1328 vdd.n1326 61.359
R35951 vdd.n1328 vdd.n1327 61.359
R35952 vdd.n1508 vdd.n1506 61.359
R35953 vdd.n1508 vdd.n1507 61.359
R35954 vdd.n1688 vdd.n1686 61.359
R35955 vdd.n1688 vdd.n1687 61.359
R35956 vdd.n1868 vdd.n1866 61.359
R35957 vdd.n1868 vdd.n1867 61.359
R35958 vdd.n2048 vdd.n2046 61.359
R35959 vdd.n2048 vdd.n2047 61.359
R35960 vdd.n2228 vdd.n2226 61.359
R35961 vdd.n2228 vdd.n2227 61.359
R35962 vdd.n2408 vdd.n2406 61.359
R35963 vdd.n2408 vdd.n2407 61.359
R35964 vdd.n2588 vdd.n2586 61.359
R35965 vdd.n2588 vdd.n2587 61.359
R35966 vdd.n2768 vdd.n2766 61.359
R35967 vdd.n2768 vdd.n2767 61.359
R35968 vdd.n2948 vdd.n2946 61.359
R35969 vdd.n2948 vdd.n2947 61.359
R35970 vdd.n3128 vdd.n3126 61.359
R35971 vdd.n3128 vdd.n3127 61.359
R35972 vdd.n3308 vdd.n3306 61.359
R35973 vdd.n3308 vdd.n3307 61.359
R35974 vdd.n3488 vdd.n3486 61.359
R35975 vdd.n3488 vdd.n3487 61.359
R35976 vdd.n3668 vdd.n3666 61.359
R35977 vdd.n3668 vdd.n3667 61.359
R35978 vdd.n3848 vdd.n3846 61.359
R35979 vdd.n3848 vdd.n3847 61.359
R35980 vdd.n4028 vdd.n4026 61.359
R35981 vdd.n4028 vdd.n4027 61.359
R35982 vdd.n4208 vdd.n4206 61.359
R35983 vdd.n4208 vdd.n4207 61.359
R35984 vdd.n4388 vdd.n4386 61.359
R35985 vdd.n4388 vdd.n4387 61.359
R35986 vdd.n4568 vdd.n4566 61.359
R35987 vdd.n4568 vdd.n4567 61.359
R35988 vdd.n4748 vdd.n4746 61.359
R35989 vdd.n4748 vdd.n4747 61.359
R35990 vdd.n4928 vdd.n4926 61.359
R35991 vdd.n4928 vdd.n4927 61.359
R35992 vdd.n5108 vdd.n5106 61.359
R35993 vdd.n5108 vdd.n5107 61.359
R35994 vdd.n5288 vdd.n5286 61.359
R35995 vdd.n5288 vdd.n5287 61.359
R35996 vdd.n5468 vdd.n5466 61.359
R35997 vdd.n5468 vdd.n5467 61.359
R35998 vdd.n5648 vdd.n5646 61.359
R35999 vdd.n5648 vdd.n5647 61.359
R36000 vdd.n5828 vdd.n5826 61.359
R36001 vdd.n5828 vdd.n5827 61.359
R36002 vdd.n6008 vdd.n6006 61.359
R36003 vdd.n6008 vdd.n6007 61.359
R36004 vdd.n6188 vdd.n6186 61.359
R36005 vdd.n6188 vdd.n6187 61.359
R36006 vdd.n6368 vdd.n6366 61.359
R36007 vdd.n6368 vdd.n6367 61.359
R36008 vdd.n6548 vdd.n6546 61.359
R36009 vdd.n6548 vdd.n6547 61.359
R36010 vdd.n6728 vdd.n6726 61.359
R36011 vdd.n6728 vdd.n6727 61.359
R36012 vdd.n6908 vdd.n6906 61.359
R36013 vdd.n6908 vdd.n6907 61.359
R36014 vdd.n7088 vdd.n7086 61.359
R36015 vdd.n7088 vdd.n7087 61.359
R36016 vdd.n7268 vdd.n7266 61.359
R36017 vdd.n7268 vdd.n7267 61.359
R36018 vdd.n7448 vdd.n7446 61.359
R36019 vdd.n7448 vdd.n7447 61.359
R36020 vdd.n7628 vdd.n7626 61.359
R36021 vdd.n7628 vdd.n7627 61.359
R36022 vdd.n7808 vdd.n7806 61.359
R36023 vdd.n7808 vdd.n7807 61.359
R36024 vdd.n7988 vdd.n7986 61.359
R36025 vdd.n7988 vdd.n7987 61.359
R36026 vdd.n8168 vdd.n8166 61.359
R36027 vdd.n8168 vdd.n8167 61.359
R36028 vdd.n8348 vdd.n8346 61.359
R36029 vdd.n8348 vdd.n8347 61.359
R36030 vdd.n8528 vdd.n8526 61.359
R36031 vdd.n8528 vdd.n8527 61.359
R36032 vdd.n8708 vdd.n8706 61.359
R36033 vdd.n8708 vdd.n8707 61.359
R36034 vdd.n8888 vdd.n8886 61.359
R36035 vdd.n8888 vdd.n8887 61.359
R36036 vdd.n9068 vdd.n9066 61.359
R36037 vdd.n9068 vdd.n9067 61.359
R36038 vdd.n9248 vdd.n9246 61.359
R36039 vdd.n9248 vdd.n9247 61.359
R36040 vdd.n9428 vdd.n9426 61.359
R36041 vdd.n9428 vdd.n9427 61.359
R36042 vdd.n9608 vdd.n9606 61.359
R36043 vdd.n9608 vdd.n9607 61.359
R36044 vdd.n9788 vdd.n9786 61.359
R36045 vdd.n9788 vdd.n9787 61.359
R36046 vdd.n9968 vdd.n9966 61.359
R36047 vdd.n9968 vdd.n9967 61.359
R36048 vdd.n10148 vdd.n10146 61.359
R36049 vdd.n10148 vdd.n10147 61.359
R36050 vdd.n10328 vdd.n10326 61.359
R36051 vdd.n10328 vdd.n10327 61.359
R36052 vdd.n10508 vdd.n10506 61.359
R36053 vdd.n10508 vdd.n10507 61.359
R36054 vdd.n10688 vdd.n10686 61.359
R36055 vdd.n10688 vdd.n10687 61.359
R36056 vdd.n10868 vdd.n10866 61.359
R36057 vdd.n10868 vdd.n10867 61.359
R36058 vdd.n11048 vdd.n11046 61.359
R36059 vdd.n11048 vdd.n11047 61.359
R36060 vdd.n11228 vdd.n11226 61.359
R36061 vdd.n11228 vdd.n11227 61.359
R36062 vdd.n13421 vdd.n13418 61.358
R36063 vdd.n13421 vdd.n13420 61.358
R36064 vdd.n13413 vdd.n13410 61.358
R36065 vdd.n13413 vdd.n13412 61.358
R36066 vdd.n13405 vdd.n13402 61.358
R36067 vdd.n13405 vdd.n13404 61.358
R36068 vdd.n13397 vdd.n13394 61.358
R36069 vdd.n13397 vdd.n13396 61.358
R36070 vdd.n13389 vdd.n13386 61.358
R36071 vdd.n13389 vdd.n13388 61.358
R36072 vdd.n13381 vdd.n13378 61.358
R36073 vdd.n13381 vdd.n13380 61.358
R36074 vdd.n13373 vdd.n13370 61.358
R36075 vdd.n13373 vdd.n13372 61.358
R36076 vdd.n13365 vdd.n13362 61.358
R36077 vdd.n13365 vdd.n13364 61.358
R36078 vdd.n13357 vdd.n13354 61.358
R36079 vdd.n13357 vdd.n13356 61.358
R36080 vdd.n13341 vdd.n13338 61.358
R36081 vdd.n13341 vdd.n13340 61.358
R36082 vdd.n13333 vdd.n13330 61.358
R36083 vdd.n13333 vdd.n13332 61.358
R36084 vdd.n13325 vdd.n13322 61.358
R36085 vdd.n13325 vdd.n13324 61.358
R36086 vdd.n13317 vdd.n13314 61.358
R36087 vdd.n13317 vdd.n13316 61.358
R36088 vdd.n13309 vdd.n13306 61.358
R36089 vdd.n13309 vdd.n13308 61.358
R36090 vdd.n13301 vdd.n13298 61.358
R36091 vdd.n13301 vdd.n13300 61.358
R36092 vdd.n13293 vdd.n13290 61.358
R36093 vdd.n13293 vdd.n13292 61.358
R36094 vdd.n13285 vdd.n13282 61.358
R36095 vdd.n13285 vdd.n13284 61.358
R36096 vdd.n13452 vdd.n13449 61.358
R36097 vdd.n13452 vdd.n13451 61.358
R36098 vdd.n13241 vdd.n13238 61.358
R36099 vdd.n13241 vdd.n13240 61.358
R36100 vdd.n13233 vdd.n13230 61.358
R36101 vdd.n13233 vdd.n13232 61.358
R36102 vdd.n13225 vdd.n13222 61.358
R36103 vdd.n13225 vdd.n13224 61.358
R36104 vdd.n13217 vdd.n13214 61.358
R36105 vdd.n13217 vdd.n13216 61.358
R36106 vdd.n13209 vdd.n13206 61.358
R36107 vdd.n13209 vdd.n13208 61.358
R36108 vdd.n13201 vdd.n13198 61.358
R36109 vdd.n13201 vdd.n13200 61.358
R36110 vdd.n13193 vdd.n13190 61.358
R36111 vdd.n13193 vdd.n13192 61.358
R36112 vdd.n13185 vdd.n13182 61.358
R36113 vdd.n13185 vdd.n13184 61.358
R36114 vdd.n13177 vdd.n13174 61.358
R36115 vdd.n13177 vdd.n13176 61.358
R36116 vdd.n13161 vdd.n13158 61.358
R36117 vdd.n13161 vdd.n13160 61.358
R36118 vdd.n13153 vdd.n13150 61.358
R36119 vdd.n13153 vdd.n13152 61.358
R36120 vdd.n13145 vdd.n13142 61.358
R36121 vdd.n13145 vdd.n13144 61.358
R36122 vdd.n13137 vdd.n13134 61.358
R36123 vdd.n13137 vdd.n13136 61.358
R36124 vdd.n13129 vdd.n13126 61.358
R36125 vdd.n13129 vdd.n13128 61.358
R36126 vdd.n13121 vdd.n13118 61.358
R36127 vdd.n13121 vdd.n13120 61.358
R36128 vdd.n13113 vdd.n13110 61.358
R36129 vdd.n13113 vdd.n13112 61.358
R36130 vdd.n13105 vdd.n13102 61.358
R36131 vdd.n13105 vdd.n13104 61.358
R36132 vdd.n13272 vdd.n13269 61.358
R36133 vdd.n13272 vdd.n13271 61.358
R36134 vdd.n13061 vdd.n13058 61.358
R36135 vdd.n13061 vdd.n13060 61.358
R36136 vdd.n13053 vdd.n13050 61.358
R36137 vdd.n13053 vdd.n13052 61.358
R36138 vdd.n13045 vdd.n13042 61.358
R36139 vdd.n13045 vdd.n13044 61.358
R36140 vdd.n13037 vdd.n13034 61.358
R36141 vdd.n13037 vdd.n13036 61.358
R36142 vdd.n13029 vdd.n13026 61.358
R36143 vdd.n13029 vdd.n13028 61.358
R36144 vdd.n13021 vdd.n13018 61.358
R36145 vdd.n13021 vdd.n13020 61.358
R36146 vdd.n13013 vdd.n13010 61.358
R36147 vdd.n13013 vdd.n13012 61.358
R36148 vdd.n13005 vdd.n13002 61.358
R36149 vdd.n13005 vdd.n13004 61.358
R36150 vdd.n12997 vdd.n12994 61.358
R36151 vdd.n12997 vdd.n12996 61.358
R36152 vdd.n12981 vdd.n12978 61.358
R36153 vdd.n12981 vdd.n12980 61.358
R36154 vdd.n12973 vdd.n12970 61.358
R36155 vdd.n12973 vdd.n12972 61.358
R36156 vdd.n12965 vdd.n12962 61.358
R36157 vdd.n12965 vdd.n12964 61.358
R36158 vdd.n12957 vdd.n12954 61.358
R36159 vdd.n12957 vdd.n12956 61.358
R36160 vdd.n12949 vdd.n12946 61.358
R36161 vdd.n12949 vdd.n12948 61.358
R36162 vdd.n12941 vdd.n12938 61.358
R36163 vdd.n12941 vdd.n12940 61.358
R36164 vdd.n12933 vdd.n12930 61.358
R36165 vdd.n12933 vdd.n12932 61.358
R36166 vdd.n12925 vdd.n12922 61.358
R36167 vdd.n12925 vdd.n12924 61.358
R36168 vdd.n13092 vdd.n13089 61.358
R36169 vdd.n13092 vdd.n13091 61.358
R36170 vdd.n12881 vdd.n12878 61.358
R36171 vdd.n12881 vdd.n12880 61.358
R36172 vdd.n12873 vdd.n12870 61.358
R36173 vdd.n12873 vdd.n12872 61.358
R36174 vdd.n12865 vdd.n12862 61.358
R36175 vdd.n12865 vdd.n12864 61.358
R36176 vdd.n12857 vdd.n12854 61.358
R36177 vdd.n12857 vdd.n12856 61.358
R36178 vdd.n12849 vdd.n12846 61.358
R36179 vdd.n12849 vdd.n12848 61.358
R36180 vdd.n12841 vdd.n12838 61.358
R36181 vdd.n12841 vdd.n12840 61.358
R36182 vdd.n12833 vdd.n12830 61.358
R36183 vdd.n12833 vdd.n12832 61.358
R36184 vdd.n12825 vdd.n12822 61.358
R36185 vdd.n12825 vdd.n12824 61.358
R36186 vdd.n12817 vdd.n12814 61.358
R36187 vdd.n12817 vdd.n12816 61.358
R36188 vdd.n12801 vdd.n12798 61.358
R36189 vdd.n12801 vdd.n12800 61.358
R36190 vdd.n12793 vdd.n12790 61.358
R36191 vdd.n12793 vdd.n12792 61.358
R36192 vdd.n12785 vdd.n12782 61.358
R36193 vdd.n12785 vdd.n12784 61.358
R36194 vdd.n12777 vdd.n12774 61.358
R36195 vdd.n12777 vdd.n12776 61.358
R36196 vdd.n12769 vdd.n12766 61.358
R36197 vdd.n12769 vdd.n12768 61.358
R36198 vdd.n12761 vdd.n12758 61.358
R36199 vdd.n12761 vdd.n12760 61.358
R36200 vdd.n12753 vdd.n12750 61.358
R36201 vdd.n12753 vdd.n12752 61.358
R36202 vdd.n12745 vdd.n12742 61.358
R36203 vdd.n12745 vdd.n12744 61.358
R36204 vdd.n12912 vdd.n12909 61.358
R36205 vdd.n12912 vdd.n12911 61.358
R36206 vdd.n12701 vdd.n12698 61.358
R36207 vdd.n12701 vdd.n12700 61.358
R36208 vdd.n12693 vdd.n12690 61.358
R36209 vdd.n12693 vdd.n12692 61.358
R36210 vdd.n12685 vdd.n12682 61.358
R36211 vdd.n12685 vdd.n12684 61.358
R36212 vdd.n12677 vdd.n12674 61.358
R36213 vdd.n12677 vdd.n12676 61.358
R36214 vdd.n12669 vdd.n12666 61.358
R36215 vdd.n12669 vdd.n12668 61.358
R36216 vdd.n12661 vdd.n12658 61.358
R36217 vdd.n12661 vdd.n12660 61.358
R36218 vdd.n12653 vdd.n12650 61.358
R36219 vdd.n12653 vdd.n12652 61.358
R36220 vdd.n12645 vdd.n12642 61.358
R36221 vdd.n12645 vdd.n12644 61.358
R36222 vdd.n12637 vdd.n12634 61.358
R36223 vdd.n12637 vdd.n12636 61.358
R36224 vdd.n12621 vdd.n12618 61.358
R36225 vdd.n12621 vdd.n12620 61.358
R36226 vdd.n12613 vdd.n12610 61.358
R36227 vdd.n12613 vdd.n12612 61.358
R36228 vdd.n12605 vdd.n12602 61.358
R36229 vdd.n12605 vdd.n12604 61.358
R36230 vdd.n12597 vdd.n12594 61.358
R36231 vdd.n12597 vdd.n12596 61.358
R36232 vdd.n12589 vdd.n12586 61.358
R36233 vdd.n12589 vdd.n12588 61.358
R36234 vdd.n12581 vdd.n12578 61.358
R36235 vdd.n12581 vdd.n12580 61.358
R36236 vdd.n12573 vdd.n12570 61.358
R36237 vdd.n12573 vdd.n12572 61.358
R36238 vdd.n12565 vdd.n12562 61.358
R36239 vdd.n12565 vdd.n12564 61.358
R36240 vdd.n12732 vdd.n12729 61.358
R36241 vdd.n12732 vdd.n12731 61.358
R36242 vdd.n12521 vdd.n12518 61.358
R36243 vdd.n12521 vdd.n12520 61.358
R36244 vdd.n12513 vdd.n12510 61.358
R36245 vdd.n12513 vdd.n12512 61.358
R36246 vdd.n12505 vdd.n12502 61.358
R36247 vdd.n12505 vdd.n12504 61.358
R36248 vdd.n12497 vdd.n12494 61.358
R36249 vdd.n12497 vdd.n12496 61.358
R36250 vdd.n12489 vdd.n12486 61.358
R36251 vdd.n12489 vdd.n12488 61.358
R36252 vdd.n12481 vdd.n12478 61.358
R36253 vdd.n12481 vdd.n12480 61.358
R36254 vdd.n12473 vdd.n12470 61.358
R36255 vdd.n12473 vdd.n12472 61.358
R36256 vdd.n12465 vdd.n12462 61.358
R36257 vdd.n12465 vdd.n12464 61.358
R36258 vdd.n12457 vdd.n12454 61.358
R36259 vdd.n12457 vdd.n12456 61.358
R36260 vdd.n12441 vdd.n12438 61.358
R36261 vdd.n12441 vdd.n12440 61.358
R36262 vdd.n12433 vdd.n12430 61.358
R36263 vdd.n12433 vdd.n12432 61.358
R36264 vdd.n12425 vdd.n12422 61.358
R36265 vdd.n12425 vdd.n12424 61.358
R36266 vdd.n12417 vdd.n12414 61.358
R36267 vdd.n12417 vdd.n12416 61.358
R36268 vdd.n12409 vdd.n12406 61.358
R36269 vdd.n12409 vdd.n12408 61.358
R36270 vdd.n12401 vdd.n12398 61.358
R36271 vdd.n12401 vdd.n12400 61.358
R36272 vdd.n12393 vdd.n12390 61.358
R36273 vdd.n12393 vdd.n12392 61.358
R36274 vdd.n12385 vdd.n12382 61.358
R36275 vdd.n12385 vdd.n12384 61.358
R36276 vdd.n12552 vdd.n12549 61.358
R36277 vdd.n12552 vdd.n12551 61.358
R36278 vdd.n12341 vdd.n12338 61.358
R36279 vdd.n12341 vdd.n12340 61.358
R36280 vdd.n12333 vdd.n12330 61.358
R36281 vdd.n12333 vdd.n12332 61.358
R36282 vdd.n12325 vdd.n12322 61.358
R36283 vdd.n12325 vdd.n12324 61.358
R36284 vdd.n12317 vdd.n12314 61.358
R36285 vdd.n12317 vdd.n12316 61.358
R36286 vdd.n12309 vdd.n12306 61.358
R36287 vdd.n12309 vdd.n12308 61.358
R36288 vdd.n12301 vdd.n12298 61.358
R36289 vdd.n12301 vdd.n12300 61.358
R36290 vdd.n12293 vdd.n12290 61.358
R36291 vdd.n12293 vdd.n12292 61.358
R36292 vdd.n12285 vdd.n12282 61.358
R36293 vdd.n12285 vdd.n12284 61.358
R36294 vdd.n12277 vdd.n12274 61.358
R36295 vdd.n12277 vdd.n12276 61.358
R36296 vdd.n12261 vdd.n12258 61.358
R36297 vdd.n12261 vdd.n12260 61.358
R36298 vdd.n12253 vdd.n12250 61.358
R36299 vdd.n12253 vdd.n12252 61.358
R36300 vdd.n12245 vdd.n12242 61.358
R36301 vdd.n12245 vdd.n12244 61.358
R36302 vdd.n12237 vdd.n12234 61.358
R36303 vdd.n12237 vdd.n12236 61.358
R36304 vdd.n12229 vdd.n12226 61.358
R36305 vdd.n12229 vdd.n12228 61.358
R36306 vdd.n12221 vdd.n12218 61.358
R36307 vdd.n12221 vdd.n12220 61.358
R36308 vdd.n12213 vdd.n12210 61.358
R36309 vdd.n12213 vdd.n12212 61.358
R36310 vdd.n12205 vdd.n12202 61.358
R36311 vdd.n12205 vdd.n12204 61.358
R36312 vdd.n12372 vdd.n12369 61.358
R36313 vdd.n12372 vdd.n12371 61.358
R36314 vdd.n12161 vdd.n12158 61.358
R36315 vdd.n12161 vdd.n12160 61.358
R36316 vdd.n12153 vdd.n12150 61.358
R36317 vdd.n12153 vdd.n12152 61.358
R36318 vdd.n12145 vdd.n12142 61.358
R36319 vdd.n12145 vdd.n12144 61.358
R36320 vdd.n12137 vdd.n12134 61.358
R36321 vdd.n12137 vdd.n12136 61.358
R36322 vdd.n12129 vdd.n12126 61.358
R36323 vdd.n12129 vdd.n12128 61.358
R36324 vdd.n12121 vdd.n12118 61.358
R36325 vdd.n12121 vdd.n12120 61.358
R36326 vdd.n12113 vdd.n12110 61.358
R36327 vdd.n12113 vdd.n12112 61.358
R36328 vdd.n12105 vdd.n12102 61.358
R36329 vdd.n12105 vdd.n12104 61.358
R36330 vdd.n12097 vdd.n12094 61.358
R36331 vdd.n12097 vdd.n12096 61.358
R36332 vdd.n12081 vdd.n12078 61.358
R36333 vdd.n12081 vdd.n12080 61.358
R36334 vdd.n12073 vdd.n12070 61.358
R36335 vdd.n12073 vdd.n12072 61.358
R36336 vdd.n12065 vdd.n12062 61.358
R36337 vdd.n12065 vdd.n12064 61.358
R36338 vdd.n12057 vdd.n12054 61.358
R36339 vdd.n12057 vdd.n12056 61.358
R36340 vdd.n12049 vdd.n12046 61.358
R36341 vdd.n12049 vdd.n12048 61.358
R36342 vdd.n12041 vdd.n12038 61.358
R36343 vdd.n12041 vdd.n12040 61.358
R36344 vdd.n12033 vdd.n12030 61.358
R36345 vdd.n12033 vdd.n12032 61.358
R36346 vdd.n12025 vdd.n12022 61.358
R36347 vdd.n12025 vdd.n12024 61.358
R36348 vdd.n12192 vdd.n12189 61.358
R36349 vdd.n12192 vdd.n12191 61.358
R36350 vdd.n11981 vdd.n11978 61.358
R36351 vdd.n11981 vdd.n11980 61.358
R36352 vdd.n11973 vdd.n11970 61.358
R36353 vdd.n11973 vdd.n11972 61.358
R36354 vdd.n11965 vdd.n11962 61.358
R36355 vdd.n11965 vdd.n11964 61.358
R36356 vdd.n11957 vdd.n11954 61.358
R36357 vdd.n11957 vdd.n11956 61.358
R36358 vdd.n11949 vdd.n11946 61.358
R36359 vdd.n11949 vdd.n11948 61.358
R36360 vdd.n11941 vdd.n11938 61.358
R36361 vdd.n11941 vdd.n11940 61.358
R36362 vdd.n11933 vdd.n11930 61.358
R36363 vdd.n11933 vdd.n11932 61.358
R36364 vdd.n11925 vdd.n11922 61.358
R36365 vdd.n11925 vdd.n11924 61.358
R36366 vdd.n11917 vdd.n11914 61.358
R36367 vdd.n11917 vdd.n11916 61.358
R36368 vdd.n11901 vdd.n11898 61.358
R36369 vdd.n11901 vdd.n11900 61.358
R36370 vdd.n11893 vdd.n11890 61.358
R36371 vdd.n11893 vdd.n11892 61.358
R36372 vdd.n11885 vdd.n11882 61.358
R36373 vdd.n11885 vdd.n11884 61.358
R36374 vdd.n11877 vdd.n11874 61.358
R36375 vdd.n11877 vdd.n11876 61.358
R36376 vdd.n11869 vdd.n11866 61.358
R36377 vdd.n11869 vdd.n11868 61.358
R36378 vdd.n11861 vdd.n11858 61.358
R36379 vdd.n11861 vdd.n11860 61.358
R36380 vdd.n11853 vdd.n11850 61.358
R36381 vdd.n11853 vdd.n11852 61.358
R36382 vdd.n11845 vdd.n11842 61.358
R36383 vdd.n11845 vdd.n11844 61.358
R36384 vdd.n12012 vdd.n12009 61.358
R36385 vdd.n12012 vdd.n12011 61.358
R36386 vdd.n11801 vdd.n11798 61.358
R36387 vdd.n11801 vdd.n11800 61.358
R36388 vdd.n11793 vdd.n11790 61.358
R36389 vdd.n11793 vdd.n11792 61.358
R36390 vdd.n11785 vdd.n11782 61.358
R36391 vdd.n11785 vdd.n11784 61.358
R36392 vdd.n11777 vdd.n11774 61.358
R36393 vdd.n11777 vdd.n11776 61.358
R36394 vdd.n11769 vdd.n11766 61.358
R36395 vdd.n11769 vdd.n11768 61.358
R36396 vdd.n11761 vdd.n11758 61.358
R36397 vdd.n11761 vdd.n11760 61.358
R36398 vdd.n11753 vdd.n11750 61.358
R36399 vdd.n11753 vdd.n11752 61.358
R36400 vdd.n11745 vdd.n11742 61.358
R36401 vdd.n11745 vdd.n11744 61.358
R36402 vdd.n11737 vdd.n11734 61.358
R36403 vdd.n11737 vdd.n11736 61.358
R36404 vdd.n11721 vdd.n11718 61.358
R36405 vdd.n11721 vdd.n11720 61.358
R36406 vdd.n11713 vdd.n11710 61.358
R36407 vdd.n11713 vdd.n11712 61.358
R36408 vdd.n11705 vdd.n11702 61.358
R36409 vdd.n11705 vdd.n11704 61.358
R36410 vdd.n11697 vdd.n11694 61.358
R36411 vdd.n11697 vdd.n11696 61.358
R36412 vdd.n11689 vdd.n11686 61.358
R36413 vdd.n11689 vdd.n11688 61.358
R36414 vdd.n11681 vdd.n11678 61.358
R36415 vdd.n11681 vdd.n11680 61.358
R36416 vdd.n11673 vdd.n11670 61.358
R36417 vdd.n11673 vdd.n11672 61.358
R36418 vdd.n11665 vdd.n11662 61.358
R36419 vdd.n11665 vdd.n11664 61.358
R36420 vdd.n11832 vdd.n11829 61.358
R36421 vdd.n11832 vdd.n11831 61.358
R36422 vdd.n11621 vdd.n11618 61.358
R36423 vdd.n11621 vdd.n11620 61.358
R36424 vdd.n11613 vdd.n11610 61.358
R36425 vdd.n11613 vdd.n11612 61.358
R36426 vdd.n11605 vdd.n11602 61.358
R36427 vdd.n11605 vdd.n11604 61.358
R36428 vdd.n11597 vdd.n11594 61.358
R36429 vdd.n11597 vdd.n11596 61.358
R36430 vdd.n11589 vdd.n11586 61.358
R36431 vdd.n11589 vdd.n11588 61.358
R36432 vdd.n11581 vdd.n11578 61.358
R36433 vdd.n11581 vdd.n11580 61.358
R36434 vdd.n11573 vdd.n11570 61.358
R36435 vdd.n11573 vdd.n11572 61.358
R36436 vdd.n11565 vdd.n11562 61.358
R36437 vdd.n11565 vdd.n11564 61.358
R36438 vdd.n11557 vdd.n11554 61.358
R36439 vdd.n11557 vdd.n11556 61.358
R36440 vdd.n11541 vdd.n11538 61.358
R36441 vdd.n11541 vdd.n11540 61.358
R36442 vdd.n11533 vdd.n11530 61.358
R36443 vdd.n11533 vdd.n11532 61.358
R36444 vdd.n11525 vdd.n11522 61.358
R36445 vdd.n11525 vdd.n11524 61.358
R36446 vdd.n11517 vdd.n11514 61.358
R36447 vdd.n11517 vdd.n11516 61.358
R36448 vdd.n11509 vdd.n11506 61.358
R36449 vdd.n11509 vdd.n11508 61.358
R36450 vdd.n11501 vdd.n11498 61.358
R36451 vdd.n11501 vdd.n11500 61.358
R36452 vdd.n11493 vdd.n11490 61.358
R36453 vdd.n11493 vdd.n11492 61.358
R36454 vdd.n11485 vdd.n11482 61.358
R36455 vdd.n11485 vdd.n11484 61.358
R36456 vdd.n11652 vdd.n11649 61.358
R36457 vdd.n11652 vdd.n11651 61.358
R36458 vdd.n142 vdd.n139 61.358
R36459 vdd.n142 vdd.n141 61.358
R36460 vdd.n134 vdd.n131 61.358
R36461 vdd.n134 vdd.n133 61.358
R36462 vdd.n126 vdd.n123 61.358
R36463 vdd.n126 vdd.n125 61.358
R36464 vdd.n118 vdd.n115 61.358
R36465 vdd.n118 vdd.n117 61.358
R36466 vdd.n110 vdd.n107 61.358
R36467 vdd.n110 vdd.n109 61.358
R36468 vdd.n102 vdd.n99 61.358
R36469 vdd.n102 vdd.n101 61.358
R36470 vdd.n94 vdd.n91 61.358
R36471 vdd.n94 vdd.n93 61.358
R36472 vdd.n86 vdd.n83 61.358
R36473 vdd.n86 vdd.n85 61.358
R36474 vdd.n78 vdd.n75 61.358
R36475 vdd.n78 vdd.n77 61.358
R36476 vdd.n62 vdd.n59 61.358
R36477 vdd.n62 vdd.n61 61.358
R36478 vdd.n54 vdd.n51 61.358
R36479 vdd.n54 vdd.n53 61.358
R36480 vdd.n46 vdd.n43 61.358
R36481 vdd.n46 vdd.n45 61.358
R36482 vdd.n38 vdd.n35 61.358
R36483 vdd.n38 vdd.n37 61.358
R36484 vdd.n30 vdd.n27 61.358
R36485 vdd.n30 vdd.n29 61.358
R36486 vdd.n22 vdd.n19 61.358
R36487 vdd.n22 vdd.n21 61.358
R36488 vdd.n14 vdd.n11 61.358
R36489 vdd.n14 vdd.n13 61.358
R36490 vdd.n6 vdd.n3 61.358
R36491 vdd.n6 vdd.n5 61.358
R36492 vdd.n173 vdd.n170 61.358
R36493 vdd.n173 vdd.n172 61.358
R36494 vdd.n322 vdd.n319 61.358
R36495 vdd.n322 vdd.n321 61.358
R36496 vdd.n314 vdd.n311 61.358
R36497 vdd.n314 vdd.n313 61.358
R36498 vdd.n306 vdd.n303 61.358
R36499 vdd.n306 vdd.n305 61.358
R36500 vdd.n298 vdd.n295 61.358
R36501 vdd.n298 vdd.n297 61.358
R36502 vdd.n290 vdd.n287 61.358
R36503 vdd.n290 vdd.n289 61.358
R36504 vdd.n282 vdd.n279 61.358
R36505 vdd.n282 vdd.n281 61.358
R36506 vdd.n274 vdd.n271 61.358
R36507 vdd.n274 vdd.n273 61.358
R36508 vdd.n266 vdd.n263 61.358
R36509 vdd.n266 vdd.n265 61.358
R36510 vdd.n258 vdd.n255 61.358
R36511 vdd.n258 vdd.n257 61.358
R36512 vdd.n242 vdd.n239 61.358
R36513 vdd.n242 vdd.n241 61.358
R36514 vdd.n234 vdd.n231 61.358
R36515 vdd.n234 vdd.n233 61.358
R36516 vdd.n226 vdd.n223 61.358
R36517 vdd.n226 vdd.n225 61.358
R36518 vdd.n218 vdd.n215 61.358
R36519 vdd.n218 vdd.n217 61.358
R36520 vdd.n210 vdd.n207 61.358
R36521 vdd.n210 vdd.n209 61.358
R36522 vdd.n202 vdd.n199 61.358
R36523 vdd.n202 vdd.n201 61.358
R36524 vdd.n194 vdd.n191 61.358
R36525 vdd.n194 vdd.n193 61.358
R36526 vdd.n186 vdd.n183 61.358
R36527 vdd.n186 vdd.n185 61.358
R36528 vdd.n353 vdd.n350 61.358
R36529 vdd.n353 vdd.n352 61.358
R36530 vdd.n502 vdd.n499 61.358
R36531 vdd.n502 vdd.n501 61.358
R36532 vdd.n494 vdd.n491 61.358
R36533 vdd.n494 vdd.n493 61.358
R36534 vdd.n486 vdd.n483 61.358
R36535 vdd.n486 vdd.n485 61.358
R36536 vdd.n478 vdd.n475 61.358
R36537 vdd.n478 vdd.n477 61.358
R36538 vdd.n470 vdd.n467 61.358
R36539 vdd.n470 vdd.n469 61.358
R36540 vdd.n462 vdd.n459 61.358
R36541 vdd.n462 vdd.n461 61.358
R36542 vdd.n454 vdd.n451 61.358
R36543 vdd.n454 vdd.n453 61.358
R36544 vdd.n446 vdd.n443 61.358
R36545 vdd.n446 vdd.n445 61.358
R36546 vdd.n438 vdd.n435 61.358
R36547 vdd.n438 vdd.n437 61.358
R36548 vdd.n422 vdd.n419 61.358
R36549 vdd.n422 vdd.n421 61.358
R36550 vdd.n414 vdd.n411 61.358
R36551 vdd.n414 vdd.n413 61.358
R36552 vdd.n406 vdd.n403 61.358
R36553 vdd.n406 vdd.n405 61.358
R36554 vdd.n398 vdd.n395 61.358
R36555 vdd.n398 vdd.n397 61.358
R36556 vdd.n390 vdd.n387 61.358
R36557 vdd.n390 vdd.n389 61.358
R36558 vdd.n382 vdd.n379 61.358
R36559 vdd.n382 vdd.n381 61.358
R36560 vdd.n374 vdd.n371 61.358
R36561 vdd.n374 vdd.n373 61.358
R36562 vdd.n366 vdd.n363 61.358
R36563 vdd.n366 vdd.n365 61.358
R36564 vdd.n533 vdd.n530 61.358
R36565 vdd.n533 vdd.n532 61.358
R36566 vdd.n682 vdd.n679 61.358
R36567 vdd.n682 vdd.n681 61.358
R36568 vdd.n674 vdd.n671 61.358
R36569 vdd.n674 vdd.n673 61.358
R36570 vdd.n666 vdd.n663 61.358
R36571 vdd.n666 vdd.n665 61.358
R36572 vdd.n658 vdd.n655 61.358
R36573 vdd.n658 vdd.n657 61.358
R36574 vdd.n650 vdd.n647 61.358
R36575 vdd.n650 vdd.n649 61.358
R36576 vdd.n642 vdd.n639 61.358
R36577 vdd.n642 vdd.n641 61.358
R36578 vdd.n634 vdd.n631 61.358
R36579 vdd.n634 vdd.n633 61.358
R36580 vdd.n626 vdd.n623 61.358
R36581 vdd.n626 vdd.n625 61.358
R36582 vdd.n618 vdd.n615 61.358
R36583 vdd.n618 vdd.n617 61.358
R36584 vdd.n602 vdd.n599 61.358
R36585 vdd.n602 vdd.n601 61.358
R36586 vdd.n594 vdd.n591 61.358
R36587 vdd.n594 vdd.n593 61.358
R36588 vdd.n586 vdd.n583 61.358
R36589 vdd.n586 vdd.n585 61.358
R36590 vdd.n578 vdd.n575 61.358
R36591 vdd.n578 vdd.n577 61.358
R36592 vdd.n570 vdd.n567 61.358
R36593 vdd.n570 vdd.n569 61.358
R36594 vdd.n562 vdd.n559 61.358
R36595 vdd.n562 vdd.n561 61.358
R36596 vdd.n554 vdd.n551 61.358
R36597 vdd.n554 vdd.n553 61.358
R36598 vdd.n546 vdd.n543 61.358
R36599 vdd.n546 vdd.n545 61.358
R36600 vdd.n713 vdd.n710 61.358
R36601 vdd.n713 vdd.n712 61.358
R36602 vdd.n862 vdd.n859 61.358
R36603 vdd.n862 vdd.n861 61.358
R36604 vdd.n854 vdd.n851 61.358
R36605 vdd.n854 vdd.n853 61.358
R36606 vdd.n846 vdd.n843 61.358
R36607 vdd.n846 vdd.n845 61.358
R36608 vdd.n838 vdd.n835 61.358
R36609 vdd.n838 vdd.n837 61.358
R36610 vdd.n830 vdd.n827 61.358
R36611 vdd.n830 vdd.n829 61.358
R36612 vdd.n822 vdd.n819 61.358
R36613 vdd.n822 vdd.n821 61.358
R36614 vdd.n814 vdd.n811 61.358
R36615 vdd.n814 vdd.n813 61.358
R36616 vdd.n806 vdd.n803 61.358
R36617 vdd.n806 vdd.n805 61.358
R36618 vdd.n798 vdd.n795 61.358
R36619 vdd.n798 vdd.n797 61.358
R36620 vdd.n782 vdd.n779 61.358
R36621 vdd.n782 vdd.n781 61.358
R36622 vdd.n774 vdd.n771 61.358
R36623 vdd.n774 vdd.n773 61.358
R36624 vdd.n766 vdd.n763 61.358
R36625 vdd.n766 vdd.n765 61.358
R36626 vdd.n758 vdd.n755 61.358
R36627 vdd.n758 vdd.n757 61.358
R36628 vdd.n750 vdd.n747 61.358
R36629 vdd.n750 vdd.n749 61.358
R36630 vdd.n742 vdd.n739 61.358
R36631 vdd.n742 vdd.n741 61.358
R36632 vdd.n734 vdd.n731 61.358
R36633 vdd.n734 vdd.n733 61.358
R36634 vdd.n726 vdd.n723 61.358
R36635 vdd.n726 vdd.n725 61.358
R36636 vdd.n893 vdd.n890 61.358
R36637 vdd.n893 vdd.n892 61.358
R36638 vdd.n1042 vdd.n1039 61.358
R36639 vdd.n1042 vdd.n1041 61.358
R36640 vdd.n1034 vdd.n1031 61.358
R36641 vdd.n1034 vdd.n1033 61.358
R36642 vdd.n1026 vdd.n1023 61.358
R36643 vdd.n1026 vdd.n1025 61.358
R36644 vdd.n1018 vdd.n1015 61.358
R36645 vdd.n1018 vdd.n1017 61.358
R36646 vdd.n1010 vdd.n1007 61.358
R36647 vdd.n1010 vdd.n1009 61.358
R36648 vdd.n1002 vdd.n999 61.358
R36649 vdd.n1002 vdd.n1001 61.358
R36650 vdd.n994 vdd.n991 61.358
R36651 vdd.n994 vdd.n993 61.358
R36652 vdd.n986 vdd.n983 61.358
R36653 vdd.n986 vdd.n985 61.358
R36654 vdd.n978 vdd.n975 61.358
R36655 vdd.n978 vdd.n977 61.358
R36656 vdd.n962 vdd.n959 61.358
R36657 vdd.n962 vdd.n961 61.358
R36658 vdd.n954 vdd.n951 61.358
R36659 vdd.n954 vdd.n953 61.358
R36660 vdd.n946 vdd.n943 61.358
R36661 vdd.n946 vdd.n945 61.358
R36662 vdd.n938 vdd.n935 61.358
R36663 vdd.n938 vdd.n937 61.358
R36664 vdd.n930 vdd.n927 61.358
R36665 vdd.n930 vdd.n929 61.358
R36666 vdd.n922 vdd.n919 61.358
R36667 vdd.n922 vdd.n921 61.358
R36668 vdd.n914 vdd.n911 61.358
R36669 vdd.n914 vdd.n913 61.358
R36670 vdd.n906 vdd.n903 61.358
R36671 vdd.n906 vdd.n905 61.358
R36672 vdd.n1073 vdd.n1070 61.358
R36673 vdd.n1073 vdd.n1072 61.358
R36674 vdd.n1222 vdd.n1219 61.358
R36675 vdd.n1222 vdd.n1221 61.358
R36676 vdd.n1214 vdd.n1211 61.358
R36677 vdd.n1214 vdd.n1213 61.358
R36678 vdd.n1206 vdd.n1203 61.358
R36679 vdd.n1206 vdd.n1205 61.358
R36680 vdd.n1198 vdd.n1195 61.358
R36681 vdd.n1198 vdd.n1197 61.358
R36682 vdd.n1190 vdd.n1187 61.358
R36683 vdd.n1190 vdd.n1189 61.358
R36684 vdd.n1182 vdd.n1179 61.358
R36685 vdd.n1182 vdd.n1181 61.358
R36686 vdd.n1174 vdd.n1171 61.358
R36687 vdd.n1174 vdd.n1173 61.358
R36688 vdd.n1166 vdd.n1163 61.358
R36689 vdd.n1166 vdd.n1165 61.358
R36690 vdd.n1158 vdd.n1155 61.358
R36691 vdd.n1158 vdd.n1157 61.358
R36692 vdd.n1142 vdd.n1139 61.358
R36693 vdd.n1142 vdd.n1141 61.358
R36694 vdd.n1134 vdd.n1131 61.358
R36695 vdd.n1134 vdd.n1133 61.358
R36696 vdd.n1126 vdd.n1123 61.358
R36697 vdd.n1126 vdd.n1125 61.358
R36698 vdd.n1118 vdd.n1115 61.358
R36699 vdd.n1118 vdd.n1117 61.358
R36700 vdd.n1110 vdd.n1107 61.358
R36701 vdd.n1110 vdd.n1109 61.358
R36702 vdd.n1102 vdd.n1099 61.358
R36703 vdd.n1102 vdd.n1101 61.358
R36704 vdd.n1094 vdd.n1091 61.358
R36705 vdd.n1094 vdd.n1093 61.358
R36706 vdd.n1086 vdd.n1083 61.358
R36707 vdd.n1086 vdd.n1085 61.358
R36708 vdd.n1253 vdd.n1250 61.358
R36709 vdd.n1253 vdd.n1252 61.358
R36710 vdd.n1402 vdd.n1399 61.358
R36711 vdd.n1402 vdd.n1401 61.358
R36712 vdd.n1394 vdd.n1391 61.358
R36713 vdd.n1394 vdd.n1393 61.358
R36714 vdd.n1386 vdd.n1383 61.358
R36715 vdd.n1386 vdd.n1385 61.358
R36716 vdd.n1378 vdd.n1375 61.358
R36717 vdd.n1378 vdd.n1377 61.358
R36718 vdd.n1370 vdd.n1367 61.358
R36719 vdd.n1370 vdd.n1369 61.358
R36720 vdd.n1362 vdd.n1359 61.358
R36721 vdd.n1362 vdd.n1361 61.358
R36722 vdd.n1354 vdd.n1351 61.358
R36723 vdd.n1354 vdd.n1353 61.358
R36724 vdd.n1346 vdd.n1343 61.358
R36725 vdd.n1346 vdd.n1345 61.358
R36726 vdd.n1338 vdd.n1335 61.358
R36727 vdd.n1338 vdd.n1337 61.358
R36728 vdd.n1322 vdd.n1319 61.358
R36729 vdd.n1322 vdd.n1321 61.358
R36730 vdd.n1314 vdd.n1311 61.358
R36731 vdd.n1314 vdd.n1313 61.358
R36732 vdd.n1306 vdd.n1303 61.358
R36733 vdd.n1306 vdd.n1305 61.358
R36734 vdd.n1298 vdd.n1295 61.358
R36735 vdd.n1298 vdd.n1297 61.358
R36736 vdd.n1290 vdd.n1287 61.358
R36737 vdd.n1290 vdd.n1289 61.358
R36738 vdd.n1282 vdd.n1279 61.358
R36739 vdd.n1282 vdd.n1281 61.358
R36740 vdd.n1274 vdd.n1271 61.358
R36741 vdd.n1274 vdd.n1273 61.358
R36742 vdd.n1266 vdd.n1263 61.358
R36743 vdd.n1266 vdd.n1265 61.358
R36744 vdd.n1433 vdd.n1430 61.358
R36745 vdd.n1433 vdd.n1432 61.358
R36746 vdd.n1582 vdd.n1579 61.358
R36747 vdd.n1582 vdd.n1581 61.358
R36748 vdd.n1574 vdd.n1571 61.358
R36749 vdd.n1574 vdd.n1573 61.358
R36750 vdd.n1566 vdd.n1563 61.358
R36751 vdd.n1566 vdd.n1565 61.358
R36752 vdd.n1558 vdd.n1555 61.358
R36753 vdd.n1558 vdd.n1557 61.358
R36754 vdd.n1550 vdd.n1547 61.358
R36755 vdd.n1550 vdd.n1549 61.358
R36756 vdd.n1542 vdd.n1539 61.358
R36757 vdd.n1542 vdd.n1541 61.358
R36758 vdd.n1534 vdd.n1531 61.358
R36759 vdd.n1534 vdd.n1533 61.358
R36760 vdd.n1526 vdd.n1523 61.358
R36761 vdd.n1526 vdd.n1525 61.358
R36762 vdd.n1518 vdd.n1515 61.358
R36763 vdd.n1518 vdd.n1517 61.358
R36764 vdd.n1502 vdd.n1499 61.358
R36765 vdd.n1502 vdd.n1501 61.358
R36766 vdd.n1494 vdd.n1491 61.358
R36767 vdd.n1494 vdd.n1493 61.358
R36768 vdd.n1486 vdd.n1483 61.358
R36769 vdd.n1486 vdd.n1485 61.358
R36770 vdd.n1478 vdd.n1475 61.358
R36771 vdd.n1478 vdd.n1477 61.358
R36772 vdd.n1470 vdd.n1467 61.358
R36773 vdd.n1470 vdd.n1469 61.358
R36774 vdd.n1462 vdd.n1459 61.358
R36775 vdd.n1462 vdd.n1461 61.358
R36776 vdd.n1454 vdd.n1451 61.358
R36777 vdd.n1454 vdd.n1453 61.358
R36778 vdd.n1446 vdd.n1443 61.358
R36779 vdd.n1446 vdd.n1445 61.358
R36780 vdd.n1613 vdd.n1610 61.358
R36781 vdd.n1613 vdd.n1612 61.358
R36782 vdd.n1762 vdd.n1759 61.358
R36783 vdd.n1762 vdd.n1761 61.358
R36784 vdd.n1754 vdd.n1751 61.358
R36785 vdd.n1754 vdd.n1753 61.358
R36786 vdd.n1746 vdd.n1743 61.358
R36787 vdd.n1746 vdd.n1745 61.358
R36788 vdd.n1738 vdd.n1735 61.358
R36789 vdd.n1738 vdd.n1737 61.358
R36790 vdd.n1730 vdd.n1727 61.358
R36791 vdd.n1730 vdd.n1729 61.358
R36792 vdd.n1722 vdd.n1719 61.358
R36793 vdd.n1722 vdd.n1721 61.358
R36794 vdd.n1714 vdd.n1711 61.358
R36795 vdd.n1714 vdd.n1713 61.358
R36796 vdd.n1706 vdd.n1703 61.358
R36797 vdd.n1706 vdd.n1705 61.358
R36798 vdd.n1698 vdd.n1695 61.358
R36799 vdd.n1698 vdd.n1697 61.358
R36800 vdd.n1682 vdd.n1679 61.358
R36801 vdd.n1682 vdd.n1681 61.358
R36802 vdd.n1674 vdd.n1671 61.358
R36803 vdd.n1674 vdd.n1673 61.358
R36804 vdd.n1666 vdd.n1663 61.358
R36805 vdd.n1666 vdd.n1665 61.358
R36806 vdd.n1658 vdd.n1655 61.358
R36807 vdd.n1658 vdd.n1657 61.358
R36808 vdd.n1650 vdd.n1647 61.358
R36809 vdd.n1650 vdd.n1649 61.358
R36810 vdd.n1642 vdd.n1639 61.358
R36811 vdd.n1642 vdd.n1641 61.358
R36812 vdd.n1634 vdd.n1631 61.358
R36813 vdd.n1634 vdd.n1633 61.358
R36814 vdd.n1626 vdd.n1623 61.358
R36815 vdd.n1626 vdd.n1625 61.358
R36816 vdd.n1793 vdd.n1790 61.358
R36817 vdd.n1793 vdd.n1792 61.358
R36818 vdd.n1942 vdd.n1939 61.358
R36819 vdd.n1942 vdd.n1941 61.358
R36820 vdd.n1934 vdd.n1931 61.358
R36821 vdd.n1934 vdd.n1933 61.358
R36822 vdd.n1926 vdd.n1923 61.358
R36823 vdd.n1926 vdd.n1925 61.358
R36824 vdd.n1918 vdd.n1915 61.358
R36825 vdd.n1918 vdd.n1917 61.358
R36826 vdd.n1910 vdd.n1907 61.358
R36827 vdd.n1910 vdd.n1909 61.358
R36828 vdd.n1902 vdd.n1899 61.358
R36829 vdd.n1902 vdd.n1901 61.358
R36830 vdd.n1894 vdd.n1891 61.358
R36831 vdd.n1894 vdd.n1893 61.358
R36832 vdd.n1886 vdd.n1883 61.358
R36833 vdd.n1886 vdd.n1885 61.358
R36834 vdd.n1878 vdd.n1875 61.358
R36835 vdd.n1878 vdd.n1877 61.358
R36836 vdd.n1862 vdd.n1859 61.358
R36837 vdd.n1862 vdd.n1861 61.358
R36838 vdd.n1854 vdd.n1851 61.358
R36839 vdd.n1854 vdd.n1853 61.358
R36840 vdd.n1846 vdd.n1843 61.358
R36841 vdd.n1846 vdd.n1845 61.358
R36842 vdd.n1838 vdd.n1835 61.358
R36843 vdd.n1838 vdd.n1837 61.358
R36844 vdd.n1830 vdd.n1827 61.358
R36845 vdd.n1830 vdd.n1829 61.358
R36846 vdd.n1822 vdd.n1819 61.358
R36847 vdd.n1822 vdd.n1821 61.358
R36848 vdd.n1814 vdd.n1811 61.358
R36849 vdd.n1814 vdd.n1813 61.358
R36850 vdd.n1806 vdd.n1803 61.358
R36851 vdd.n1806 vdd.n1805 61.358
R36852 vdd.n1973 vdd.n1970 61.358
R36853 vdd.n1973 vdd.n1972 61.358
R36854 vdd.n2122 vdd.n2119 61.358
R36855 vdd.n2122 vdd.n2121 61.358
R36856 vdd.n2114 vdd.n2111 61.358
R36857 vdd.n2114 vdd.n2113 61.358
R36858 vdd.n2106 vdd.n2103 61.358
R36859 vdd.n2106 vdd.n2105 61.358
R36860 vdd.n2098 vdd.n2095 61.358
R36861 vdd.n2098 vdd.n2097 61.358
R36862 vdd.n2090 vdd.n2087 61.358
R36863 vdd.n2090 vdd.n2089 61.358
R36864 vdd.n2082 vdd.n2079 61.358
R36865 vdd.n2082 vdd.n2081 61.358
R36866 vdd.n2074 vdd.n2071 61.358
R36867 vdd.n2074 vdd.n2073 61.358
R36868 vdd.n2066 vdd.n2063 61.358
R36869 vdd.n2066 vdd.n2065 61.358
R36870 vdd.n2058 vdd.n2055 61.358
R36871 vdd.n2058 vdd.n2057 61.358
R36872 vdd.n2042 vdd.n2039 61.358
R36873 vdd.n2042 vdd.n2041 61.358
R36874 vdd.n2034 vdd.n2031 61.358
R36875 vdd.n2034 vdd.n2033 61.358
R36876 vdd.n2026 vdd.n2023 61.358
R36877 vdd.n2026 vdd.n2025 61.358
R36878 vdd.n2018 vdd.n2015 61.358
R36879 vdd.n2018 vdd.n2017 61.358
R36880 vdd.n2010 vdd.n2007 61.358
R36881 vdd.n2010 vdd.n2009 61.358
R36882 vdd.n2002 vdd.n1999 61.358
R36883 vdd.n2002 vdd.n2001 61.358
R36884 vdd.n1994 vdd.n1991 61.358
R36885 vdd.n1994 vdd.n1993 61.358
R36886 vdd.n1986 vdd.n1983 61.358
R36887 vdd.n1986 vdd.n1985 61.358
R36888 vdd.n2153 vdd.n2150 61.358
R36889 vdd.n2153 vdd.n2152 61.358
R36890 vdd.n2302 vdd.n2299 61.358
R36891 vdd.n2302 vdd.n2301 61.358
R36892 vdd.n2294 vdd.n2291 61.358
R36893 vdd.n2294 vdd.n2293 61.358
R36894 vdd.n2286 vdd.n2283 61.358
R36895 vdd.n2286 vdd.n2285 61.358
R36896 vdd.n2278 vdd.n2275 61.358
R36897 vdd.n2278 vdd.n2277 61.358
R36898 vdd.n2270 vdd.n2267 61.358
R36899 vdd.n2270 vdd.n2269 61.358
R36900 vdd.n2262 vdd.n2259 61.358
R36901 vdd.n2262 vdd.n2261 61.358
R36902 vdd.n2254 vdd.n2251 61.358
R36903 vdd.n2254 vdd.n2253 61.358
R36904 vdd.n2246 vdd.n2243 61.358
R36905 vdd.n2246 vdd.n2245 61.358
R36906 vdd.n2238 vdd.n2235 61.358
R36907 vdd.n2238 vdd.n2237 61.358
R36908 vdd.n2222 vdd.n2219 61.358
R36909 vdd.n2222 vdd.n2221 61.358
R36910 vdd.n2214 vdd.n2211 61.358
R36911 vdd.n2214 vdd.n2213 61.358
R36912 vdd.n2206 vdd.n2203 61.358
R36913 vdd.n2206 vdd.n2205 61.358
R36914 vdd.n2198 vdd.n2195 61.358
R36915 vdd.n2198 vdd.n2197 61.358
R36916 vdd.n2190 vdd.n2187 61.358
R36917 vdd.n2190 vdd.n2189 61.358
R36918 vdd.n2182 vdd.n2179 61.358
R36919 vdd.n2182 vdd.n2181 61.358
R36920 vdd.n2174 vdd.n2171 61.358
R36921 vdd.n2174 vdd.n2173 61.358
R36922 vdd.n2166 vdd.n2163 61.358
R36923 vdd.n2166 vdd.n2165 61.358
R36924 vdd.n2333 vdd.n2330 61.358
R36925 vdd.n2333 vdd.n2332 61.358
R36926 vdd.n2482 vdd.n2479 61.358
R36927 vdd.n2482 vdd.n2481 61.358
R36928 vdd.n2474 vdd.n2471 61.358
R36929 vdd.n2474 vdd.n2473 61.358
R36930 vdd.n2466 vdd.n2463 61.358
R36931 vdd.n2466 vdd.n2465 61.358
R36932 vdd.n2458 vdd.n2455 61.358
R36933 vdd.n2458 vdd.n2457 61.358
R36934 vdd.n2450 vdd.n2447 61.358
R36935 vdd.n2450 vdd.n2449 61.358
R36936 vdd.n2442 vdd.n2439 61.358
R36937 vdd.n2442 vdd.n2441 61.358
R36938 vdd.n2434 vdd.n2431 61.358
R36939 vdd.n2434 vdd.n2433 61.358
R36940 vdd.n2426 vdd.n2423 61.358
R36941 vdd.n2426 vdd.n2425 61.358
R36942 vdd.n2418 vdd.n2415 61.358
R36943 vdd.n2418 vdd.n2417 61.358
R36944 vdd.n2402 vdd.n2399 61.358
R36945 vdd.n2402 vdd.n2401 61.358
R36946 vdd.n2394 vdd.n2391 61.358
R36947 vdd.n2394 vdd.n2393 61.358
R36948 vdd.n2386 vdd.n2383 61.358
R36949 vdd.n2386 vdd.n2385 61.358
R36950 vdd.n2378 vdd.n2375 61.358
R36951 vdd.n2378 vdd.n2377 61.358
R36952 vdd.n2370 vdd.n2367 61.358
R36953 vdd.n2370 vdd.n2369 61.358
R36954 vdd.n2362 vdd.n2359 61.358
R36955 vdd.n2362 vdd.n2361 61.358
R36956 vdd.n2354 vdd.n2351 61.358
R36957 vdd.n2354 vdd.n2353 61.358
R36958 vdd.n2346 vdd.n2343 61.358
R36959 vdd.n2346 vdd.n2345 61.358
R36960 vdd.n2513 vdd.n2510 61.358
R36961 vdd.n2513 vdd.n2512 61.358
R36962 vdd.n2662 vdd.n2659 61.358
R36963 vdd.n2662 vdd.n2661 61.358
R36964 vdd.n2654 vdd.n2651 61.358
R36965 vdd.n2654 vdd.n2653 61.358
R36966 vdd.n2646 vdd.n2643 61.358
R36967 vdd.n2646 vdd.n2645 61.358
R36968 vdd.n2638 vdd.n2635 61.358
R36969 vdd.n2638 vdd.n2637 61.358
R36970 vdd.n2630 vdd.n2627 61.358
R36971 vdd.n2630 vdd.n2629 61.358
R36972 vdd.n2622 vdd.n2619 61.358
R36973 vdd.n2622 vdd.n2621 61.358
R36974 vdd.n2614 vdd.n2611 61.358
R36975 vdd.n2614 vdd.n2613 61.358
R36976 vdd.n2606 vdd.n2603 61.358
R36977 vdd.n2606 vdd.n2605 61.358
R36978 vdd.n2598 vdd.n2595 61.358
R36979 vdd.n2598 vdd.n2597 61.358
R36980 vdd.n2582 vdd.n2579 61.358
R36981 vdd.n2582 vdd.n2581 61.358
R36982 vdd.n2574 vdd.n2571 61.358
R36983 vdd.n2574 vdd.n2573 61.358
R36984 vdd.n2566 vdd.n2563 61.358
R36985 vdd.n2566 vdd.n2565 61.358
R36986 vdd.n2558 vdd.n2555 61.358
R36987 vdd.n2558 vdd.n2557 61.358
R36988 vdd.n2550 vdd.n2547 61.358
R36989 vdd.n2550 vdd.n2549 61.358
R36990 vdd.n2542 vdd.n2539 61.358
R36991 vdd.n2542 vdd.n2541 61.358
R36992 vdd.n2534 vdd.n2531 61.358
R36993 vdd.n2534 vdd.n2533 61.358
R36994 vdd.n2526 vdd.n2523 61.358
R36995 vdd.n2526 vdd.n2525 61.358
R36996 vdd.n2693 vdd.n2690 61.358
R36997 vdd.n2693 vdd.n2692 61.358
R36998 vdd.n2842 vdd.n2839 61.358
R36999 vdd.n2842 vdd.n2841 61.358
R37000 vdd.n2834 vdd.n2831 61.358
R37001 vdd.n2834 vdd.n2833 61.358
R37002 vdd.n2826 vdd.n2823 61.358
R37003 vdd.n2826 vdd.n2825 61.358
R37004 vdd.n2818 vdd.n2815 61.358
R37005 vdd.n2818 vdd.n2817 61.358
R37006 vdd.n2810 vdd.n2807 61.358
R37007 vdd.n2810 vdd.n2809 61.358
R37008 vdd.n2802 vdd.n2799 61.358
R37009 vdd.n2802 vdd.n2801 61.358
R37010 vdd.n2794 vdd.n2791 61.358
R37011 vdd.n2794 vdd.n2793 61.358
R37012 vdd.n2786 vdd.n2783 61.358
R37013 vdd.n2786 vdd.n2785 61.358
R37014 vdd.n2778 vdd.n2775 61.358
R37015 vdd.n2778 vdd.n2777 61.358
R37016 vdd.n2762 vdd.n2759 61.358
R37017 vdd.n2762 vdd.n2761 61.358
R37018 vdd.n2754 vdd.n2751 61.358
R37019 vdd.n2754 vdd.n2753 61.358
R37020 vdd.n2746 vdd.n2743 61.358
R37021 vdd.n2746 vdd.n2745 61.358
R37022 vdd.n2738 vdd.n2735 61.358
R37023 vdd.n2738 vdd.n2737 61.358
R37024 vdd.n2730 vdd.n2727 61.358
R37025 vdd.n2730 vdd.n2729 61.358
R37026 vdd.n2722 vdd.n2719 61.358
R37027 vdd.n2722 vdd.n2721 61.358
R37028 vdd.n2714 vdd.n2711 61.358
R37029 vdd.n2714 vdd.n2713 61.358
R37030 vdd.n2706 vdd.n2703 61.358
R37031 vdd.n2706 vdd.n2705 61.358
R37032 vdd.n2873 vdd.n2870 61.358
R37033 vdd.n2873 vdd.n2872 61.358
R37034 vdd.n3022 vdd.n3019 61.358
R37035 vdd.n3022 vdd.n3021 61.358
R37036 vdd.n3014 vdd.n3011 61.358
R37037 vdd.n3014 vdd.n3013 61.358
R37038 vdd.n3006 vdd.n3003 61.358
R37039 vdd.n3006 vdd.n3005 61.358
R37040 vdd.n2998 vdd.n2995 61.358
R37041 vdd.n2998 vdd.n2997 61.358
R37042 vdd.n2990 vdd.n2987 61.358
R37043 vdd.n2990 vdd.n2989 61.358
R37044 vdd.n2982 vdd.n2979 61.358
R37045 vdd.n2982 vdd.n2981 61.358
R37046 vdd.n2974 vdd.n2971 61.358
R37047 vdd.n2974 vdd.n2973 61.358
R37048 vdd.n2966 vdd.n2963 61.358
R37049 vdd.n2966 vdd.n2965 61.358
R37050 vdd.n2958 vdd.n2955 61.358
R37051 vdd.n2958 vdd.n2957 61.358
R37052 vdd.n2942 vdd.n2939 61.358
R37053 vdd.n2942 vdd.n2941 61.358
R37054 vdd.n2934 vdd.n2931 61.358
R37055 vdd.n2934 vdd.n2933 61.358
R37056 vdd.n2926 vdd.n2923 61.358
R37057 vdd.n2926 vdd.n2925 61.358
R37058 vdd.n2918 vdd.n2915 61.358
R37059 vdd.n2918 vdd.n2917 61.358
R37060 vdd.n2910 vdd.n2907 61.358
R37061 vdd.n2910 vdd.n2909 61.358
R37062 vdd.n2902 vdd.n2899 61.358
R37063 vdd.n2902 vdd.n2901 61.358
R37064 vdd.n2894 vdd.n2891 61.358
R37065 vdd.n2894 vdd.n2893 61.358
R37066 vdd.n2886 vdd.n2883 61.358
R37067 vdd.n2886 vdd.n2885 61.358
R37068 vdd.n3053 vdd.n3050 61.358
R37069 vdd.n3053 vdd.n3052 61.358
R37070 vdd.n3202 vdd.n3199 61.358
R37071 vdd.n3202 vdd.n3201 61.358
R37072 vdd.n3194 vdd.n3191 61.358
R37073 vdd.n3194 vdd.n3193 61.358
R37074 vdd.n3186 vdd.n3183 61.358
R37075 vdd.n3186 vdd.n3185 61.358
R37076 vdd.n3178 vdd.n3175 61.358
R37077 vdd.n3178 vdd.n3177 61.358
R37078 vdd.n3170 vdd.n3167 61.358
R37079 vdd.n3170 vdd.n3169 61.358
R37080 vdd.n3162 vdd.n3159 61.358
R37081 vdd.n3162 vdd.n3161 61.358
R37082 vdd.n3154 vdd.n3151 61.358
R37083 vdd.n3154 vdd.n3153 61.358
R37084 vdd.n3146 vdd.n3143 61.358
R37085 vdd.n3146 vdd.n3145 61.358
R37086 vdd.n3138 vdd.n3135 61.358
R37087 vdd.n3138 vdd.n3137 61.358
R37088 vdd.n3122 vdd.n3119 61.358
R37089 vdd.n3122 vdd.n3121 61.358
R37090 vdd.n3114 vdd.n3111 61.358
R37091 vdd.n3114 vdd.n3113 61.358
R37092 vdd.n3106 vdd.n3103 61.358
R37093 vdd.n3106 vdd.n3105 61.358
R37094 vdd.n3098 vdd.n3095 61.358
R37095 vdd.n3098 vdd.n3097 61.358
R37096 vdd.n3090 vdd.n3087 61.358
R37097 vdd.n3090 vdd.n3089 61.358
R37098 vdd.n3082 vdd.n3079 61.358
R37099 vdd.n3082 vdd.n3081 61.358
R37100 vdd.n3074 vdd.n3071 61.358
R37101 vdd.n3074 vdd.n3073 61.358
R37102 vdd.n3066 vdd.n3063 61.358
R37103 vdd.n3066 vdd.n3065 61.358
R37104 vdd.n3233 vdd.n3230 61.358
R37105 vdd.n3233 vdd.n3232 61.358
R37106 vdd.n3382 vdd.n3379 61.358
R37107 vdd.n3382 vdd.n3381 61.358
R37108 vdd.n3374 vdd.n3371 61.358
R37109 vdd.n3374 vdd.n3373 61.358
R37110 vdd.n3366 vdd.n3363 61.358
R37111 vdd.n3366 vdd.n3365 61.358
R37112 vdd.n3358 vdd.n3355 61.358
R37113 vdd.n3358 vdd.n3357 61.358
R37114 vdd.n3350 vdd.n3347 61.358
R37115 vdd.n3350 vdd.n3349 61.358
R37116 vdd.n3342 vdd.n3339 61.358
R37117 vdd.n3342 vdd.n3341 61.358
R37118 vdd.n3334 vdd.n3331 61.358
R37119 vdd.n3334 vdd.n3333 61.358
R37120 vdd.n3326 vdd.n3323 61.358
R37121 vdd.n3326 vdd.n3325 61.358
R37122 vdd.n3318 vdd.n3315 61.358
R37123 vdd.n3318 vdd.n3317 61.358
R37124 vdd.n3302 vdd.n3299 61.358
R37125 vdd.n3302 vdd.n3301 61.358
R37126 vdd.n3294 vdd.n3291 61.358
R37127 vdd.n3294 vdd.n3293 61.358
R37128 vdd.n3286 vdd.n3283 61.358
R37129 vdd.n3286 vdd.n3285 61.358
R37130 vdd.n3278 vdd.n3275 61.358
R37131 vdd.n3278 vdd.n3277 61.358
R37132 vdd.n3270 vdd.n3267 61.358
R37133 vdd.n3270 vdd.n3269 61.358
R37134 vdd.n3262 vdd.n3259 61.358
R37135 vdd.n3262 vdd.n3261 61.358
R37136 vdd.n3254 vdd.n3251 61.358
R37137 vdd.n3254 vdd.n3253 61.358
R37138 vdd.n3246 vdd.n3243 61.358
R37139 vdd.n3246 vdd.n3245 61.358
R37140 vdd.n3413 vdd.n3410 61.358
R37141 vdd.n3413 vdd.n3412 61.358
R37142 vdd.n3562 vdd.n3559 61.358
R37143 vdd.n3562 vdd.n3561 61.358
R37144 vdd.n3554 vdd.n3551 61.358
R37145 vdd.n3554 vdd.n3553 61.358
R37146 vdd.n3546 vdd.n3543 61.358
R37147 vdd.n3546 vdd.n3545 61.358
R37148 vdd.n3538 vdd.n3535 61.358
R37149 vdd.n3538 vdd.n3537 61.358
R37150 vdd.n3530 vdd.n3527 61.358
R37151 vdd.n3530 vdd.n3529 61.358
R37152 vdd.n3522 vdd.n3519 61.358
R37153 vdd.n3522 vdd.n3521 61.358
R37154 vdd.n3514 vdd.n3511 61.358
R37155 vdd.n3514 vdd.n3513 61.358
R37156 vdd.n3506 vdd.n3503 61.358
R37157 vdd.n3506 vdd.n3505 61.358
R37158 vdd.n3498 vdd.n3495 61.358
R37159 vdd.n3498 vdd.n3497 61.358
R37160 vdd.n3482 vdd.n3479 61.358
R37161 vdd.n3482 vdd.n3481 61.358
R37162 vdd.n3474 vdd.n3471 61.358
R37163 vdd.n3474 vdd.n3473 61.358
R37164 vdd.n3466 vdd.n3463 61.358
R37165 vdd.n3466 vdd.n3465 61.358
R37166 vdd.n3458 vdd.n3455 61.358
R37167 vdd.n3458 vdd.n3457 61.358
R37168 vdd.n3450 vdd.n3447 61.358
R37169 vdd.n3450 vdd.n3449 61.358
R37170 vdd.n3442 vdd.n3439 61.358
R37171 vdd.n3442 vdd.n3441 61.358
R37172 vdd.n3434 vdd.n3431 61.358
R37173 vdd.n3434 vdd.n3433 61.358
R37174 vdd.n3426 vdd.n3423 61.358
R37175 vdd.n3426 vdd.n3425 61.358
R37176 vdd.n3593 vdd.n3590 61.358
R37177 vdd.n3593 vdd.n3592 61.358
R37178 vdd.n3742 vdd.n3739 61.358
R37179 vdd.n3742 vdd.n3741 61.358
R37180 vdd.n3734 vdd.n3731 61.358
R37181 vdd.n3734 vdd.n3733 61.358
R37182 vdd.n3726 vdd.n3723 61.358
R37183 vdd.n3726 vdd.n3725 61.358
R37184 vdd.n3718 vdd.n3715 61.358
R37185 vdd.n3718 vdd.n3717 61.358
R37186 vdd.n3710 vdd.n3707 61.358
R37187 vdd.n3710 vdd.n3709 61.358
R37188 vdd.n3702 vdd.n3699 61.358
R37189 vdd.n3702 vdd.n3701 61.358
R37190 vdd.n3694 vdd.n3691 61.358
R37191 vdd.n3694 vdd.n3693 61.358
R37192 vdd.n3686 vdd.n3683 61.358
R37193 vdd.n3686 vdd.n3685 61.358
R37194 vdd.n3678 vdd.n3675 61.358
R37195 vdd.n3678 vdd.n3677 61.358
R37196 vdd.n3662 vdd.n3659 61.358
R37197 vdd.n3662 vdd.n3661 61.358
R37198 vdd.n3654 vdd.n3651 61.358
R37199 vdd.n3654 vdd.n3653 61.358
R37200 vdd.n3646 vdd.n3643 61.358
R37201 vdd.n3646 vdd.n3645 61.358
R37202 vdd.n3638 vdd.n3635 61.358
R37203 vdd.n3638 vdd.n3637 61.358
R37204 vdd.n3630 vdd.n3627 61.358
R37205 vdd.n3630 vdd.n3629 61.358
R37206 vdd.n3622 vdd.n3619 61.358
R37207 vdd.n3622 vdd.n3621 61.358
R37208 vdd.n3614 vdd.n3611 61.358
R37209 vdd.n3614 vdd.n3613 61.358
R37210 vdd.n3606 vdd.n3603 61.358
R37211 vdd.n3606 vdd.n3605 61.358
R37212 vdd.n3773 vdd.n3770 61.358
R37213 vdd.n3773 vdd.n3772 61.358
R37214 vdd.n3922 vdd.n3919 61.358
R37215 vdd.n3922 vdd.n3921 61.358
R37216 vdd.n3914 vdd.n3911 61.358
R37217 vdd.n3914 vdd.n3913 61.358
R37218 vdd.n3906 vdd.n3903 61.358
R37219 vdd.n3906 vdd.n3905 61.358
R37220 vdd.n3898 vdd.n3895 61.358
R37221 vdd.n3898 vdd.n3897 61.358
R37222 vdd.n3890 vdd.n3887 61.358
R37223 vdd.n3890 vdd.n3889 61.358
R37224 vdd.n3882 vdd.n3879 61.358
R37225 vdd.n3882 vdd.n3881 61.358
R37226 vdd.n3874 vdd.n3871 61.358
R37227 vdd.n3874 vdd.n3873 61.358
R37228 vdd.n3866 vdd.n3863 61.358
R37229 vdd.n3866 vdd.n3865 61.358
R37230 vdd.n3858 vdd.n3855 61.358
R37231 vdd.n3858 vdd.n3857 61.358
R37232 vdd.n3842 vdd.n3839 61.358
R37233 vdd.n3842 vdd.n3841 61.358
R37234 vdd.n3834 vdd.n3831 61.358
R37235 vdd.n3834 vdd.n3833 61.358
R37236 vdd.n3826 vdd.n3823 61.358
R37237 vdd.n3826 vdd.n3825 61.358
R37238 vdd.n3818 vdd.n3815 61.358
R37239 vdd.n3818 vdd.n3817 61.358
R37240 vdd.n3810 vdd.n3807 61.358
R37241 vdd.n3810 vdd.n3809 61.358
R37242 vdd.n3802 vdd.n3799 61.358
R37243 vdd.n3802 vdd.n3801 61.358
R37244 vdd.n3794 vdd.n3791 61.358
R37245 vdd.n3794 vdd.n3793 61.358
R37246 vdd.n3786 vdd.n3783 61.358
R37247 vdd.n3786 vdd.n3785 61.358
R37248 vdd.n3953 vdd.n3950 61.358
R37249 vdd.n3953 vdd.n3952 61.358
R37250 vdd.n4102 vdd.n4099 61.358
R37251 vdd.n4102 vdd.n4101 61.358
R37252 vdd.n4094 vdd.n4091 61.358
R37253 vdd.n4094 vdd.n4093 61.358
R37254 vdd.n4086 vdd.n4083 61.358
R37255 vdd.n4086 vdd.n4085 61.358
R37256 vdd.n4078 vdd.n4075 61.358
R37257 vdd.n4078 vdd.n4077 61.358
R37258 vdd.n4070 vdd.n4067 61.358
R37259 vdd.n4070 vdd.n4069 61.358
R37260 vdd.n4062 vdd.n4059 61.358
R37261 vdd.n4062 vdd.n4061 61.358
R37262 vdd.n4054 vdd.n4051 61.358
R37263 vdd.n4054 vdd.n4053 61.358
R37264 vdd.n4046 vdd.n4043 61.358
R37265 vdd.n4046 vdd.n4045 61.358
R37266 vdd.n4038 vdd.n4035 61.358
R37267 vdd.n4038 vdd.n4037 61.358
R37268 vdd.n4022 vdd.n4019 61.358
R37269 vdd.n4022 vdd.n4021 61.358
R37270 vdd.n4014 vdd.n4011 61.358
R37271 vdd.n4014 vdd.n4013 61.358
R37272 vdd.n4006 vdd.n4003 61.358
R37273 vdd.n4006 vdd.n4005 61.358
R37274 vdd.n3998 vdd.n3995 61.358
R37275 vdd.n3998 vdd.n3997 61.358
R37276 vdd.n3990 vdd.n3987 61.358
R37277 vdd.n3990 vdd.n3989 61.358
R37278 vdd.n3982 vdd.n3979 61.358
R37279 vdd.n3982 vdd.n3981 61.358
R37280 vdd.n3974 vdd.n3971 61.358
R37281 vdd.n3974 vdd.n3973 61.358
R37282 vdd.n3966 vdd.n3963 61.358
R37283 vdd.n3966 vdd.n3965 61.358
R37284 vdd.n4133 vdd.n4130 61.358
R37285 vdd.n4133 vdd.n4132 61.358
R37286 vdd.n4282 vdd.n4279 61.358
R37287 vdd.n4282 vdd.n4281 61.358
R37288 vdd.n4274 vdd.n4271 61.358
R37289 vdd.n4274 vdd.n4273 61.358
R37290 vdd.n4266 vdd.n4263 61.358
R37291 vdd.n4266 vdd.n4265 61.358
R37292 vdd.n4258 vdd.n4255 61.358
R37293 vdd.n4258 vdd.n4257 61.358
R37294 vdd.n4250 vdd.n4247 61.358
R37295 vdd.n4250 vdd.n4249 61.358
R37296 vdd.n4242 vdd.n4239 61.358
R37297 vdd.n4242 vdd.n4241 61.358
R37298 vdd.n4234 vdd.n4231 61.358
R37299 vdd.n4234 vdd.n4233 61.358
R37300 vdd.n4226 vdd.n4223 61.358
R37301 vdd.n4226 vdd.n4225 61.358
R37302 vdd.n4218 vdd.n4215 61.358
R37303 vdd.n4218 vdd.n4217 61.358
R37304 vdd.n4202 vdd.n4199 61.358
R37305 vdd.n4202 vdd.n4201 61.358
R37306 vdd.n4194 vdd.n4191 61.358
R37307 vdd.n4194 vdd.n4193 61.358
R37308 vdd.n4186 vdd.n4183 61.358
R37309 vdd.n4186 vdd.n4185 61.358
R37310 vdd.n4178 vdd.n4175 61.358
R37311 vdd.n4178 vdd.n4177 61.358
R37312 vdd.n4170 vdd.n4167 61.358
R37313 vdd.n4170 vdd.n4169 61.358
R37314 vdd.n4162 vdd.n4159 61.358
R37315 vdd.n4162 vdd.n4161 61.358
R37316 vdd.n4154 vdd.n4151 61.358
R37317 vdd.n4154 vdd.n4153 61.358
R37318 vdd.n4146 vdd.n4143 61.358
R37319 vdd.n4146 vdd.n4145 61.358
R37320 vdd.n4313 vdd.n4310 61.358
R37321 vdd.n4313 vdd.n4312 61.358
R37322 vdd.n4462 vdd.n4459 61.358
R37323 vdd.n4462 vdd.n4461 61.358
R37324 vdd.n4454 vdd.n4451 61.358
R37325 vdd.n4454 vdd.n4453 61.358
R37326 vdd.n4446 vdd.n4443 61.358
R37327 vdd.n4446 vdd.n4445 61.358
R37328 vdd.n4438 vdd.n4435 61.358
R37329 vdd.n4438 vdd.n4437 61.358
R37330 vdd.n4430 vdd.n4427 61.358
R37331 vdd.n4430 vdd.n4429 61.358
R37332 vdd.n4422 vdd.n4419 61.358
R37333 vdd.n4422 vdd.n4421 61.358
R37334 vdd.n4414 vdd.n4411 61.358
R37335 vdd.n4414 vdd.n4413 61.358
R37336 vdd.n4406 vdd.n4403 61.358
R37337 vdd.n4406 vdd.n4405 61.358
R37338 vdd.n4398 vdd.n4395 61.358
R37339 vdd.n4398 vdd.n4397 61.358
R37340 vdd.n4382 vdd.n4379 61.358
R37341 vdd.n4382 vdd.n4381 61.358
R37342 vdd.n4374 vdd.n4371 61.358
R37343 vdd.n4374 vdd.n4373 61.358
R37344 vdd.n4366 vdd.n4363 61.358
R37345 vdd.n4366 vdd.n4365 61.358
R37346 vdd.n4358 vdd.n4355 61.358
R37347 vdd.n4358 vdd.n4357 61.358
R37348 vdd.n4350 vdd.n4347 61.358
R37349 vdd.n4350 vdd.n4349 61.358
R37350 vdd.n4342 vdd.n4339 61.358
R37351 vdd.n4342 vdd.n4341 61.358
R37352 vdd.n4334 vdd.n4331 61.358
R37353 vdd.n4334 vdd.n4333 61.358
R37354 vdd.n4326 vdd.n4323 61.358
R37355 vdd.n4326 vdd.n4325 61.358
R37356 vdd.n4493 vdd.n4490 61.358
R37357 vdd.n4493 vdd.n4492 61.358
R37358 vdd.n4642 vdd.n4639 61.358
R37359 vdd.n4642 vdd.n4641 61.358
R37360 vdd.n4634 vdd.n4631 61.358
R37361 vdd.n4634 vdd.n4633 61.358
R37362 vdd.n4626 vdd.n4623 61.358
R37363 vdd.n4626 vdd.n4625 61.358
R37364 vdd.n4618 vdd.n4615 61.358
R37365 vdd.n4618 vdd.n4617 61.358
R37366 vdd.n4610 vdd.n4607 61.358
R37367 vdd.n4610 vdd.n4609 61.358
R37368 vdd.n4602 vdd.n4599 61.358
R37369 vdd.n4602 vdd.n4601 61.358
R37370 vdd.n4594 vdd.n4591 61.358
R37371 vdd.n4594 vdd.n4593 61.358
R37372 vdd.n4586 vdd.n4583 61.358
R37373 vdd.n4586 vdd.n4585 61.358
R37374 vdd.n4578 vdd.n4575 61.358
R37375 vdd.n4578 vdd.n4577 61.358
R37376 vdd.n4562 vdd.n4559 61.358
R37377 vdd.n4562 vdd.n4561 61.358
R37378 vdd.n4554 vdd.n4551 61.358
R37379 vdd.n4554 vdd.n4553 61.358
R37380 vdd.n4546 vdd.n4543 61.358
R37381 vdd.n4546 vdd.n4545 61.358
R37382 vdd.n4538 vdd.n4535 61.358
R37383 vdd.n4538 vdd.n4537 61.358
R37384 vdd.n4530 vdd.n4527 61.358
R37385 vdd.n4530 vdd.n4529 61.358
R37386 vdd.n4522 vdd.n4519 61.358
R37387 vdd.n4522 vdd.n4521 61.358
R37388 vdd.n4514 vdd.n4511 61.358
R37389 vdd.n4514 vdd.n4513 61.358
R37390 vdd.n4506 vdd.n4503 61.358
R37391 vdd.n4506 vdd.n4505 61.358
R37392 vdd.n4673 vdd.n4670 61.358
R37393 vdd.n4673 vdd.n4672 61.358
R37394 vdd.n4822 vdd.n4819 61.358
R37395 vdd.n4822 vdd.n4821 61.358
R37396 vdd.n4814 vdd.n4811 61.358
R37397 vdd.n4814 vdd.n4813 61.358
R37398 vdd.n4806 vdd.n4803 61.358
R37399 vdd.n4806 vdd.n4805 61.358
R37400 vdd.n4798 vdd.n4795 61.358
R37401 vdd.n4798 vdd.n4797 61.358
R37402 vdd.n4790 vdd.n4787 61.358
R37403 vdd.n4790 vdd.n4789 61.358
R37404 vdd.n4782 vdd.n4779 61.358
R37405 vdd.n4782 vdd.n4781 61.358
R37406 vdd.n4774 vdd.n4771 61.358
R37407 vdd.n4774 vdd.n4773 61.358
R37408 vdd.n4766 vdd.n4763 61.358
R37409 vdd.n4766 vdd.n4765 61.358
R37410 vdd.n4758 vdd.n4755 61.358
R37411 vdd.n4758 vdd.n4757 61.358
R37412 vdd.n4742 vdd.n4739 61.358
R37413 vdd.n4742 vdd.n4741 61.358
R37414 vdd.n4734 vdd.n4731 61.358
R37415 vdd.n4734 vdd.n4733 61.358
R37416 vdd.n4726 vdd.n4723 61.358
R37417 vdd.n4726 vdd.n4725 61.358
R37418 vdd.n4718 vdd.n4715 61.358
R37419 vdd.n4718 vdd.n4717 61.358
R37420 vdd.n4710 vdd.n4707 61.358
R37421 vdd.n4710 vdd.n4709 61.358
R37422 vdd.n4702 vdd.n4699 61.358
R37423 vdd.n4702 vdd.n4701 61.358
R37424 vdd.n4694 vdd.n4691 61.358
R37425 vdd.n4694 vdd.n4693 61.358
R37426 vdd.n4686 vdd.n4683 61.358
R37427 vdd.n4686 vdd.n4685 61.358
R37428 vdd.n4853 vdd.n4850 61.358
R37429 vdd.n4853 vdd.n4852 61.358
R37430 vdd.n5002 vdd.n4999 61.358
R37431 vdd.n5002 vdd.n5001 61.358
R37432 vdd.n4994 vdd.n4991 61.358
R37433 vdd.n4994 vdd.n4993 61.358
R37434 vdd.n4986 vdd.n4983 61.358
R37435 vdd.n4986 vdd.n4985 61.358
R37436 vdd.n4978 vdd.n4975 61.358
R37437 vdd.n4978 vdd.n4977 61.358
R37438 vdd.n4970 vdd.n4967 61.358
R37439 vdd.n4970 vdd.n4969 61.358
R37440 vdd.n4962 vdd.n4959 61.358
R37441 vdd.n4962 vdd.n4961 61.358
R37442 vdd.n4954 vdd.n4951 61.358
R37443 vdd.n4954 vdd.n4953 61.358
R37444 vdd.n4946 vdd.n4943 61.358
R37445 vdd.n4946 vdd.n4945 61.358
R37446 vdd.n4938 vdd.n4935 61.358
R37447 vdd.n4938 vdd.n4937 61.358
R37448 vdd.n4922 vdd.n4919 61.358
R37449 vdd.n4922 vdd.n4921 61.358
R37450 vdd.n4914 vdd.n4911 61.358
R37451 vdd.n4914 vdd.n4913 61.358
R37452 vdd.n4906 vdd.n4903 61.358
R37453 vdd.n4906 vdd.n4905 61.358
R37454 vdd.n4898 vdd.n4895 61.358
R37455 vdd.n4898 vdd.n4897 61.358
R37456 vdd.n4890 vdd.n4887 61.358
R37457 vdd.n4890 vdd.n4889 61.358
R37458 vdd.n4882 vdd.n4879 61.358
R37459 vdd.n4882 vdd.n4881 61.358
R37460 vdd.n4874 vdd.n4871 61.358
R37461 vdd.n4874 vdd.n4873 61.358
R37462 vdd.n4866 vdd.n4863 61.358
R37463 vdd.n4866 vdd.n4865 61.358
R37464 vdd.n5033 vdd.n5030 61.358
R37465 vdd.n5033 vdd.n5032 61.358
R37466 vdd.n5182 vdd.n5179 61.358
R37467 vdd.n5182 vdd.n5181 61.358
R37468 vdd.n5174 vdd.n5171 61.358
R37469 vdd.n5174 vdd.n5173 61.358
R37470 vdd.n5166 vdd.n5163 61.358
R37471 vdd.n5166 vdd.n5165 61.358
R37472 vdd.n5158 vdd.n5155 61.358
R37473 vdd.n5158 vdd.n5157 61.358
R37474 vdd.n5150 vdd.n5147 61.358
R37475 vdd.n5150 vdd.n5149 61.358
R37476 vdd.n5142 vdd.n5139 61.358
R37477 vdd.n5142 vdd.n5141 61.358
R37478 vdd.n5134 vdd.n5131 61.358
R37479 vdd.n5134 vdd.n5133 61.358
R37480 vdd.n5126 vdd.n5123 61.358
R37481 vdd.n5126 vdd.n5125 61.358
R37482 vdd.n5118 vdd.n5115 61.358
R37483 vdd.n5118 vdd.n5117 61.358
R37484 vdd.n5102 vdd.n5099 61.358
R37485 vdd.n5102 vdd.n5101 61.358
R37486 vdd.n5094 vdd.n5091 61.358
R37487 vdd.n5094 vdd.n5093 61.358
R37488 vdd.n5086 vdd.n5083 61.358
R37489 vdd.n5086 vdd.n5085 61.358
R37490 vdd.n5078 vdd.n5075 61.358
R37491 vdd.n5078 vdd.n5077 61.358
R37492 vdd.n5070 vdd.n5067 61.358
R37493 vdd.n5070 vdd.n5069 61.358
R37494 vdd.n5062 vdd.n5059 61.358
R37495 vdd.n5062 vdd.n5061 61.358
R37496 vdd.n5054 vdd.n5051 61.358
R37497 vdd.n5054 vdd.n5053 61.358
R37498 vdd.n5046 vdd.n5043 61.358
R37499 vdd.n5046 vdd.n5045 61.358
R37500 vdd.n5213 vdd.n5210 61.358
R37501 vdd.n5213 vdd.n5212 61.358
R37502 vdd.n5362 vdd.n5359 61.358
R37503 vdd.n5362 vdd.n5361 61.358
R37504 vdd.n5354 vdd.n5351 61.358
R37505 vdd.n5354 vdd.n5353 61.358
R37506 vdd.n5346 vdd.n5343 61.358
R37507 vdd.n5346 vdd.n5345 61.358
R37508 vdd.n5338 vdd.n5335 61.358
R37509 vdd.n5338 vdd.n5337 61.358
R37510 vdd.n5330 vdd.n5327 61.358
R37511 vdd.n5330 vdd.n5329 61.358
R37512 vdd.n5322 vdd.n5319 61.358
R37513 vdd.n5322 vdd.n5321 61.358
R37514 vdd.n5314 vdd.n5311 61.358
R37515 vdd.n5314 vdd.n5313 61.358
R37516 vdd.n5306 vdd.n5303 61.358
R37517 vdd.n5306 vdd.n5305 61.358
R37518 vdd.n5298 vdd.n5295 61.358
R37519 vdd.n5298 vdd.n5297 61.358
R37520 vdd.n5282 vdd.n5279 61.358
R37521 vdd.n5282 vdd.n5281 61.358
R37522 vdd.n5274 vdd.n5271 61.358
R37523 vdd.n5274 vdd.n5273 61.358
R37524 vdd.n5266 vdd.n5263 61.358
R37525 vdd.n5266 vdd.n5265 61.358
R37526 vdd.n5258 vdd.n5255 61.358
R37527 vdd.n5258 vdd.n5257 61.358
R37528 vdd.n5250 vdd.n5247 61.358
R37529 vdd.n5250 vdd.n5249 61.358
R37530 vdd.n5242 vdd.n5239 61.358
R37531 vdd.n5242 vdd.n5241 61.358
R37532 vdd.n5234 vdd.n5231 61.358
R37533 vdd.n5234 vdd.n5233 61.358
R37534 vdd.n5226 vdd.n5223 61.358
R37535 vdd.n5226 vdd.n5225 61.358
R37536 vdd.n5393 vdd.n5390 61.358
R37537 vdd.n5393 vdd.n5392 61.358
R37538 vdd.n5542 vdd.n5539 61.358
R37539 vdd.n5542 vdd.n5541 61.358
R37540 vdd.n5534 vdd.n5531 61.358
R37541 vdd.n5534 vdd.n5533 61.358
R37542 vdd.n5526 vdd.n5523 61.358
R37543 vdd.n5526 vdd.n5525 61.358
R37544 vdd.n5518 vdd.n5515 61.358
R37545 vdd.n5518 vdd.n5517 61.358
R37546 vdd.n5510 vdd.n5507 61.358
R37547 vdd.n5510 vdd.n5509 61.358
R37548 vdd.n5502 vdd.n5499 61.358
R37549 vdd.n5502 vdd.n5501 61.358
R37550 vdd.n5494 vdd.n5491 61.358
R37551 vdd.n5494 vdd.n5493 61.358
R37552 vdd.n5486 vdd.n5483 61.358
R37553 vdd.n5486 vdd.n5485 61.358
R37554 vdd.n5478 vdd.n5475 61.358
R37555 vdd.n5478 vdd.n5477 61.358
R37556 vdd.n5462 vdd.n5459 61.358
R37557 vdd.n5462 vdd.n5461 61.358
R37558 vdd.n5454 vdd.n5451 61.358
R37559 vdd.n5454 vdd.n5453 61.358
R37560 vdd.n5446 vdd.n5443 61.358
R37561 vdd.n5446 vdd.n5445 61.358
R37562 vdd.n5438 vdd.n5435 61.358
R37563 vdd.n5438 vdd.n5437 61.358
R37564 vdd.n5430 vdd.n5427 61.358
R37565 vdd.n5430 vdd.n5429 61.358
R37566 vdd.n5422 vdd.n5419 61.358
R37567 vdd.n5422 vdd.n5421 61.358
R37568 vdd.n5414 vdd.n5411 61.358
R37569 vdd.n5414 vdd.n5413 61.358
R37570 vdd.n5406 vdd.n5403 61.358
R37571 vdd.n5406 vdd.n5405 61.358
R37572 vdd.n5573 vdd.n5570 61.358
R37573 vdd.n5573 vdd.n5572 61.358
R37574 vdd.n5722 vdd.n5719 61.358
R37575 vdd.n5722 vdd.n5721 61.358
R37576 vdd.n5714 vdd.n5711 61.358
R37577 vdd.n5714 vdd.n5713 61.358
R37578 vdd.n5706 vdd.n5703 61.358
R37579 vdd.n5706 vdd.n5705 61.358
R37580 vdd.n5698 vdd.n5695 61.358
R37581 vdd.n5698 vdd.n5697 61.358
R37582 vdd.n5690 vdd.n5687 61.358
R37583 vdd.n5690 vdd.n5689 61.358
R37584 vdd.n5682 vdd.n5679 61.358
R37585 vdd.n5682 vdd.n5681 61.358
R37586 vdd.n5674 vdd.n5671 61.358
R37587 vdd.n5674 vdd.n5673 61.358
R37588 vdd.n5666 vdd.n5663 61.358
R37589 vdd.n5666 vdd.n5665 61.358
R37590 vdd.n5658 vdd.n5655 61.358
R37591 vdd.n5658 vdd.n5657 61.358
R37592 vdd.n5642 vdd.n5639 61.358
R37593 vdd.n5642 vdd.n5641 61.358
R37594 vdd.n5634 vdd.n5631 61.358
R37595 vdd.n5634 vdd.n5633 61.358
R37596 vdd.n5626 vdd.n5623 61.358
R37597 vdd.n5626 vdd.n5625 61.358
R37598 vdd.n5618 vdd.n5615 61.358
R37599 vdd.n5618 vdd.n5617 61.358
R37600 vdd.n5610 vdd.n5607 61.358
R37601 vdd.n5610 vdd.n5609 61.358
R37602 vdd.n5602 vdd.n5599 61.358
R37603 vdd.n5602 vdd.n5601 61.358
R37604 vdd.n5594 vdd.n5591 61.358
R37605 vdd.n5594 vdd.n5593 61.358
R37606 vdd.n5586 vdd.n5583 61.358
R37607 vdd.n5586 vdd.n5585 61.358
R37608 vdd.n5753 vdd.n5750 61.358
R37609 vdd.n5753 vdd.n5752 61.358
R37610 vdd.n5902 vdd.n5899 61.358
R37611 vdd.n5902 vdd.n5901 61.358
R37612 vdd.n5894 vdd.n5891 61.358
R37613 vdd.n5894 vdd.n5893 61.358
R37614 vdd.n5886 vdd.n5883 61.358
R37615 vdd.n5886 vdd.n5885 61.358
R37616 vdd.n5878 vdd.n5875 61.358
R37617 vdd.n5878 vdd.n5877 61.358
R37618 vdd.n5870 vdd.n5867 61.358
R37619 vdd.n5870 vdd.n5869 61.358
R37620 vdd.n5862 vdd.n5859 61.358
R37621 vdd.n5862 vdd.n5861 61.358
R37622 vdd.n5854 vdd.n5851 61.358
R37623 vdd.n5854 vdd.n5853 61.358
R37624 vdd.n5846 vdd.n5843 61.358
R37625 vdd.n5846 vdd.n5845 61.358
R37626 vdd.n5838 vdd.n5835 61.358
R37627 vdd.n5838 vdd.n5837 61.358
R37628 vdd.n5822 vdd.n5819 61.358
R37629 vdd.n5822 vdd.n5821 61.358
R37630 vdd.n5814 vdd.n5811 61.358
R37631 vdd.n5814 vdd.n5813 61.358
R37632 vdd.n5806 vdd.n5803 61.358
R37633 vdd.n5806 vdd.n5805 61.358
R37634 vdd.n5798 vdd.n5795 61.358
R37635 vdd.n5798 vdd.n5797 61.358
R37636 vdd.n5790 vdd.n5787 61.358
R37637 vdd.n5790 vdd.n5789 61.358
R37638 vdd.n5782 vdd.n5779 61.358
R37639 vdd.n5782 vdd.n5781 61.358
R37640 vdd.n5774 vdd.n5771 61.358
R37641 vdd.n5774 vdd.n5773 61.358
R37642 vdd.n5766 vdd.n5763 61.358
R37643 vdd.n5766 vdd.n5765 61.358
R37644 vdd.n5933 vdd.n5930 61.358
R37645 vdd.n5933 vdd.n5932 61.358
R37646 vdd.n6082 vdd.n6079 61.358
R37647 vdd.n6082 vdd.n6081 61.358
R37648 vdd.n6074 vdd.n6071 61.358
R37649 vdd.n6074 vdd.n6073 61.358
R37650 vdd.n6066 vdd.n6063 61.358
R37651 vdd.n6066 vdd.n6065 61.358
R37652 vdd.n6058 vdd.n6055 61.358
R37653 vdd.n6058 vdd.n6057 61.358
R37654 vdd.n6050 vdd.n6047 61.358
R37655 vdd.n6050 vdd.n6049 61.358
R37656 vdd.n6042 vdd.n6039 61.358
R37657 vdd.n6042 vdd.n6041 61.358
R37658 vdd.n6034 vdd.n6031 61.358
R37659 vdd.n6034 vdd.n6033 61.358
R37660 vdd.n6026 vdd.n6023 61.358
R37661 vdd.n6026 vdd.n6025 61.358
R37662 vdd.n6018 vdd.n6015 61.358
R37663 vdd.n6018 vdd.n6017 61.358
R37664 vdd.n6002 vdd.n5999 61.358
R37665 vdd.n6002 vdd.n6001 61.358
R37666 vdd.n5994 vdd.n5991 61.358
R37667 vdd.n5994 vdd.n5993 61.358
R37668 vdd.n5986 vdd.n5983 61.358
R37669 vdd.n5986 vdd.n5985 61.358
R37670 vdd.n5978 vdd.n5975 61.358
R37671 vdd.n5978 vdd.n5977 61.358
R37672 vdd.n5970 vdd.n5967 61.358
R37673 vdd.n5970 vdd.n5969 61.358
R37674 vdd.n5962 vdd.n5959 61.358
R37675 vdd.n5962 vdd.n5961 61.358
R37676 vdd.n5954 vdd.n5951 61.358
R37677 vdd.n5954 vdd.n5953 61.358
R37678 vdd.n5946 vdd.n5943 61.358
R37679 vdd.n5946 vdd.n5945 61.358
R37680 vdd.n6113 vdd.n6110 61.358
R37681 vdd.n6113 vdd.n6112 61.358
R37682 vdd.n6262 vdd.n6259 61.358
R37683 vdd.n6262 vdd.n6261 61.358
R37684 vdd.n6254 vdd.n6251 61.358
R37685 vdd.n6254 vdd.n6253 61.358
R37686 vdd.n6246 vdd.n6243 61.358
R37687 vdd.n6246 vdd.n6245 61.358
R37688 vdd.n6238 vdd.n6235 61.358
R37689 vdd.n6238 vdd.n6237 61.358
R37690 vdd.n6230 vdd.n6227 61.358
R37691 vdd.n6230 vdd.n6229 61.358
R37692 vdd.n6222 vdd.n6219 61.358
R37693 vdd.n6222 vdd.n6221 61.358
R37694 vdd.n6214 vdd.n6211 61.358
R37695 vdd.n6214 vdd.n6213 61.358
R37696 vdd.n6206 vdd.n6203 61.358
R37697 vdd.n6206 vdd.n6205 61.358
R37698 vdd.n6198 vdd.n6195 61.358
R37699 vdd.n6198 vdd.n6197 61.358
R37700 vdd.n6182 vdd.n6179 61.358
R37701 vdd.n6182 vdd.n6181 61.358
R37702 vdd.n6174 vdd.n6171 61.358
R37703 vdd.n6174 vdd.n6173 61.358
R37704 vdd.n6166 vdd.n6163 61.358
R37705 vdd.n6166 vdd.n6165 61.358
R37706 vdd.n6158 vdd.n6155 61.358
R37707 vdd.n6158 vdd.n6157 61.358
R37708 vdd.n6150 vdd.n6147 61.358
R37709 vdd.n6150 vdd.n6149 61.358
R37710 vdd.n6142 vdd.n6139 61.358
R37711 vdd.n6142 vdd.n6141 61.358
R37712 vdd.n6134 vdd.n6131 61.358
R37713 vdd.n6134 vdd.n6133 61.358
R37714 vdd.n6126 vdd.n6123 61.358
R37715 vdd.n6126 vdd.n6125 61.358
R37716 vdd.n6293 vdd.n6290 61.358
R37717 vdd.n6293 vdd.n6292 61.358
R37718 vdd.n6442 vdd.n6439 61.358
R37719 vdd.n6442 vdd.n6441 61.358
R37720 vdd.n6434 vdd.n6431 61.358
R37721 vdd.n6434 vdd.n6433 61.358
R37722 vdd.n6426 vdd.n6423 61.358
R37723 vdd.n6426 vdd.n6425 61.358
R37724 vdd.n6418 vdd.n6415 61.358
R37725 vdd.n6418 vdd.n6417 61.358
R37726 vdd.n6410 vdd.n6407 61.358
R37727 vdd.n6410 vdd.n6409 61.358
R37728 vdd.n6402 vdd.n6399 61.358
R37729 vdd.n6402 vdd.n6401 61.358
R37730 vdd.n6394 vdd.n6391 61.358
R37731 vdd.n6394 vdd.n6393 61.358
R37732 vdd.n6386 vdd.n6383 61.358
R37733 vdd.n6386 vdd.n6385 61.358
R37734 vdd.n6378 vdd.n6375 61.358
R37735 vdd.n6378 vdd.n6377 61.358
R37736 vdd.n6362 vdd.n6359 61.358
R37737 vdd.n6362 vdd.n6361 61.358
R37738 vdd.n6354 vdd.n6351 61.358
R37739 vdd.n6354 vdd.n6353 61.358
R37740 vdd.n6346 vdd.n6343 61.358
R37741 vdd.n6346 vdd.n6345 61.358
R37742 vdd.n6338 vdd.n6335 61.358
R37743 vdd.n6338 vdd.n6337 61.358
R37744 vdd.n6330 vdd.n6327 61.358
R37745 vdd.n6330 vdd.n6329 61.358
R37746 vdd.n6322 vdd.n6319 61.358
R37747 vdd.n6322 vdd.n6321 61.358
R37748 vdd.n6314 vdd.n6311 61.358
R37749 vdd.n6314 vdd.n6313 61.358
R37750 vdd.n6306 vdd.n6303 61.358
R37751 vdd.n6306 vdd.n6305 61.358
R37752 vdd.n6473 vdd.n6470 61.358
R37753 vdd.n6473 vdd.n6472 61.358
R37754 vdd.n6622 vdd.n6619 61.358
R37755 vdd.n6622 vdd.n6621 61.358
R37756 vdd.n6614 vdd.n6611 61.358
R37757 vdd.n6614 vdd.n6613 61.358
R37758 vdd.n6606 vdd.n6603 61.358
R37759 vdd.n6606 vdd.n6605 61.358
R37760 vdd.n6598 vdd.n6595 61.358
R37761 vdd.n6598 vdd.n6597 61.358
R37762 vdd.n6590 vdd.n6587 61.358
R37763 vdd.n6590 vdd.n6589 61.358
R37764 vdd.n6582 vdd.n6579 61.358
R37765 vdd.n6582 vdd.n6581 61.358
R37766 vdd.n6574 vdd.n6571 61.358
R37767 vdd.n6574 vdd.n6573 61.358
R37768 vdd.n6566 vdd.n6563 61.358
R37769 vdd.n6566 vdd.n6565 61.358
R37770 vdd.n6558 vdd.n6555 61.358
R37771 vdd.n6558 vdd.n6557 61.358
R37772 vdd.n6542 vdd.n6539 61.358
R37773 vdd.n6542 vdd.n6541 61.358
R37774 vdd.n6534 vdd.n6531 61.358
R37775 vdd.n6534 vdd.n6533 61.358
R37776 vdd.n6526 vdd.n6523 61.358
R37777 vdd.n6526 vdd.n6525 61.358
R37778 vdd.n6518 vdd.n6515 61.358
R37779 vdd.n6518 vdd.n6517 61.358
R37780 vdd.n6510 vdd.n6507 61.358
R37781 vdd.n6510 vdd.n6509 61.358
R37782 vdd.n6502 vdd.n6499 61.358
R37783 vdd.n6502 vdd.n6501 61.358
R37784 vdd.n6494 vdd.n6491 61.358
R37785 vdd.n6494 vdd.n6493 61.358
R37786 vdd.n6486 vdd.n6483 61.358
R37787 vdd.n6486 vdd.n6485 61.358
R37788 vdd.n6653 vdd.n6650 61.358
R37789 vdd.n6653 vdd.n6652 61.358
R37790 vdd.n6802 vdd.n6799 61.358
R37791 vdd.n6802 vdd.n6801 61.358
R37792 vdd.n6794 vdd.n6791 61.358
R37793 vdd.n6794 vdd.n6793 61.358
R37794 vdd.n6786 vdd.n6783 61.358
R37795 vdd.n6786 vdd.n6785 61.358
R37796 vdd.n6778 vdd.n6775 61.358
R37797 vdd.n6778 vdd.n6777 61.358
R37798 vdd.n6770 vdd.n6767 61.358
R37799 vdd.n6770 vdd.n6769 61.358
R37800 vdd.n6762 vdd.n6759 61.358
R37801 vdd.n6762 vdd.n6761 61.358
R37802 vdd.n6754 vdd.n6751 61.358
R37803 vdd.n6754 vdd.n6753 61.358
R37804 vdd.n6746 vdd.n6743 61.358
R37805 vdd.n6746 vdd.n6745 61.358
R37806 vdd.n6738 vdd.n6735 61.358
R37807 vdd.n6738 vdd.n6737 61.358
R37808 vdd.n6722 vdd.n6719 61.358
R37809 vdd.n6722 vdd.n6721 61.358
R37810 vdd.n6714 vdd.n6711 61.358
R37811 vdd.n6714 vdd.n6713 61.358
R37812 vdd.n6706 vdd.n6703 61.358
R37813 vdd.n6706 vdd.n6705 61.358
R37814 vdd.n6698 vdd.n6695 61.358
R37815 vdd.n6698 vdd.n6697 61.358
R37816 vdd.n6690 vdd.n6687 61.358
R37817 vdd.n6690 vdd.n6689 61.358
R37818 vdd.n6682 vdd.n6679 61.358
R37819 vdd.n6682 vdd.n6681 61.358
R37820 vdd.n6674 vdd.n6671 61.358
R37821 vdd.n6674 vdd.n6673 61.358
R37822 vdd.n6666 vdd.n6663 61.358
R37823 vdd.n6666 vdd.n6665 61.358
R37824 vdd.n6833 vdd.n6830 61.358
R37825 vdd.n6833 vdd.n6832 61.358
R37826 vdd.n6982 vdd.n6979 61.358
R37827 vdd.n6982 vdd.n6981 61.358
R37828 vdd.n6974 vdd.n6971 61.358
R37829 vdd.n6974 vdd.n6973 61.358
R37830 vdd.n6966 vdd.n6963 61.358
R37831 vdd.n6966 vdd.n6965 61.358
R37832 vdd.n6958 vdd.n6955 61.358
R37833 vdd.n6958 vdd.n6957 61.358
R37834 vdd.n6950 vdd.n6947 61.358
R37835 vdd.n6950 vdd.n6949 61.358
R37836 vdd.n6942 vdd.n6939 61.358
R37837 vdd.n6942 vdd.n6941 61.358
R37838 vdd.n6934 vdd.n6931 61.358
R37839 vdd.n6934 vdd.n6933 61.358
R37840 vdd.n6926 vdd.n6923 61.358
R37841 vdd.n6926 vdd.n6925 61.358
R37842 vdd.n6918 vdd.n6915 61.358
R37843 vdd.n6918 vdd.n6917 61.358
R37844 vdd.n6902 vdd.n6899 61.358
R37845 vdd.n6902 vdd.n6901 61.358
R37846 vdd.n6894 vdd.n6891 61.358
R37847 vdd.n6894 vdd.n6893 61.358
R37848 vdd.n6886 vdd.n6883 61.358
R37849 vdd.n6886 vdd.n6885 61.358
R37850 vdd.n6878 vdd.n6875 61.358
R37851 vdd.n6878 vdd.n6877 61.358
R37852 vdd.n6870 vdd.n6867 61.358
R37853 vdd.n6870 vdd.n6869 61.358
R37854 vdd.n6862 vdd.n6859 61.358
R37855 vdd.n6862 vdd.n6861 61.358
R37856 vdd.n6854 vdd.n6851 61.358
R37857 vdd.n6854 vdd.n6853 61.358
R37858 vdd.n6846 vdd.n6843 61.358
R37859 vdd.n6846 vdd.n6845 61.358
R37860 vdd.n7013 vdd.n7010 61.358
R37861 vdd.n7013 vdd.n7012 61.358
R37862 vdd.n7162 vdd.n7159 61.358
R37863 vdd.n7162 vdd.n7161 61.358
R37864 vdd.n7154 vdd.n7151 61.358
R37865 vdd.n7154 vdd.n7153 61.358
R37866 vdd.n7146 vdd.n7143 61.358
R37867 vdd.n7146 vdd.n7145 61.358
R37868 vdd.n7138 vdd.n7135 61.358
R37869 vdd.n7138 vdd.n7137 61.358
R37870 vdd.n7130 vdd.n7127 61.358
R37871 vdd.n7130 vdd.n7129 61.358
R37872 vdd.n7122 vdd.n7119 61.358
R37873 vdd.n7122 vdd.n7121 61.358
R37874 vdd.n7114 vdd.n7111 61.358
R37875 vdd.n7114 vdd.n7113 61.358
R37876 vdd.n7106 vdd.n7103 61.358
R37877 vdd.n7106 vdd.n7105 61.358
R37878 vdd.n7098 vdd.n7095 61.358
R37879 vdd.n7098 vdd.n7097 61.358
R37880 vdd.n7082 vdd.n7079 61.358
R37881 vdd.n7082 vdd.n7081 61.358
R37882 vdd.n7074 vdd.n7071 61.358
R37883 vdd.n7074 vdd.n7073 61.358
R37884 vdd.n7066 vdd.n7063 61.358
R37885 vdd.n7066 vdd.n7065 61.358
R37886 vdd.n7058 vdd.n7055 61.358
R37887 vdd.n7058 vdd.n7057 61.358
R37888 vdd.n7050 vdd.n7047 61.358
R37889 vdd.n7050 vdd.n7049 61.358
R37890 vdd.n7042 vdd.n7039 61.358
R37891 vdd.n7042 vdd.n7041 61.358
R37892 vdd.n7034 vdd.n7031 61.358
R37893 vdd.n7034 vdd.n7033 61.358
R37894 vdd.n7026 vdd.n7023 61.358
R37895 vdd.n7026 vdd.n7025 61.358
R37896 vdd.n7193 vdd.n7190 61.358
R37897 vdd.n7193 vdd.n7192 61.358
R37898 vdd.n7342 vdd.n7339 61.358
R37899 vdd.n7342 vdd.n7341 61.358
R37900 vdd.n7334 vdd.n7331 61.358
R37901 vdd.n7334 vdd.n7333 61.358
R37902 vdd.n7326 vdd.n7323 61.358
R37903 vdd.n7326 vdd.n7325 61.358
R37904 vdd.n7318 vdd.n7315 61.358
R37905 vdd.n7318 vdd.n7317 61.358
R37906 vdd.n7310 vdd.n7307 61.358
R37907 vdd.n7310 vdd.n7309 61.358
R37908 vdd.n7302 vdd.n7299 61.358
R37909 vdd.n7302 vdd.n7301 61.358
R37910 vdd.n7294 vdd.n7291 61.358
R37911 vdd.n7294 vdd.n7293 61.358
R37912 vdd.n7286 vdd.n7283 61.358
R37913 vdd.n7286 vdd.n7285 61.358
R37914 vdd.n7278 vdd.n7275 61.358
R37915 vdd.n7278 vdd.n7277 61.358
R37916 vdd.n7262 vdd.n7259 61.358
R37917 vdd.n7262 vdd.n7261 61.358
R37918 vdd.n7254 vdd.n7251 61.358
R37919 vdd.n7254 vdd.n7253 61.358
R37920 vdd.n7246 vdd.n7243 61.358
R37921 vdd.n7246 vdd.n7245 61.358
R37922 vdd.n7238 vdd.n7235 61.358
R37923 vdd.n7238 vdd.n7237 61.358
R37924 vdd.n7230 vdd.n7227 61.358
R37925 vdd.n7230 vdd.n7229 61.358
R37926 vdd.n7222 vdd.n7219 61.358
R37927 vdd.n7222 vdd.n7221 61.358
R37928 vdd.n7214 vdd.n7211 61.358
R37929 vdd.n7214 vdd.n7213 61.358
R37930 vdd.n7206 vdd.n7203 61.358
R37931 vdd.n7206 vdd.n7205 61.358
R37932 vdd.n7373 vdd.n7370 61.358
R37933 vdd.n7373 vdd.n7372 61.358
R37934 vdd.n7522 vdd.n7519 61.358
R37935 vdd.n7522 vdd.n7521 61.358
R37936 vdd.n7514 vdd.n7511 61.358
R37937 vdd.n7514 vdd.n7513 61.358
R37938 vdd.n7506 vdd.n7503 61.358
R37939 vdd.n7506 vdd.n7505 61.358
R37940 vdd.n7498 vdd.n7495 61.358
R37941 vdd.n7498 vdd.n7497 61.358
R37942 vdd.n7490 vdd.n7487 61.358
R37943 vdd.n7490 vdd.n7489 61.358
R37944 vdd.n7482 vdd.n7479 61.358
R37945 vdd.n7482 vdd.n7481 61.358
R37946 vdd.n7474 vdd.n7471 61.358
R37947 vdd.n7474 vdd.n7473 61.358
R37948 vdd.n7466 vdd.n7463 61.358
R37949 vdd.n7466 vdd.n7465 61.358
R37950 vdd.n7458 vdd.n7455 61.358
R37951 vdd.n7458 vdd.n7457 61.358
R37952 vdd.n7442 vdd.n7439 61.358
R37953 vdd.n7442 vdd.n7441 61.358
R37954 vdd.n7434 vdd.n7431 61.358
R37955 vdd.n7434 vdd.n7433 61.358
R37956 vdd.n7426 vdd.n7423 61.358
R37957 vdd.n7426 vdd.n7425 61.358
R37958 vdd.n7418 vdd.n7415 61.358
R37959 vdd.n7418 vdd.n7417 61.358
R37960 vdd.n7410 vdd.n7407 61.358
R37961 vdd.n7410 vdd.n7409 61.358
R37962 vdd.n7402 vdd.n7399 61.358
R37963 vdd.n7402 vdd.n7401 61.358
R37964 vdd.n7394 vdd.n7391 61.358
R37965 vdd.n7394 vdd.n7393 61.358
R37966 vdd.n7386 vdd.n7383 61.358
R37967 vdd.n7386 vdd.n7385 61.358
R37968 vdd.n7553 vdd.n7550 61.358
R37969 vdd.n7553 vdd.n7552 61.358
R37970 vdd.n7702 vdd.n7699 61.358
R37971 vdd.n7702 vdd.n7701 61.358
R37972 vdd.n7694 vdd.n7691 61.358
R37973 vdd.n7694 vdd.n7693 61.358
R37974 vdd.n7686 vdd.n7683 61.358
R37975 vdd.n7686 vdd.n7685 61.358
R37976 vdd.n7678 vdd.n7675 61.358
R37977 vdd.n7678 vdd.n7677 61.358
R37978 vdd.n7670 vdd.n7667 61.358
R37979 vdd.n7670 vdd.n7669 61.358
R37980 vdd.n7662 vdd.n7659 61.358
R37981 vdd.n7662 vdd.n7661 61.358
R37982 vdd.n7654 vdd.n7651 61.358
R37983 vdd.n7654 vdd.n7653 61.358
R37984 vdd.n7646 vdd.n7643 61.358
R37985 vdd.n7646 vdd.n7645 61.358
R37986 vdd.n7638 vdd.n7635 61.358
R37987 vdd.n7638 vdd.n7637 61.358
R37988 vdd.n7622 vdd.n7619 61.358
R37989 vdd.n7622 vdd.n7621 61.358
R37990 vdd.n7614 vdd.n7611 61.358
R37991 vdd.n7614 vdd.n7613 61.358
R37992 vdd.n7606 vdd.n7603 61.358
R37993 vdd.n7606 vdd.n7605 61.358
R37994 vdd.n7598 vdd.n7595 61.358
R37995 vdd.n7598 vdd.n7597 61.358
R37996 vdd.n7590 vdd.n7587 61.358
R37997 vdd.n7590 vdd.n7589 61.358
R37998 vdd.n7582 vdd.n7579 61.358
R37999 vdd.n7582 vdd.n7581 61.358
R38000 vdd.n7574 vdd.n7571 61.358
R38001 vdd.n7574 vdd.n7573 61.358
R38002 vdd.n7566 vdd.n7563 61.358
R38003 vdd.n7566 vdd.n7565 61.358
R38004 vdd.n7733 vdd.n7730 61.358
R38005 vdd.n7733 vdd.n7732 61.358
R38006 vdd.n7882 vdd.n7879 61.358
R38007 vdd.n7882 vdd.n7881 61.358
R38008 vdd.n7874 vdd.n7871 61.358
R38009 vdd.n7874 vdd.n7873 61.358
R38010 vdd.n7866 vdd.n7863 61.358
R38011 vdd.n7866 vdd.n7865 61.358
R38012 vdd.n7858 vdd.n7855 61.358
R38013 vdd.n7858 vdd.n7857 61.358
R38014 vdd.n7850 vdd.n7847 61.358
R38015 vdd.n7850 vdd.n7849 61.358
R38016 vdd.n7842 vdd.n7839 61.358
R38017 vdd.n7842 vdd.n7841 61.358
R38018 vdd.n7834 vdd.n7831 61.358
R38019 vdd.n7834 vdd.n7833 61.358
R38020 vdd.n7826 vdd.n7823 61.358
R38021 vdd.n7826 vdd.n7825 61.358
R38022 vdd.n7818 vdd.n7815 61.358
R38023 vdd.n7818 vdd.n7817 61.358
R38024 vdd.n7802 vdd.n7799 61.358
R38025 vdd.n7802 vdd.n7801 61.358
R38026 vdd.n7794 vdd.n7791 61.358
R38027 vdd.n7794 vdd.n7793 61.358
R38028 vdd.n7786 vdd.n7783 61.358
R38029 vdd.n7786 vdd.n7785 61.358
R38030 vdd.n7778 vdd.n7775 61.358
R38031 vdd.n7778 vdd.n7777 61.358
R38032 vdd.n7770 vdd.n7767 61.358
R38033 vdd.n7770 vdd.n7769 61.358
R38034 vdd.n7762 vdd.n7759 61.358
R38035 vdd.n7762 vdd.n7761 61.358
R38036 vdd.n7754 vdd.n7751 61.358
R38037 vdd.n7754 vdd.n7753 61.358
R38038 vdd.n7746 vdd.n7743 61.358
R38039 vdd.n7746 vdd.n7745 61.358
R38040 vdd.n7913 vdd.n7910 61.358
R38041 vdd.n7913 vdd.n7912 61.358
R38042 vdd.n8062 vdd.n8059 61.358
R38043 vdd.n8062 vdd.n8061 61.358
R38044 vdd.n8054 vdd.n8051 61.358
R38045 vdd.n8054 vdd.n8053 61.358
R38046 vdd.n8046 vdd.n8043 61.358
R38047 vdd.n8046 vdd.n8045 61.358
R38048 vdd.n8038 vdd.n8035 61.358
R38049 vdd.n8038 vdd.n8037 61.358
R38050 vdd.n8030 vdd.n8027 61.358
R38051 vdd.n8030 vdd.n8029 61.358
R38052 vdd.n8022 vdd.n8019 61.358
R38053 vdd.n8022 vdd.n8021 61.358
R38054 vdd.n8014 vdd.n8011 61.358
R38055 vdd.n8014 vdd.n8013 61.358
R38056 vdd.n8006 vdd.n8003 61.358
R38057 vdd.n8006 vdd.n8005 61.358
R38058 vdd.n7998 vdd.n7995 61.358
R38059 vdd.n7998 vdd.n7997 61.358
R38060 vdd.n7982 vdd.n7979 61.358
R38061 vdd.n7982 vdd.n7981 61.358
R38062 vdd.n7974 vdd.n7971 61.358
R38063 vdd.n7974 vdd.n7973 61.358
R38064 vdd.n7966 vdd.n7963 61.358
R38065 vdd.n7966 vdd.n7965 61.358
R38066 vdd.n7958 vdd.n7955 61.358
R38067 vdd.n7958 vdd.n7957 61.358
R38068 vdd.n7950 vdd.n7947 61.358
R38069 vdd.n7950 vdd.n7949 61.358
R38070 vdd.n7942 vdd.n7939 61.358
R38071 vdd.n7942 vdd.n7941 61.358
R38072 vdd.n7934 vdd.n7931 61.358
R38073 vdd.n7934 vdd.n7933 61.358
R38074 vdd.n7926 vdd.n7923 61.358
R38075 vdd.n7926 vdd.n7925 61.358
R38076 vdd.n8093 vdd.n8090 61.358
R38077 vdd.n8093 vdd.n8092 61.358
R38078 vdd.n8242 vdd.n8239 61.358
R38079 vdd.n8242 vdd.n8241 61.358
R38080 vdd.n8234 vdd.n8231 61.358
R38081 vdd.n8234 vdd.n8233 61.358
R38082 vdd.n8226 vdd.n8223 61.358
R38083 vdd.n8226 vdd.n8225 61.358
R38084 vdd.n8218 vdd.n8215 61.358
R38085 vdd.n8218 vdd.n8217 61.358
R38086 vdd.n8210 vdd.n8207 61.358
R38087 vdd.n8210 vdd.n8209 61.358
R38088 vdd.n8202 vdd.n8199 61.358
R38089 vdd.n8202 vdd.n8201 61.358
R38090 vdd.n8194 vdd.n8191 61.358
R38091 vdd.n8194 vdd.n8193 61.358
R38092 vdd.n8186 vdd.n8183 61.358
R38093 vdd.n8186 vdd.n8185 61.358
R38094 vdd.n8178 vdd.n8175 61.358
R38095 vdd.n8178 vdd.n8177 61.358
R38096 vdd.n8162 vdd.n8159 61.358
R38097 vdd.n8162 vdd.n8161 61.358
R38098 vdd.n8154 vdd.n8151 61.358
R38099 vdd.n8154 vdd.n8153 61.358
R38100 vdd.n8146 vdd.n8143 61.358
R38101 vdd.n8146 vdd.n8145 61.358
R38102 vdd.n8138 vdd.n8135 61.358
R38103 vdd.n8138 vdd.n8137 61.358
R38104 vdd.n8130 vdd.n8127 61.358
R38105 vdd.n8130 vdd.n8129 61.358
R38106 vdd.n8122 vdd.n8119 61.358
R38107 vdd.n8122 vdd.n8121 61.358
R38108 vdd.n8114 vdd.n8111 61.358
R38109 vdd.n8114 vdd.n8113 61.358
R38110 vdd.n8106 vdd.n8103 61.358
R38111 vdd.n8106 vdd.n8105 61.358
R38112 vdd.n8273 vdd.n8270 61.358
R38113 vdd.n8273 vdd.n8272 61.358
R38114 vdd.n8422 vdd.n8419 61.358
R38115 vdd.n8422 vdd.n8421 61.358
R38116 vdd.n8414 vdd.n8411 61.358
R38117 vdd.n8414 vdd.n8413 61.358
R38118 vdd.n8406 vdd.n8403 61.358
R38119 vdd.n8406 vdd.n8405 61.358
R38120 vdd.n8398 vdd.n8395 61.358
R38121 vdd.n8398 vdd.n8397 61.358
R38122 vdd.n8390 vdd.n8387 61.358
R38123 vdd.n8390 vdd.n8389 61.358
R38124 vdd.n8382 vdd.n8379 61.358
R38125 vdd.n8382 vdd.n8381 61.358
R38126 vdd.n8374 vdd.n8371 61.358
R38127 vdd.n8374 vdd.n8373 61.358
R38128 vdd.n8366 vdd.n8363 61.358
R38129 vdd.n8366 vdd.n8365 61.358
R38130 vdd.n8358 vdd.n8355 61.358
R38131 vdd.n8358 vdd.n8357 61.358
R38132 vdd.n8342 vdd.n8339 61.358
R38133 vdd.n8342 vdd.n8341 61.358
R38134 vdd.n8334 vdd.n8331 61.358
R38135 vdd.n8334 vdd.n8333 61.358
R38136 vdd.n8326 vdd.n8323 61.358
R38137 vdd.n8326 vdd.n8325 61.358
R38138 vdd.n8318 vdd.n8315 61.358
R38139 vdd.n8318 vdd.n8317 61.358
R38140 vdd.n8310 vdd.n8307 61.358
R38141 vdd.n8310 vdd.n8309 61.358
R38142 vdd.n8302 vdd.n8299 61.358
R38143 vdd.n8302 vdd.n8301 61.358
R38144 vdd.n8294 vdd.n8291 61.358
R38145 vdd.n8294 vdd.n8293 61.358
R38146 vdd.n8286 vdd.n8283 61.358
R38147 vdd.n8286 vdd.n8285 61.358
R38148 vdd.n8453 vdd.n8450 61.358
R38149 vdd.n8453 vdd.n8452 61.358
R38150 vdd.n8602 vdd.n8599 61.358
R38151 vdd.n8602 vdd.n8601 61.358
R38152 vdd.n8594 vdd.n8591 61.358
R38153 vdd.n8594 vdd.n8593 61.358
R38154 vdd.n8586 vdd.n8583 61.358
R38155 vdd.n8586 vdd.n8585 61.358
R38156 vdd.n8578 vdd.n8575 61.358
R38157 vdd.n8578 vdd.n8577 61.358
R38158 vdd.n8570 vdd.n8567 61.358
R38159 vdd.n8570 vdd.n8569 61.358
R38160 vdd.n8562 vdd.n8559 61.358
R38161 vdd.n8562 vdd.n8561 61.358
R38162 vdd.n8554 vdd.n8551 61.358
R38163 vdd.n8554 vdd.n8553 61.358
R38164 vdd.n8546 vdd.n8543 61.358
R38165 vdd.n8546 vdd.n8545 61.358
R38166 vdd.n8538 vdd.n8535 61.358
R38167 vdd.n8538 vdd.n8537 61.358
R38168 vdd.n8522 vdd.n8519 61.358
R38169 vdd.n8522 vdd.n8521 61.358
R38170 vdd.n8514 vdd.n8511 61.358
R38171 vdd.n8514 vdd.n8513 61.358
R38172 vdd.n8506 vdd.n8503 61.358
R38173 vdd.n8506 vdd.n8505 61.358
R38174 vdd.n8498 vdd.n8495 61.358
R38175 vdd.n8498 vdd.n8497 61.358
R38176 vdd.n8490 vdd.n8487 61.358
R38177 vdd.n8490 vdd.n8489 61.358
R38178 vdd.n8482 vdd.n8479 61.358
R38179 vdd.n8482 vdd.n8481 61.358
R38180 vdd.n8474 vdd.n8471 61.358
R38181 vdd.n8474 vdd.n8473 61.358
R38182 vdd.n8466 vdd.n8463 61.358
R38183 vdd.n8466 vdd.n8465 61.358
R38184 vdd.n8633 vdd.n8630 61.358
R38185 vdd.n8633 vdd.n8632 61.358
R38186 vdd.n8782 vdd.n8779 61.358
R38187 vdd.n8782 vdd.n8781 61.358
R38188 vdd.n8774 vdd.n8771 61.358
R38189 vdd.n8774 vdd.n8773 61.358
R38190 vdd.n8766 vdd.n8763 61.358
R38191 vdd.n8766 vdd.n8765 61.358
R38192 vdd.n8758 vdd.n8755 61.358
R38193 vdd.n8758 vdd.n8757 61.358
R38194 vdd.n8750 vdd.n8747 61.358
R38195 vdd.n8750 vdd.n8749 61.358
R38196 vdd.n8742 vdd.n8739 61.358
R38197 vdd.n8742 vdd.n8741 61.358
R38198 vdd.n8734 vdd.n8731 61.358
R38199 vdd.n8734 vdd.n8733 61.358
R38200 vdd.n8726 vdd.n8723 61.358
R38201 vdd.n8726 vdd.n8725 61.358
R38202 vdd.n8718 vdd.n8715 61.358
R38203 vdd.n8718 vdd.n8717 61.358
R38204 vdd.n8702 vdd.n8699 61.358
R38205 vdd.n8702 vdd.n8701 61.358
R38206 vdd.n8694 vdd.n8691 61.358
R38207 vdd.n8694 vdd.n8693 61.358
R38208 vdd.n8686 vdd.n8683 61.358
R38209 vdd.n8686 vdd.n8685 61.358
R38210 vdd.n8678 vdd.n8675 61.358
R38211 vdd.n8678 vdd.n8677 61.358
R38212 vdd.n8670 vdd.n8667 61.358
R38213 vdd.n8670 vdd.n8669 61.358
R38214 vdd.n8662 vdd.n8659 61.358
R38215 vdd.n8662 vdd.n8661 61.358
R38216 vdd.n8654 vdd.n8651 61.358
R38217 vdd.n8654 vdd.n8653 61.358
R38218 vdd.n8646 vdd.n8643 61.358
R38219 vdd.n8646 vdd.n8645 61.358
R38220 vdd.n8813 vdd.n8810 61.358
R38221 vdd.n8813 vdd.n8812 61.358
R38222 vdd.n8962 vdd.n8959 61.358
R38223 vdd.n8962 vdd.n8961 61.358
R38224 vdd.n8954 vdd.n8951 61.358
R38225 vdd.n8954 vdd.n8953 61.358
R38226 vdd.n8946 vdd.n8943 61.358
R38227 vdd.n8946 vdd.n8945 61.358
R38228 vdd.n8938 vdd.n8935 61.358
R38229 vdd.n8938 vdd.n8937 61.358
R38230 vdd.n8930 vdd.n8927 61.358
R38231 vdd.n8930 vdd.n8929 61.358
R38232 vdd.n8922 vdd.n8919 61.358
R38233 vdd.n8922 vdd.n8921 61.358
R38234 vdd.n8914 vdd.n8911 61.358
R38235 vdd.n8914 vdd.n8913 61.358
R38236 vdd.n8906 vdd.n8903 61.358
R38237 vdd.n8906 vdd.n8905 61.358
R38238 vdd.n8898 vdd.n8895 61.358
R38239 vdd.n8898 vdd.n8897 61.358
R38240 vdd.n8882 vdd.n8879 61.358
R38241 vdd.n8882 vdd.n8881 61.358
R38242 vdd.n8874 vdd.n8871 61.358
R38243 vdd.n8874 vdd.n8873 61.358
R38244 vdd.n8866 vdd.n8863 61.358
R38245 vdd.n8866 vdd.n8865 61.358
R38246 vdd.n8858 vdd.n8855 61.358
R38247 vdd.n8858 vdd.n8857 61.358
R38248 vdd.n8850 vdd.n8847 61.358
R38249 vdd.n8850 vdd.n8849 61.358
R38250 vdd.n8842 vdd.n8839 61.358
R38251 vdd.n8842 vdd.n8841 61.358
R38252 vdd.n8834 vdd.n8831 61.358
R38253 vdd.n8834 vdd.n8833 61.358
R38254 vdd.n8826 vdd.n8823 61.358
R38255 vdd.n8826 vdd.n8825 61.358
R38256 vdd.n8993 vdd.n8990 61.358
R38257 vdd.n8993 vdd.n8992 61.358
R38258 vdd.n9142 vdd.n9139 61.358
R38259 vdd.n9142 vdd.n9141 61.358
R38260 vdd.n9134 vdd.n9131 61.358
R38261 vdd.n9134 vdd.n9133 61.358
R38262 vdd.n9126 vdd.n9123 61.358
R38263 vdd.n9126 vdd.n9125 61.358
R38264 vdd.n9118 vdd.n9115 61.358
R38265 vdd.n9118 vdd.n9117 61.358
R38266 vdd.n9110 vdd.n9107 61.358
R38267 vdd.n9110 vdd.n9109 61.358
R38268 vdd.n9102 vdd.n9099 61.358
R38269 vdd.n9102 vdd.n9101 61.358
R38270 vdd.n9094 vdd.n9091 61.358
R38271 vdd.n9094 vdd.n9093 61.358
R38272 vdd.n9086 vdd.n9083 61.358
R38273 vdd.n9086 vdd.n9085 61.358
R38274 vdd.n9078 vdd.n9075 61.358
R38275 vdd.n9078 vdd.n9077 61.358
R38276 vdd.n9062 vdd.n9059 61.358
R38277 vdd.n9062 vdd.n9061 61.358
R38278 vdd.n9054 vdd.n9051 61.358
R38279 vdd.n9054 vdd.n9053 61.358
R38280 vdd.n9046 vdd.n9043 61.358
R38281 vdd.n9046 vdd.n9045 61.358
R38282 vdd.n9038 vdd.n9035 61.358
R38283 vdd.n9038 vdd.n9037 61.358
R38284 vdd.n9030 vdd.n9027 61.358
R38285 vdd.n9030 vdd.n9029 61.358
R38286 vdd.n9022 vdd.n9019 61.358
R38287 vdd.n9022 vdd.n9021 61.358
R38288 vdd.n9014 vdd.n9011 61.358
R38289 vdd.n9014 vdd.n9013 61.358
R38290 vdd.n9006 vdd.n9003 61.358
R38291 vdd.n9006 vdd.n9005 61.358
R38292 vdd.n9173 vdd.n9170 61.358
R38293 vdd.n9173 vdd.n9172 61.358
R38294 vdd.n9322 vdd.n9319 61.358
R38295 vdd.n9322 vdd.n9321 61.358
R38296 vdd.n9314 vdd.n9311 61.358
R38297 vdd.n9314 vdd.n9313 61.358
R38298 vdd.n9306 vdd.n9303 61.358
R38299 vdd.n9306 vdd.n9305 61.358
R38300 vdd.n9298 vdd.n9295 61.358
R38301 vdd.n9298 vdd.n9297 61.358
R38302 vdd.n9290 vdd.n9287 61.358
R38303 vdd.n9290 vdd.n9289 61.358
R38304 vdd.n9282 vdd.n9279 61.358
R38305 vdd.n9282 vdd.n9281 61.358
R38306 vdd.n9274 vdd.n9271 61.358
R38307 vdd.n9274 vdd.n9273 61.358
R38308 vdd.n9266 vdd.n9263 61.358
R38309 vdd.n9266 vdd.n9265 61.358
R38310 vdd.n9258 vdd.n9255 61.358
R38311 vdd.n9258 vdd.n9257 61.358
R38312 vdd.n9242 vdd.n9239 61.358
R38313 vdd.n9242 vdd.n9241 61.358
R38314 vdd.n9234 vdd.n9231 61.358
R38315 vdd.n9234 vdd.n9233 61.358
R38316 vdd.n9226 vdd.n9223 61.358
R38317 vdd.n9226 vdd.n9225 61.358
R38318 vdd.n9218 vdd.n9215 61.358
R38319 vdd.n9218 vdd.n9217 61.358
R38320 vdd.n9210 vdd.n9207 61.358
R38321 vdd.n9210 vdd.n9209 61.358
R38322 vdd.n9202 vdd.n9199 61.358
R38323 vdd.n9202 vdd.n9201 61.358
R38324 vdd.n9194 vdd.n9191 61.358
R38325 vdd.n9194 vdd.n9193 61.358
R38326 vdd.n9186 vdd.n9183 61.358
R38327 vdd.n9186 vdd.n9185 61.358
R38328 vdd.n9353 vdd.n9350 61.358
R38329 vdd.n9353 vdd.n9352 61.358
R38330 vdd.n9502 vdd.n9499 61.358
R38331 vdd.n9502 vdd.n9501 61.358
R38332 vdd.n9494 vdd.n9491 61.358
R38333 vdd.n9494 vdd.n9493 61.358
R38334 vdd.n9486 vdd.n9483 61.358
R38335 vdd.n9486 vdd.n9485 61.358
R38336 vdd.n9478 vdd.n9475 61.358
R38337 vdd.n9478 vdd.n9477 61.358
R38338 vdd.n9470 vdd.n9467 61.358
R38339 vdd.n9470 vdd.n9469 61.358
R38340 vdd.n9462 vdd.n9459 61.358
R38341 vdd.n9462 vdd.n9461 61.358
R38342 vdd.n9454 vdd.n9451 61.358
R38343 vdd.n9454 vdd.n9453 61.358
R38344 vdd.n9446 vdd.n9443 61.358
R38345 vdd.n9446 vdd.n9445 61.358
R38346 vdd.n9438 vdd.n9435 61.358
R38347 vdd.n9438 vdd.n9437 61.358
R38348 vdd.n9422 vdd.n9419 61.358
R38349 vdd.n9422 vdd.n9421 61.358
R38350 vdd.n9414 vdd.n9411 61.358
R38351 vdd.n9414 vdd.n9413 61.358
R38352 vdd.n9406 vdd.n9403 61.358
R38353 vdd.n9406 vdd.n9405 61.358
R38354 vdd.n9398 vdd.n9395 61.358
R38355 vdd.n9398 vdd.n9397 61.358
R38356 vdd.n9390 vdd.n9387 61.358
R38357 vdd.n9390 vdd.n9389 61.358
R38358 vdd.n9382 vdd.n9379 61.358
R38359 vdd.n9382 vdd.n9381 61.358
R38360 vdd.n9374 vdd.n9371 61.358
R38361 vdd.n9374 vdd.n9373 61.358
R38362 vdd.n9366 vdd.n9363 61.358
R38363 vdd.n9366 vdd.n9365 61.358
R38364 vdd.n9533 vdd.n9530 61.358
R38365 vdd.n9533 vdd.n9532 61.358
R38366 vdd.n9682 vdd.n9679 61.358
R38367 vdd.n9682 vdd.n9681 61.358
R38368 vdd.n9674 vdd.n9671 61.358
R38369 vdd.n9674 vdd.n9673 61.358
R38370 vdd.n9666 vdd.n9663 61.358
R38371 vdd.n9666 vdd.n9665 61.358
R38372 vdd.n9658 vdd.n9655 61.358
R38373 vdd.n9658 vdd.n9657 61.358
R38374 vdd.n9650 vdd.n9647 61.358
R38375 vdd.n9650 vdd.n9649 61.358
R38376 vdd.n9642 vdd.n9639 61.358
R38377 vdd.n9642 vdd.n9641 61.358
R38378 vdd.n9634 vdd.n9631 61.358
R38379 vdd.n9634 vdd.n9633 61.358
R38380 vdd.n9626 vdd.n9623 61.358
R38381 vdd.n9626 vdd.n9625 61.358
R38382 vdd.n9618 vdd.n9615 61.358
R38383 vdd.n9618 vdd.n9617 61.358
R38384 vdd.n9602 vdd.n9599 61.358
R38385 vdd.n9602 vdd.n9601 61.358
R38386 vdd.n9594 vdd.n9591 61.358
R38387 vdd.n9594 vdd.n9593 61.358
R38388 vdd.n9586 vdd.n9583 61.358
R38389 vdd.n9586 vdd.n9585 61.358
R38390 vdd.n9578 vdd.n9575 61.358
R38391 vdd.n9578 vdd.n9577 61.358
R38392 vdd.n9570 vdd.n9567 61.358
R38393 vdd.n9570 vdd.n9569 61.358
R38394 vdd.n9562 vdd.n9559 61.358
R38395 vdd.n9562 vdd.n9561 61.358
R38396 vdd.n9554 vdd.n9551 61.358
R38397 vdd.n9554 vdd.n9553 61.358
R38398 vdd.n9546 vdd.n9543 61.358
R38399 vdd.n9546 vdd.n9545 61.358
R38400 vdd.n9713 vdd.n9710 61.358
R38401 vdd.n9713 vdd.n9712 61.358
R38402 vdd.n9862 vdd.n9859 61.358
R38403 vdd.n9862 vdd.n9861 61.358
R38404 vdd.n9854 vdd.n9851 61.358
R38405 vdd.n9854 vdd.n9853 61.358
R38406 vdd.n9846 vdd.n9843 61.358
R38407 vdd.n9846 vdd.n9845 61.358
R38408 vdd.n9838 vdd.n9835 61.358
R38409 vdd.n9838 vdd.n9837 61.358
R38410 vdd.n9830 vdd.n9827 61.358
R38411 vdd.n9830 vdd.n9829 61.358
R38412 vdd.n9822 vdd.n9819 61.358
R38413 vdd.n9822 vdd.n9821 61.358
R38414 vdd.n9814 vdd.n9811 61.358
R38415 vdd.n9814 vdd.n9813 61.358
R38416 vdd.n9806 vdd.n9803 61.358
R38417 vdd.n9806 vdd.n9805 61.358
R38418 vdd.n9798 vdd.n9795 61.358
R38419 vdd.n9798 vdd.n9797 61.358
R38420 vdd.n9782 vdd.n9779 61.358
R38421 vdd.n9782 vdd.n9781 61.358
R38422 vdd.n9774 vdd.n9771 61.358
R38423 vdd.n9774 vdd.n9773 61.358
R38424 vdd.n9766 vdd.n9763 61.358
R38425 vdd.n9766 vdd.n9765 61.358
R38426 vdd.n9758 vdd.n9755 61.358
R38427 vdd.n9758 vdd.n9757 61.358
R38428 vdd.n9750 vdd.n9747 61.358
R38429 vdd.n9750 vdd.n9749 61.358
R38430 vdd.n9742 vdd.n9739 61.358
R38431 vdd.n9742 vdd.n9741 61.358
R38432 vdd.n9734 vdd.n9731 61.358
R38433 vdd.n9734 vdd.n9733 61.358
R38434 vdd.n9726 vdd.n9723 61.358
R38435 vdd.n9726 vdd.n9725 61.358
R38436 vdd.n9893 vdd.n9890 61.358
R38437 vdd.n9893 vdd.n9892 61.358
R38438 vdd.n10042 vdd.n10039 61.358
R38439 vdd.n10042 vdd.n10041 61.358
R38440 vdd.n10034 vdd.n10031 61.358
R38441 vdd.n10034 vdd.n10033 61.358
R38442 vdd.n10026 vdd.n10023 61.358
R38443 vdd.n10026 vdd.n10025 61.358
R38444 vdd.n10018 vdd.n10015 61.358
R38445 vdd.n10018 vdd.n10017 61.358
R38446 vdd.n10010 vdd.n10007 61.358
R38447 vdd.n10010 vdd.n10009 61.358
R38448 vdd.n10002 vdd.n9999 61.358
R38449 vdd.n10002 vdd.n10001 61.358
R38450 vdd.n9994 vdd.n9991 61.358
R38451 vdd.n9994 vdd.n9993 61.358
R38452 vdd.n9986 vdd.n9983 61.358
R38453 vdd.n9986 vdd.n9985 61.358
R38454 vdd.n9978 vdd.n9975 61.358
R38455 vdd.n9978 vdd.n9977 61.358
R38456 vdd.n9962 vdd.n9959 61.358
R38457 vdd.n9962 vdd.n9961 61.358
R38458 vdd.n9954 vdd.n9951 61.358
R38459 vdd.n9954 vdd.n9953 61.358
R38460 vdd.n9946 vdd.n9943 61.358
R38461 vdd.n9946 vdd.n9945 61.358
R38462 vdd.n9938 vdd.n9935 61.358
R38463 vdd.n9938 vdd.n9937 61.358
R38464 vdd.n9930 vdd.n9927 61.358
R38465 vdd.n9930 vdd.n9929 61.358
R38466 vdd.n9922 vdd.n9919 61.358
R38467 vdd.n9922 vdd.n9921 61.358
R38468 vdd.n9914 vdd.n9911 61.358
R38469 vdd.n9914 vdd.n9913 61.358
R38470 vdd.n9906 vdd.n9903 61.358
R38471 vdd.n9906 vdd.n9905 61.358
R38472 vdd.n10073 vdd.n10070 61.358
R38473 vdd.n10073 vdd.n10072 61.358
R38474 vdd.n10222 vdd.n10219 61.358
R38475 vdd.n10222 vdd.n10221 61.358
R38476 vdd.n10214 vdd.n10211 61.358
R38477 vdd.n10214 vdd.n10213 61.358
R38478 vdd.n10206 vdd.n10203 61.358
R38479 vdd.n10206 vdd.n10205 61.358
R38480 vdd.n10198 vdd.n10195 61.358
R38481 vdd.n10198 vdd.n10197 61.358
R38482 vdd.n10190 vdd.n10187 61.358
R38483 vdd.n10190 vdd.n10189 61.358
R38484 vdd.n10182 vdd.n10179 61.358
R38485 vdd.n10182 vdd.n10181 61.358
R38486 vdd.n10174 vdd.n10171 61.358
R38487 vdd.n10174 vdd.n10173 61.358
R38488 vdd.n10166 vdd.n10163 61.358
R38489 vdd.n10166 vdd.n10165 61.358
R38490 vdd.n10158 vdd.n10155 61.358
R38491 vdd.n10158 vdd.n10157 61.358
R38492 vdd.n10142 vdd.n10139 61.358
R38493 vdd.n10142 vdd.n10141 61.358
R38494 vdd.n10134 vdd.n10131 61.358
R38495 vdd.n10134 vdd.n10133 61.358
R38496 vdd.n10126 vdd.n10123 61.358
R38497 vdd.n10126 vdd.n10125 61.358
R38498 vdd.n10118 vdd.n10115 61.358
R38499 vdd.n10118 vdd.n10117 61.358
R38500 vdd.n10110 vdd.n10107 61.358
R38501 vdd.n10110 vdd.n10109 61.358
R38502 vdd.n10102 vdd.n10099 61.358
R38503 vdd.n10102 vdd.n10101 61.358
R38504 vdd.n10094 vdd.n10091 61.358
R38505 vdd.n10094 vdd.n10093 61.358
R38506 vdd.n10086 vdd.n10083 61.358
R38507 vdd.n10086 vdd.n10085 61.358
R38508 vdd.n10253 vdd.n10250 61.358
R38509 vdd.n10253 vdd.n10252 61.358
R38510 vdd.n10402 vdd.n10399 61.358
R38511 vdd.n10402 vdd.n10401 61.358
R38512 vdd.n10394 vdd.n10391 61.358
R38513 vdd.n10394 vdd.n10393 61.358
R38514 vdd.n10386 vdd.n10383 61.358
R38515 vdd.n10386 vdd.n10385 61.358
R38516 vdd.n10378 vdd.n10375 61.358
R38517 vdd.n10378 vdd.n10377 61.358
R38518 vdd.n10370 vdd.n10367 61.358
R38519 vdd.n10370 vdd.n10369 61.358
R38520 vdd.n10362 vdd.n10359 61.358
R38521 vdd.n10362 vdd.n10361 61.358
R38522 vdd.n10354 vdd.n10351 61.358
R38523 vdd.n10354 vdd.n10353 61.358
R38524 vdd.n10346 vdd.n10343 61.358
R38525 vdd.n10346 vdd.n10345 61.358
R38526 vdd.n10338 vdd.n10335 61.358
R38527 vdd.n10338 vdd.n10337 61.358
R38528 vdd.n10322 vdd.n10319 61.358
R38529 vdd.n10322 vdd.n10321 61.358
R38530 vdd.n10314 vdd.n10311 61.358
R38531 vdd.n10314 vdd.n10313 61.358
R38532 vdd.n10306 vdd.n10303 61.358
R38533 vdd.n10306 vdd.n10305 61.358
R38534 vdd.n10298 vdd.n10295 61.358
R38535 vdd.n10298 vdd.n10297 61.358
R38536 vdd.n10290 vdd.n10287 61.358
R38537 vdd.n10290 vdd.n10289 61.358
R38538 vdd.n10282 vdd.n10279 61.358
R38539 vdd.n10282 vdd.n10281 61.358
R38540 vdd.n10274 vdd.n10271 61.358
R38541 vdd.n10274 vdd.n10273 61.358
R38542 vdd.n10266 vdd.n10263 61.358
R38543 vdd.n10266 vdd.n10265 61.358
R38544 vdd.n10433 vdd.n10430 61.358
R38545 vdd.n10433 vdd.n10432 61.358
R38546 vdd.n10582 vdd.n10579 61.358
R38547 vdd.n10582 vdd.n10581 61.358
R38548 vdd.n10574 vdd.n10571 61.358
R38549 vdd.n10574 vdd.n10573 61.358
R38550 vdd.n10566 vdd.n10563 61.358
R38551 vdd.n10566 vdd.n10565 61.358
R38552 vdd.n10558 vdd.n10555 61.358
R38553 vdd.n10558 vdd.n10557 61.358
R38554 vdd.n10550 vdd.n10547 61.358
R38555 vdd.n10550 vdd.n10549 61.358
R38556 vdd.n10542 vdd.n10539 61.358
R38557 vdd.n10542 vdd.n10541 61.358
R38558 vdd.n10534 vdd.n10531 61.358
R38559 vdd.n10534 vdd.n10533 61.358
R38560 vdd.n10526 vdd.n10523 61.358
R38561 vdd.n10526 vdd.n10525 61.358
R38562 vdd.n10518 vdd.n10515 61.358
R38563 vdd.n10518 vdd.n10517 61.358
R38564 vdd.n10502 vdd.n10499 61.358
R38565 vdd.n10502 vdd.n10501 61.358
R38566 vdd.n10494 vdd.n10491 61.358
R38567 vdd.n10494 vdd.n10493 61.358
R38568 vdd.n10486 vdd.n10483 61.358
R38569 vdd.n10486 vdd.n10485 61.358
R38570 vdd.n10478 vdd.n10475 61.358
R38571 vdd.n10478 vdd.n10477 61.358
R38572 vdd.n10470 vdd.n10467 61.358
R38573 vdd.n10470 vdd.n10469 61.358
R38574 vdd.n10462 vdd.n10459 61.358
R38575 vdd.n10462 vdd.n10461 61.358
R38576 vdd.n10454 vdd.n10451 61.358
R38577 vdd.n10454 vdd.n10453 61.358
R38578 vdd.n10446 vdd.n10443 61.358
R38579 vdd.n10446 vdd.n10445 61.358
R38580 vdd.n10613 vdd.n10610 61.358
R38581 vdd.n10613 vdd.n10612 61.358
R38582 vdd.n10762 vdd.n10759 61.358
R38583 vdd.n10762 vdd.n10761 61.358
R38584 vdd.n10754 vdd.n10751 61.358
R38585 vdd.n10754 vdd.n10753 61.358
R38586 vdd.n10746 vdd.n10743 61.358
R38587 vdd.n10746 vdd.n10745 61.358
R38588 vdd.n10738 vdd.n10735 61.358
R38589 vdd.n10738 vdd.n10737 61.358
R38590 vdd.n10730 vdd.n10727 61.358
R38591 vdd.n10730 vdd.n10729 61.358
R38592 vdd.n10722 vdd.n10719 61.358
R38593 vdd.n10722 vdd.n10721 61.358
R38594 vdd.n10714 vdd.n10711 61.358
R38595 vdd.n10714 vdd.n10713 61.358
R38596 vdd.n10706 vdd.n10703 61.358
R38597 vdd.n10706 vdd.n10705 61.358
R38598 vdd.n10698 vdd.n10695 61.358
R38599 vdd.n10698 vdd.n10697 61.358
R38600 vdd.n10682 vdd.n10679 61.358
R38601 vdd.n10682 vdd.n10681 61.358
R38602 vdd.n10674 vdd.n10671 61.358
R38603 vdd.n10674 vdd.n10673 61.358
R38604 vdd.n10666 vdd.n10663 61.358
R38605 vdd.n10666 vdd.n10665 61.358
R38606 vdd.n10658 vdd.n10655 61.358
R38607 vdd.n10658 vdd.n10657 61.358
R38608 vdd.n10650 vdd.n10647 61.358
R38609 vdd.n10650 vdd.n10649 61.358
R38610 vdd.n10642 vdd.n10639 61.358
R38611 vdd.n10642 vdd.n10641 61.358
R38612 vdd.n10634 vdd.n10631 61.358
R38613 vdd.n10634 vdd.n10633 61.358
R38614 vdd.n10626 vdd.n10623 61.358
R38615 vdd.n10626 vdd.n10625 61.358
R38616 vdd.n10793 vdd.n10790 61.358
R38617 vdd.n10793 vdd.n10792 61.358
R38618 vdd.n10942 vdd.n10939 61.358
R38619 vdd.n10942 vdd.n10941 61.358
R38620 vdd.n10934 vdd.n10931 61.358
R38621 vdd.n10934 vdd.n10933 61.358
R38622 vdd.n10926 vdd.n10923 61.358
R38623 vdd.n10926 vdd.n10925 61.358
R38624 vdd.n10918 vdd.n10915 61.358
R38625 vdd.n10918 vdd.n10917 61.358
R38626 vdd.n10910 vdd.n10907 61.358
R38627 vdd.n10910 vdd.n10909 61.358
R38628 vdd.n10902 vdd.n10899 61.358
R38629 vdd.n10902 vdd.n10901 61.358
R38630 vdd.n10894 vdd.n10891 61.358
R38631 vdd.n10894 vdd.n10893 61.358
R38632 vdd.n10886 vdd.n10883 61.358
R38633 vdd.n10886 vdd.n10885 61.358
R38634 vdd.n10878 vdd.n10875 61.358
R38635 vdd.n10878 vdd.n10877 61.358
R38636 vdd.n10862 vdd.n10859 61.358
R38637 vdd.n10862 vdd.n10861 61.358
R38638 vdd.n10854 vdd.n10851 61.358
R38639 vdd.n10854 vdd.n10853 61.358
R38640 vdd.n10846 vdd.n10843 61.358
R38641 vdd.n10846 vdd.n10845 61.358
R38642 vdd.n10838 vdd.n10835 61.358
R38643 vdd.n10838 vdd.n10837 61.358
R38644 vdd.n10830 vdd.n10827 61.358
R38645 vdd.n10830 vdd.n10829 61.358
R38646 vdd.n10822 vdd.n10819 61.358
R38647 vdd.n10822 vdd.n10821 61.358
R38648 vdd.n10814 vdd.n10811 61.358
R38649 vdd.n10814 vdd.n10813 61.358
R38650 vdd.n10806 vdd.n10803 61.358
R38651 vdd.n10806 vdd.n10805 61.358
R38652 vdd.n10973 vdd.n10970 61.358
R38653 vdd.n10973 vdd.n10972 61.358
R38654 vdd.n11122 vdd.n11119 61.358
R38655 vdd.n11122 vdd.n11121 61.358
R38656 vdd.n11114 vdd.n11111 61.358
R38657 vdd.n11114 vdd.n11113 61.358
R38658 vdd.n11106 vdd.n11103 61.358
R38659 vdd.n11106 vdd.n11105 61.358
R38660 vdd.n11098 vdd.n11095 61.358
R38661 vdd.n11098 vdd.n11097 61.358
R38662 vdd.n11090 vdd.n11087 61.358
R38663 vdd.n11090 vdd.n11089 61.358
R38664 vdd.n11082 vdd.n11079 61.358
R38665 vdd.n11082 vdd.n11081 61.358
R38666 vdd.n11074 vdd.n11071 61.358
R38667 vdd.n11074 vdd.n11073 61.358
R38668 vdd.n11066 vdd.n11063 61.358
R38669 vdd.n11066 vdd.n11065 61.358
R38670 vdd.n11058 vdd.n11055 61.358
R38671 vdd.n11058 vdd.n11057 61.358
R38672 vdd.n11042 vdd.n11039 61.358
R38673 vdd.n11042 vdd.n11041 61.358
R38674 vdd.n11034 vdd.n11031 61.358
R38675 vdd.n11034 vdd.n11033 61.358
R38676 vdd.n11026 vdd.n11023 61.358
R38677 vdd.n11026 vdd.n11025 61.358
R38678 vdd.n11018 vdd.n11015 61.358
R38679 vdd.n11018 vdd.n11017 61.358
R38680 vdd.n11010 vdd.n11007 61.358
R38681 vdd.n11010 vdd.n11009 61.358
R38682 vdd.n11002 vdd.n10999 61.358
R38683 vdd.n11002 vdd.n11001 61.358
R38684 vdd.n10994 vdd.n10991 61.358
R38685 vdd.n10994 vdd.n10993 61.358
R38686 vdd.n10986 vdd.n10983 61.358
R38687 vdd.n10986 vdd.n10985 61.358
R38688 vdd.n11153 vdd.n11150 61.358
R38689 vdd.n11153 vdd.n11152 61.358
R38690 vdd.n11302 vdd.n11299 61.358
R38691 vdd.n11302 vdd.n11301 61.358
R38692 vdd.n11294 vdd.n11291 61.358
R38693 vdd.n11294 vdd.n11293 61.358
R38694 vdd.n11286 vdd.n11283 61.358
R38695 vdd.n11286 vdd.n11285 61.358
R38696 vdd.n11278 vdd.n11275 61.358
R38697 vdd.n11278 vdd.n11277 61.358
R38698 vdd.n11270 vdd.n11267 61.358
R38699 vdd.n11270 vdd.n11269 61.358
R38700 vdd.n11262 vdd.n11259 61.358
R38701 vdd.n11262 vdd.n11261 61.358
R38702 vdd.n11254 vdd.n11251 61.358
R38703 vdd.n11254 vdd.n11253 61.358
R38704 vdd.n11246 vdd.n11243 61.358
R38705 vdd.n11246 vdd.n11245 61.358
R38706 vdd.n11238 vdd.n11235 61.358
R38707 vdd.n11238 vdd.n11237 61.358
R38708 vdd.n11222 vdd.n11219 61.358
R38709 vdd.n11222 vdd.n11221 61.358
R38710 vdd.n11214 vdd.n11211 61.358
R38711 vdd.n11214 vdd.n11213 61.358
R38712 vdd.n11206 vdd.n11203 61.358
R38713 vdd.n11206 vdd.n11205 61.358
R38714 vdd.n11198 vdd.n11195 61.358
R38715 vdd.n11198 vdd.n11197 61.358
R38716 vdd.n11190 vdd.n11187 61.358
R38717 vdd.n11190 vdd.n11189 61.358
R38718 vdd.n11182 vdd.n11179 61.358
R38719 vdd.n11182 vdd.n11181 61.358
R38720 vdd.n11174 vdd.n11171 61.358
R38721 vdd.n11174 vdd.n11173 61.358
R38722 vdd.n11166 vdd.n11163 61.358
R38723 vdd.n11166 vdd.n11165 61.358
R38724 vdd.n11333 vdd.n11330 61.358
R38725 vdd.n11333 vdd.n11332 61.358
R38726 vdd.n13351 vdd.n13350 61
R38727 vdd.n13351 vdd.n13349 61
R38728 vdd.n13171 vdd.n13170 61
R38729 vdd.n13171 vdd.n13169 61
R38730 vdd.n12991 vdd.n12990 61
R38731 vdd.n12991 vdd.n12989 61
R38732 vdd.n12811 vdd.n12810 61
R38733 vdd.n12811 vdd.n12809 61
R38734 vdd.n12631 vdd.n12630 61
R38735 vdd.n12631 vdd.n12629 61
R38736 vdd.n12451 vdd.n12450 61
R38737 vdd.n12451 vdd.n12449 61
R38738 vdd.n12271 vdd.n12270 61
R38739 vdd.n12271 vdd.n12269 61
R38740 vdd.n12091 vdd.n12090 61
R38741 vdd.n12091 vdd.n12089 61
R38742 vdd.n11911 vdd.n11910 61
R38743 vdd.n11911 vdd.n11909 61
R38744 vdd.n11731 vdd.n11730 61
R38745 vdd.n11731 vdd.n11729 61
R38746 vdd.n11551 vdd.n11550 61
R38747 vdd.n11551 vdd.n11549 61
R38748 vdd.n72 vdd.n71 61
R38749 vdd.n72 vdd.n70 61
R38750 vdd.n252 vdd.n251 61
R38751 vdd.n252 vdd.n250 61
R38752 vdd.n432 vdd.n431 61
R38753 vdd.n432 vdd.n430 61
R38754 vdd.n612 vdd.n611 61
R38755 vdd.n612 vdd.n610 61
R38756 vdd.n792 vdd.n791 61
R38757 vdd.n792 vdd.n790 61
R38758 vdd.n972 vdd.n971 61
R38759 vdd.n972 vdd.n970 61
R38760 vdd.n1152 vdd.n1151 61
R38761 vdd.n1152 vdd.n1150 61
R38762 vdd.n1332 vdd.n1331 61
R38763 vdd.n1332 vdd.n1330 61
R38764 vdd.n1512 vdd.n1511 61
R38765 vdd.n1512 vdd.n1510 61
R38766 vdd.n1692 vdd.n1691 61
R38767 vdd.n1692 vdd.n1690 61
R38768 vdd.n1872 vdd.n1871 61
R38769 vdd.n1872 vdd.n1870 61
R38770 vdd.n2052 vdd.n2051 61
R38771 vdd.n2052 vdd.n2050 61
R38772 vdd.n2232 vdd.n2231 61
R38773 vdd.n2232 vdd.n2230 61
R38774 vdd.n2412 vdd.n2411 61
R38775 vdd.n2412 vdd.n2410 61
R38776 vdd.n2592 vdd.n2591 61
R38777 vdd.n2592 vdd.n2590 61
R38778 vdd.n2772 vdd.n2771 61
R38779 vdd.n2772 vdd.n2770 61
R38780 vdd.n2952 vdd.n2951 61
R38781 vdd.n2952 vdd.n2950 61
R38782 vdd.n3132 vdd.n3131 61
R38783 vdd.n3132 vdd.n3130 61
R38784 vdd.n3312 vdd.n3311 61
R38785 vdd.n3312 vdd.n3310 61
R38786 vdd.n3492 vdd.n3491 61
R38787 vdd.n3492 vdd.n3490 61
R38788 vdd.n3672 vdd.n3671 61
R38789 vdd.n3672 vdd.n3670 61
R38790 vdd.n3852 vdd.n3851 61
R38791 vdd.n3852 vdd.n3850 61
R38792 vdd.n4032 vdd.n4031 61
R38793 vdd.n4032 vdd.n4030 61
R38794 vdd.n4212 vdd.n4211 61
R38795 vdd.n4212 vdd.n4210 61
R38796 vdd.n4392 vdd.n4391 61
R38797 vdd.n4392 vdd.n4390 61
R38798 vdd.n4572 vdd.n4571 61
R38799 vdd.n4572 vdd.n4570 61
R38800 vdd.n4752 vdd.n4751 61
R38801 vdd.n4752 vdd.n4750 61
R38802 vdd.n4932 vdd.n4931 61
R38803 vdd.n4932 vdd.n4930 61
R38804 vdd.n5112 vdd.n5111 61
R38805 vdd.n5112 vdd.n5110 61
R38806 vdd.n5292 vdd.n5291 61
R38807 vdd.n5292 vdd.n5290 61
R38808 vdd.n5472 vdd.n5471 61
R38809 vdd.n5472 vdd.n5470 61
R38810 vdd.n5652 vdd.n5651 61
R38811 vdd.n5652 vdd.n5650 61
R38812 vdd.n5832 vdd.n5831 61
R38813 vdd.n5832 vdd.n5830 61
R38814 vdd.n6012 vdd.n6011 61
R38815 vdd.n6012 vdd.n6010 61
R38816 vdd.n6192 vdd.n6191 61
R38817 vdd.n6192 vdd.n6190 61
R38818 vdd.n6372 vdd.n6371 61
R38819 vdd.n6372 vdd.n6370 61
R38820 vdd.n6552 vdd.n6551 61
R38821 vdd.n6552 vdd.n6550 61
R38822 vdd.n6732 vdd.n6731 61
R38823 vdd.n6732 vdd.n6730 61
R38824 vdd.n6912 vdd.n6911 61
R38825 vdd.n6912 vdd.n6910 61
R38826 vdd.n7092 vdd.n7091 61
R38827 vdd.n7092 vdd.n7090 61
R38828 vdd.n7272 vdd.n7271 61
R38829 vdd.n7272 vdd.n7270 61
R38830 vdd.n7452 vdd.n7451 61
R38831 vdd.n7452 vdd.n7450 61
R38832 vdd.n7632 vdd.n7631 61
R38833 vdd.n7632 vdd.n7630 61
R38834 vdd.n7812 vdd.n7811 61
R38835 vdd.n7812 vdd.n7810 61
R38836 vdd.n7992 vdd.n7991 61
R38837 vdd.n7992 vdd.n7990 61
R38838 vdd.n8172 vdd.n8171 61
R38839 vdd.n8172 vdd.n8170 61
R38840 vdd.n8352 vdd.n8351 61
R38841 vdd.n8352 vdd.n8350 61
R38842 vdd.n8532 vdd.n8531 61
R38843 vdd.n8532 vdd.n8530 61
R38844 vdd.n8712 vdd.n8711 61
R38845 vdd.n8712 vdd.n8710 61
R38846 vdd.n8892 vdd.n8891 61
R38847 vdd.n8892 vdd.n8890 61
R38848 vdd.n9072 vdd.n9071 61
R38849 vdd.n9072 vdd.n9070 61
R38850 vdd.n9252 vdd.n9251 61
R38851 vdd.n9252 vdd.n9250 61
R38852 vdd.n9432 vdd.n9431 61
R38853 vdd.n9432 vdd.n9430 61
R38854 vdd.n9612 vdd.n9611 61
R38855 vdd.n9612 vdd.n9610 61
R38856 vdd.n9792 vdd.n9791 61
R38857 vdd.n9792 vdd.n9790 61
R38858 vdd.n9972 vdd.n9971 61
R38859 vdd.n9972 vdd.n9970 61
R38860 vdd.n10152 vdd.n10151 61
R38861 vdd.n10152 vdd.n10150 61
R38862 vdd.n10332 vdd.n10331 61
R38863 vdd.n10332 vdd.n10330 61
R38864 vdd.n10512 vdd.n10511 61
R38865 vdd.n10512 vdd.n10510 61
R38866 vdd.n10692 vdd.n10691 61
R38867 vdd.n10692 vdd.n10690 61
R38868 vdd.n10872 vdd.n10871 61
R38869 vdd.n10872 vdd.n10870 61
R38870 vdd.n11052 vdd.n11051 61
R38871 vdd.n11052 vdd.n11050 61
R38872 vdd.n11232 vdd.n11231 61
R38873 vdd.n11232 vdd.n11230 61
R38874 vdd.n11360 vdd.n11357 53.134
R38875 vdd.n11363 vdd.n11356 53.134
R38876 vdd.n11366 vdd.n11355 53.134
R38877 vdd.n11369 vdd.n11354 53.134
R38878 vdd.n11372 vdd.n11353 53.134
R38879 vdd.n11375 vdd.n11352 53.134
R38880 vdd.n11378 vdd.n11351 53.134
R38881 vdd.n11381 vdd.n11350 53.134
R38882 vdd.n11384 vdd.n11349 53.134
R38883 vdd.n11388 vdd.n11347 53.134
R38884 vdd.n11391 vdd.n11346 53.134
R38885 vdd.n11394 vdd.n11345 53.134
R38886 vdd.n11397 vdd.n11344 53.134
R38887 vdd.n11400 vdd.n11343 53.134
R38888 vdd.n11403 vdd.n11342 53.134
R38889 vdd.n11406 vdd.n11341 53.134
R38890 vdd.n11409 vdd.n11340 53.134
R38891 vdd.n11413 vdd.n11412 53.134
R38892 vdd.n13482 vdd.n13475 51.368
R38893 vdd.n13485 vdd.n13474 51.368
R38894 vdd.n13488 vdd.n13473 51.368
R38895 vdd.n13491 vdd.n13472 51.368
R38896 vdd.n13494 vdd.n13471 51.368
R38897 vdd.n13497 vdd.n13470 51.368
R38898 vdd.n13500 vdd.n13469 51.368
R38899 vdd.n13503 vdd.n13468 51.368
R38900 vdd.n13507 vdd.n13466 51.368
R38901 vdd.n13510 vdd.n13465 51.368
R38902 vdd.n13513 vdd.n13464 51.368
R38903 vdd.n13516 vdd.n13463 51.368
R38904 vdd.n13519 vdd.n13462 51.368
R38905 vdd.n13522 vdd.n13461 51.368
R38906 vdd.n13525 vdd.n13460 51.368
R38907 vdd.n13528 vdd.n13459 51.368
R38908 vdd.n13532 vdd.n13531 51.368
R38909 vdd.n13479 vdd.n13476 51.368
R38910 vdd.n13426 vdd.n13424 25.477
R38911 vdd.n13426 vdd.n13425 25.477
R38912 vdd.n13246 vdd.n13244 25.477
R38913 vdd.n13246 vdd.n13245 25.477
R38914 vdd.n13066 vdd.n13064 25.477
R38915 vdd.n13066 vdd.n13065 25.477
R38916 vdd.n12886 vdd.n12884 25.477
R38917 vdd.n12886 vdd.n12885 25.477
R38918 vdd.n12706 vdd.n12704 25.477
R38919 vdd.n12706 vdd.n12705 25.477
R38920 vdd.n12526 vdd.n12524 25.477
R38921 vdd.n12526 vdd.n12525 25.477
R38922 vdd.n12346 vdd.n12344 25.477
R38923 vdd.n12346 vdd.n12345 25.477
R38924 vdd.n12166 vdd.n12164 25.477
R38925 vdd.n12166 vdd.n12165 25.477
R38926 vdd.n11986 vdd.n11984 25.477
R38927 vdd.n11986 vdd.n11985 25.477
R38928 vdd.n11806 vdd.n11804 25.477
R38929 vdd.n11806 vdd.n11805 25.477
R38930 vdd.n11626 vdd.n11624 25.477
R38931 vdd.n11626 vdd.n11625 25.477
R38932 vdd.n147 vdd.n145 25.477
R38933 vdd.n147 vdd.n146 25.477
R38934 vdd.n327 vdd.n325 25.477
R38935 vdd.n327 vdd.n326 25.477
R38936 vdd.n507 vdd.n505 25.477
R38937 vdd.n507 vdd.n506 25.477
R38938 vdd.n687 vdd.n685 25.477
R38939 vdd.n687 vdd.n686 25.477
R38940 vdd.n867 vdd.n865 25.477
R38941 vdd.n867 vdd.n866 25.477
R38942 vdd.n1047 vdd.n1045 25.477
R38943 vdd.n1047 vdd.n1046 25.477
R38944 vdd.n1227 vdd.n1225 25.477
R38945 vdd.n1227 vdd.n1226 25.477
R38946 vdd.n1407 vdd.n1405 25.477
R38947 vdd.n1407 vdd.n1406 25.477
R38948 vdd.n1587 vdd.n1585 25.477
R38949 vdd.n1587 vdd.n1586 25.477
R38950 vdd.n1767 vdd.n1765 25.477
R38951 vdd.n1767 vdd.n1766 25.477
R38952 vdd.n1947 vdd.n1945 25.477
R38953 vdd.n1947 vdd.n1946 25.477
R38954 vdd.n2127 vdd.n2125 25.477
R38955 vdd.n2127 vdd.n2126 25.477
R38956 vdd.n2307 vdd.n2305 25.477
R38957 vdd.n2307 vdd.n2306 25.477
R38958 vdd.n2487 vdd.n2485 25.477
R38959 vdd.n2487 vdd.n2486 25.477
R38960 vdd.n2667 vdd.n2665 25.477
R38961 vdd.n2667 vdd.n2666 25.477
R38962 vdd.n2847 vdd.n2845 25.477
R38963 vdd.n2847 vdd.n2846 25.477
R38964 vdd.n3027 vdd.n3025 25.477
R38965 vdd.n3027 vdd.n3026 25.477
R38966 vdd.n3207 vdd.n3205 25.477
R38967 vdd.n3207 vdd.n3206 25.477
R38968 vdd.n3387 vdd.n3385 25.477
R38969 vdd.n3387 vdd.n3386 25.477
R38970 vdd.n3567 vdd.n3565 25.477
R38971 vdd.n3567 vdd.n3566 25.477
R38972 vdd.n3747 vdd.n3745 25.477
R38973 vdd.n3747 vdd.n3746 25.477
R38974 vdd.n3927 vdd.n3925 25.477
R38975 vdd.n3927 vdd.n3926 25.477
R38976 vdd.n4107 vdd.n4105 25.477
R38977 vdd.n4107 vdd.n4106 25.477
R38978 vdd.n4287 vdd.n4285 25.477
R38979 vdd.n4287 vdd.n4286 25.477
R38980 vdd.n4467 vdd.n4465 25.477
R38981 vdd.n4467 vdd.n4466 25.477
R38982 vdd.n4647 vdd.n4645 25.477
R38983 vdd.n4647 vdd.n4646 25.477
R38984 vdd.n4827 vdd.n4825 25.477
R38985 vdd.n4827 vdd.n4826 25.477
R38986 vdd.n5007 vdd.n5005 25.477
R38987 vdd.n5007 vdd.n5006 25.477
R38988 vdd.n5187 vdd.n5185 25.477
R38989 vdd.n5187 vdd.n5186 25.477
R38990 vdd.n5367 vdd.n5365 25.477
R38991 vdd.n5367 vdd.n5366 25.477
R38992 vdd.n5547 vdd.n5545 25.477
R38993 vdd.n5547 vdd.n5546 25.477
R38994 vdd.n5727 vdd.n5725 25.477
R38995 vdd.n5727 vdd.n5726 25.477
R38996 vdd.n5907 vdd.n5905 25.477
R38997 vdd.n5907 vdd.n5906 25.477
R38998 vdd.n6087 vdd.n6085 25.477
R38999 vdd.n6087 vdd.n6086 25.477
R39000 vdd.n6267 vdd.n6265 25.477
R39001 vdd.n6267 vdd.n6266 25.477
R39002 vdd.n6447 vdd.n6445 25.477
R39003 vdd.n6447 vdd.n6446 25.477
R39004 vdd.n6627 vdd.n6625 25.477
R39005 vdd.n6627 vdd.n6626 25.477
R39006 vdd.n6807 vdd.n6805 25.477
R39007 vdd.n6807 vdd.n6806 25.477
R39008 vdd.n6987 vdd.n6985 25.477
R39009 vdd.n6987 vdd.n6986 25.477
R39010 vdd.n7167 vdd.n7165 25.477
R39011 vdd.n7167 vdd.n7166 25.477
R39012 vdd.n7347 vdd.n7345 25.477
R39013 vdd.n7347 vdd.n7346 25.477
R39014 vdd.n7527 vdd.n7525 25.477
R39015 vdd.n7527 vdd.n7526 25.477
R39016 vdd.n7707 vdd.n7705 25.477
R39017 vdd.n7707 vdd.n7706 25.477
R39018 vdd.n7887 vdd.n7885 25.477
R39019 vdd.n7887 vdd.n7886 25.477
R39020 vdd.n8067 vdd.n8065 25.477
R39021 vdd.n8067 vdd.n8066 25.477
R39022 vdd.n8247 vdd.n8245 25.477
R39023 vdd.n8247 vdd.n8246 25.477
R39024 vdd.n8427 vdd.n8425 25.477
R39025 vdd.n8427 vdd.n8426 25.477
R39026 vdd.n8607 vdd.n8605 25.477
R39027 vdd.n8607 vdd.n8606 25.477
R39028 vdd.n8787 vdd.n8785 25.477
R39029 vdd.n8787 vdd.n8786 25.477
R39030 vdd.n8967 vdd.n8965 25.477
R39031 vdd.n8967 vdd.n8966 25.477
R39032 vdd.n9147 vdd.n9145 25.477
R39033 vdd.n9147 vdd.n9146 25.477
R39034 vdd.n9327 vdd.n9325 25.477
R39035 vdd.n9327 vdd.n9326 25.477
R39036 vdd.n9507 vdd.n9505 25.477
R39037 vdd.n9507 vdd.n9506 25.477
R39038 vdd.n9687 vdd.n9685 25.477
R39039 vdd.n9687 vdd.n9686 25.477
R39040 vdd.n9867 vdd.n9865 25.477
R39041 vdd.n9867 vdd.n9866 25.477
R39042 vdd.n10047 vdd.n10045 25.477
R39043 vdd.n10047 vdd.n10046 25.477
R39044 vdd.n10227 vdd.n10225 25.477
R39045 vdd.n10227 vdd.n10226 25.477
R39046 vdd.n10407 vdd.n10405 25.477
R39047 vdd.n10407 vdd.n10406 25.477
R39048 vdd.n10587 vdd.n10585 25.477
R39049 vdd.n10587 vdd.n10586 25.477
R39050 vdd.n10767 vdd.n10765 25.477
R39051 vdd.n10767 vdd.n10766 25.477
R39052 vdd.n10947 vdd.n10945 25.477
R39053 vdd.n10947 vdd.n10946 25.477
R39054 vdd.n11127 vdd.n11125 25.477
R39055 vdd.n11127 vdd.n11126 25.477
R39056 vdd.n11307 vdd.n11305 25.477
R39057 vdd.n11307 vdd.n11306 25.477
R39058 vdd.n13457 vdd.n13455 24.759
R39059 vdd.n13457 vdd.n13456 24.759
R39060 vdd.n13277 vdd.n13275 24.759
R39061 vdd.n13277 vdd.n13276 24.759
R39062 vdd.n13097 vdd.n13095 24.759
R39063 vdd.n13097 vdd.n13096 24.759
R39064 vdd.n12917 vdd.n12915 24.759
R39065 vdd.n12917 vdd.n12916 24.759
R39066 vdd.n12737 vdd.n12735 24.759
R39067 vdd.n12737 vdd.n12736 24.759
R39068 vdd.n12557 vdd.n12555 24.759
R39069 vdd.n12557 vdd.n12556 24.759
R39070 vdd.n12377 vdd.n12375 24.759
R39071 vdd.n12377 vdd.n12376 24.759
R39072 vdd.n12197 vdd.n12195 24.759
R39073 vdd.n12197 vdd.n12196 24.759
R39074 vdd.n12017 vdd.n12015 24.759
R39075 vdd.n12017 vdd.n12016 24.759
R39076 vdd.n11837 vdd.n11835 24.759
R39077 vdd.n11837 vdd.n11836 24.759
R39078 vdd.n11657 vdd.n11655 24.759
R39079 vdd.n11657 vdd.n11656 24.759
R39080 vdd.n178 vdd.n176 24.759
R39081 vdd.n178 vdd.n177 24.759
R39082 vdd.n358 vdd.n356 24.759
R39083 vdd.n358 vdd.n357 24.759
R39084 vdd.n538 vdd.n536 24.759
R39085 vdd.n538 vdd.n537 24.759
R39086 vdd.n718 vdd.n716 24.759
R39087 vdd.n718 vdd.n717 24.759
R39088 vdd.n898 vdd.n896 24.759
R39089 vdd.n898 vdd.n897 24.759
R39090 vdd.n1078 vdd.n1076 24.759
R39091 vdd.n1078 vdd.n1077 24.759
R39092 vdd.n1258 vdd.n1256 24.759
R39093 vdd.n1258 vdd.n1257 24.759
R39094 vdd.n1438 vdd.n1436 24.759
R39095 vdd.n1438 vdd.n1437 24.759
R39096 vdd.n1618 vdd.n1616 24.759
R39097 vdd.n1618 vdd.n1617 24.759
R39098 vdd.n1798 vdd.n1796 24.759
R39099 vdd.n1798 vdd.n1797 24.759
R39100 vdd.n1978 vdd.n1976 24.759
R39101 vdd.n1978 vdd.n1977 24.759
R39102 vdd.n2158 vdd.n2156 24.759
R39103 vdd.n2158 vdd.n2157 24.759
R39104 vdd.n2338 vdd.n2336 24.759
R39105 vdd.n2338 vdd.n2337 24.759
R39106 vdd.n2518 vdd.n2516 24.759
R39107 vdd.n2518 vdd.n2517 24.759
R39108 vdd.n2698 vdd.n2696 24.759
R39109 vdd.n2698 vdd.n2697 24.759
R39110 vdd.n2878 vdd.n2876 24.759
R39111 vdd.n2878 vdd.n2877 24.759
R39112 vdd.n3058 vdd.n3056 24.759
R39113 vdd.n3058 vdd.n3057 24.759
R39114 vdd.n3238 vdd.n3236 24.759
R39115 vdd.n3238 vdd.n3237 24.759
R39116 vdd.n3418 vdd.n3416 24.759
R39117 vdd.n3418 vdd.n3417 24.759
R39118 vdd.n3598 vdd.n3596 24.759
R39119 vdd.n3598 vdd.n3597 24.759
R39120 vdd.n3778 vdd.n3776 24.759
R39121 vdd.n3778 vdd.n3777 24.759
R39122 vdd.n3958 vdd.n3956 24.759
R39123 vdd.n3958 vdd.n3957 24.759
R39124 vdd.n4138 vdd.n4136 24.759
R39125 vdd.n4138 vdd.n4137 24.759
R39126 vdd.n4318 vdd.n4316 24.759
R39127 vdd.n4318 vdd.n4317 24.759
R39128 vdd.n4498 vdd.n4496 24.759
R39129 vdd.n4498 vdd.n4497 24.759
R39130 vdd.n4678 vdd.n4676 24.759
R39131 vdd.n4678 vdd.n4677 24.759
R39132 vdd.n4858 vdd.n4856 24.759
R39133 vdd.n4858 vdd.n4857 24.759
R39134 vdd.n5038 vdd.n5036 24.759
R39135 vdd.n5038 vdd.n5037 24.759
R39136 vdd.n5218 vdd.n5216 24.759
R39137 vdd.n5218 vdd.n5217 24.759
R39138 vdd.n5398 vdd.n5396 24.759
R39139 vdd.n5398 vdd.n5397 24.759
R39140 vdd.n5578 vdd.n5576 24.759
R39141 vdd.n5578 vdd.n5577 24.759
R39142 vdd.n5758 vdd.n5756 24.759
R39143 vdd.n5758 vdd.n5757 24.759
R39144 vdd.n5938 vdd.n5936 24.759
R39145 vdd.n5938 vdd.n5937 24.759
R39146 vdd.n6118 vdd.n6116 24.759
R39147 vdd.n6118 vdd.n6117 24.759
R39148 vdd.n6298 vdd.n6296 24.759
R39149 vdd.n6298 vdd.n6297 24.759
R39150 vdd.n6478 vdd.n6476 24.759
R39151 vdd.n6478 vdd.n6477 24.759
R39152 vdd.n6658 vdd.n6656 24.759
R39153 vdd.n6658 vdd.n6657 24.759
R39154 vdd.n6838 vdd.n6836 24.759
R39155 vdd.n6838 vdd.n6837 24.759
R39156 vdd.n7018 vdd.n7016 24.759
R39157 vdd.n7018 vdd.n7017 24.759
R39158 vdd.n7198 vdd.n7196 24.759
R39159 vdd.n7198 vdd.n7197 24.759
R39160 vdd.n7378 vdd.n7376 24.759
R39161 vdd.n7378 vdd.n7377 24.759
R39162 vdd.n7558 vdd.n7556 24.759
R39163 vdd.n7558 vdd.n7557 24.759
R39164 vdd.n7738 vdd.n7736 24.759
R39165 vdd.n7738 vdd.n7737 24.759
R39166 vdd.n7918 vdd.n7916 24.759
R39167 vdd.n7918 vdd.n7917 24.759
R39168 vdd.n8098 vdd.n8096 24.759
R39169 vdd.n8098 vdd.n8097 24.759
R39170 vdd.n8278 vdd.n8276 24.759
R39171 vdd.n8278 vdd.n8277 24.759
R39172 vdd.n8458 vdd.n8456 24.759
R39173 vdd.n8458 vdd.n8457 24.759
R39174 vdd.n8638 vdd.n8636 24.759
R39175 vdd.n8638 vdd.n8637 24.759
R39176 vdd.n8818 vdd.n8816 24.759
R39177 vdd.n8818 vdd.n8817 24.759
R39178 vdd.n8998 vdd.n8996 24.759
R39179 vdd.n8998 vdd.n8997 24.759
R39180 vdd.n9178 vdd.n9176 24.759
R39181 vdd.n9178 vdd.n9177 24.759
R39182 vdd.n9358 vdd.n9356 24.759
R39183 vdd.n9358 vdd.n9357 24.759
R39184 vdd.n9538 vdd.n9536 24.759
R39185 vdd.n9538 vdd.n9537 24.759
R39186 vdd.n9718 vdd.n9716 24.759
R39187 vdd.n9718 vdd.n9717 24.759
R39188 vdd.n9898 vdd.n9896 24.759
R39189 vdd.n9898 vdd.n9897 24.759
R39190 vdd.n10078 vdd.n10076 24.759
R39191 vdd.n10078 vdd.n10077 24.759
R39192 vdd.n10258 vdd.n10256 24.759
R39193 vdd.n10258 vdd.n10257 24.759
R39194 vdd.n10438 vdd.n10436 24.759
R39195 vdd.n10438 vdd.n10437 24.759
R39196 vdd.n10618 vdd.n10616 24.759
R39197 vdd.n10618 vdd.n10617 24.759
R39198 vdd.n10798 vdd.n10796 24.759
R39199 vdd.n10798 vdd.n10797 24.759
R39200 vdd.n10978 vdd.n10976 24.759
R39201 vdd.n10978 vdd.n10977 24.759
R39202 vdd.n11158 vdd.n11156 24.759
R39203 vdd.n11158 vdd.n11157 24.759
R39204 vdd.n11338 vdd.n11336 24.759
R39205 vdd.n11338 vdd.n11337 24.759
R39206 vdd.n13429 vdd.n13428 23.783
R39207 vdd.n13429 vdd.n13426 23.783
R39208 vdd.n13430 vdd.n13415 23.783
R39209 vdd.n13430 vdd.n13421 23.783
R39210 vdd.n13431 vdd.n13407 23.783
R39211 vdd.n13431 vdd.n13413 23.783
R39212 vdd.n13432 vdd.n13399 23.783
R39213 vdd.n13432 vdd.n13405 23.783
R39214 vdd.n13433 vdd.n13391 23.783
R39215 vdd.n13433 vdd.n13397 23.783
R39216 vdd.n13434 vdd.n13383 23.783
R39217 vdd.n13434 vdd.n13389 23.783
R39218 vdd.n13435 vdd.n13375 23.783
R39219 vdd.n13435 vdd.n13381 23.783
R39220 vdd.n13436 vdd.n13367 23.783
R39221 vdd.n13436 vdd.n13373 23.783
R39222 vdd.n13437 vdd.n13359 23.783
R39223 vdd.n13437 vdd.n13365 23.783
R39224 vdd.n13438 vdd.n13351 23.783
R39225 vdd.n13438 vdd.n13357 23.783
R39226 vdd.n13439 vdd.n13343 23.783
R39227 vdd.n13439 vdd.n13347 23.783
R39228 vdd.n13440 vdd.n13335 23.783
R39229 vdd.n13440 vdd.n13341 23.783
R39230 vdd.n13441 vdd.n13327 23.783
R39231 vdd.n13441 vdd.n13333 23.783
R39232 vdd.n13442 vdd.n13319 23.783
R39233 vdd.n13442 vdd.n13325 23.783
R39234 vdd.n13443 vdd.n13311 23.783
R39235 vdd.n13443 vdd.n13317 23.783
R39236 vdd.n13444 vdd.n13303 23.783
R39237 vdd.n13444 vdd.n13309 23.783
R39238 vdd.n13445 vdd.n13295 23.783
R39239 vdd.n13445 vdd.n13301 23.783
R39240 vdd.n13446 vdd.n13287 23.783
R39241 vdd.n13446 vdd.n13293 23.783
R39242 vdd.n13447 vdd.n13279 23.783
R39243 vdd.n13447 vdd.n13285 23.783
R39244 vdd.n13458 vdd.n13457 23.783
R39245 vdd.n13458 vdd.n13452 23.783
R39246 vdd.n13249 vdd.n13248 23.783
R39247 vdd.n13249 vdd.n13246 23.783
R39248 vdd.n13250 vdd.n13235 23.783
R39249 vdd.n13250 vdd.n13241 23.783
R39250 vdd.n13251 vdd.n13227 23.783
R39251 vdd.n13251 vdd.n13233 23.783
R39252 vdd.n13252 vdd.n13219 23.783
R39253 vdd.n13252 vdd.n13225 23.783
R39254 vdd.n13253 vdd.n13211 23.783
R39255 vdd.n13253 vdd.n13217 23.783
R39256 vdd.n13254 vdd.n13203 23.783
R39257 vdd.n13254 vdd.n13209 23.783
R39258 vdd.n13255 vdd.n13195 23.783
R39259 vdd.n13255 vdd.n13201 23.783
R39260 vdd.n13256 vdd.n13187 23.783
R39261 vdd.n13256 vdd.n13193 23.783
R39262 vdd.n13257 vdd.n13179 23.783
R39263 vdd.n13257 vdd.n13185 23.783
R39264 vdd.n13258 vdd.n13171 23.783
R39265 vdd.n13258 vdd.n13177 23.783
R39266 vdd.n13259 vdd.n13163 23.783
R39267 vdd.n13259 vdd.n13167 23.783
R39268 vdd.n13260 vdd.n13155 23.783
R39269 vdd.n13260 vdd.n13161 23.783
R39270 vdd.n13261 vdd.n13147 23.783
R39271 vdd.n13261 vdd.n13153 23.783
R39272 vdd.n13262 vdd.n13139 23.783
R39273 vdd.n13262 vdd.n13145 23.783
R39274 vdd.n13263 vdd.n13131 23.783
R39275 vdd.n13263 vdd.n13137 23.783
R39276 vdd.n13264 vdd.n13123 23.783
R39277 vdd.n13264 vdd.n13129 23.783
R39278 vdd.n13265 vdd.n13115 23.783
R39279 vdd.n13265 vdd.n13121 23.783
R39280 vdd.n13266 vdd.n13107 23.783
R39281 vdd.n13266 vdd.n13113 23.783
R39282 vdd.n13267 vdd.n13099 23.783
R39283 vdd.n13267 vdd.n13105 23.783
R39284 vdd.n13278 vdd.n13277 23.783
R39285 vdd.n13278 vdd.n13272 23.783
R39286 vdd.n13069 vdd.n13068 23.783
R39287 vdd.n13069 vdd.n13066 23.783
R39288 vdd.n13070 vdd.n13055 23.783
R39289 vdd.n13070 vdd.n13061 23.783
R39290 vdd.n13071 vdd.n13047 23.783
R39291 vdd.n13071 vdd.n13053 23.783
R39292 vdd.n13072 vdd.n13039 23.783
R39293 vdd.n13072 vdd.n13045 23.783
R39294 vdd.n13073 vdd.n13031 23.783
R39295 vdd.n13073 vdd.n13037 23.783
R39296 vdd.n13074 vdd.n13023 23.783
R39297 vdd.n13074 vdd.n13029 23.783
R39298 vdd.n13075 vdd.n13015 23.783
R39299 vdd.n13075 vdd.n13021 23.783
R39300 vdd.n13076 vdd.n13007 23.783
R39301 vdd.n13076 vdd.n13013 23.783
R39302 vdd.n13077 vdd.n12999 23.783
R39303 vdd.n13077 vdd.n13005 23.783
R39304 vdd.n13078 vdd.n12991 23.783
R39305 vdd.n13078 vdd.n12997 23.783
R39306 vdd.n13079 vdd.n12983 23.783
R39307 vdd.n13079 vdd.n12987 23.783
R39308 vdd.n13080 vdd.n12975 23.783
R39309 vdd.n13080 vdd.n12981 23.783
R39310 vdd.n13081 vdd.n12967 23.783
R39311 vdd.n13081 vdd.n12973 23.783
R39312 vdd.n13082 vdd.n12959 23.783
R39313 vdd.n13082 vdd.n12965 23.783
R39314 vdd.n13083 vdd.n12951 23.783
R39315 vdd.n13083 vdd.n12957 23.783
R39316 vdd.n13084 vdd.n12943 23.783
R39317 vdd.n13084 vdd.n12949 23.783
R39318 vdd.n13085 vdd.n12935 23.783
R39319 vdd.n13085 vdd.n12941 23.783
R39320 vdd.n13086 vdd.n12927 23.783
R39321 vdd.n13086 vdd.n12933 23.783
R39322 vdd.n13087 vdd.n12919 23.783
R39323 vdd.n13087 vdd.n12925 23.783
R39324 vdd.n13098 vdd.n13097 23.783
R39325 vdd.n13098 vdd.n13092 23.783
R39326 vdd.n12889 vdd.n12888 23.783
R39327 vdd.n12889 vdd.n12886 23.783
R39328 vdd.n12890 vdd.n12875 23.783
R39329 vdd.n12890 vdd.n12881 23.783
R39330 vdd.n12891 vdd.n12867 23.783
R39331 vdd.n12891 vdd.n12873 23.783
R39332 vdd.n12892 vdd.n12859 23.783
R39333 vdd.n12892 vdd.n12865 23.783
R39334 vdd.n12893 vdd.n12851 23.783
R39335 vdd.n12893 vdd.n12857 23.783
R39336 vdd.n12894 vdd.n12843 23.783
R39337 vdd.n12894 vdd.n12849 23.783
R39338 vdd.n12895 vdd.n12835 23.783
R39339 vdd.n12895 vdd.n12841 23.783
R39340 vdd.n12896 vdd.n12827 23.783
R39341 vdd.n12896 vdd.n12833 23.783
R39342 vdd.n12897 vdd.n12819 23.783
R39343 vdd.n12897 vdd.n12825 23.783
R39344 vdd.n12898 vdd.n12811 23.783
R39345 vdd.n12898 vdd.n12817 23.783
R39346 vdd.n12899 vdd.n12803 23.783
R39347 vdd.n12899 vdd.n12807 23.783
R39348 vdd.n12900 vdd.n12795 23.783
R39349 vdd.n12900 vdd.n12801 23.783
R39350 vdd.n12901 vdd.n12787 23.783
R39351 vdd.n12901 vdd.n12793 23.783
R39352 vdd.n12902 vdd.n12779 23.783
R39353 vdd.n12902 vdd.n12785 23.783
R39354 vdd.n12903 vdd.n12771 23.783
R39355 vdd.n12903 vdd.n12777 23.783
R39356 vdd.n12904 vdd.n12763 23.783
R39357 vdd.n12904 vdd.n12769 23.783
R39358 vdd.n12905 vdd.n12755 23.783
R39359 vdd.n12905 vdd.n12761 23.783
R39360 vdd.n12906 vdd.n12747 23.783
R39361 vdd.n12906 vdd.n12753 23.783
R39362 vdd.n12907 vdd.n12739 23.783
R39363 vdd.n12907 vdd.n12745 23.783
R39364 vdd.n12918 vdd.n12917 23.783
R39365 vdd.n12918 vdd.n12912 23.783
R39366 vdd.n12709 vdd.n12708 23.783
R39367 vdd.n12709 vdd.n12706 23.783
R39368 vdd.n12710 vdd.n12695 23.783
R39369 vdd.n12710 vdd.n12701 23.783
R39370 vdd.n12711 vdd.n12687 23.783
R39371 vdd.n12711 vdd.n12693 23.783
R39372 vdd.n12712 vdd.n12679 23.783
R39373 vdd.n12712 vdd.n12685 23.783
R39374 vdd.n12713 vdd.n12671 23.783
R39375 vdd.n12713 vdd.n12677 23.783
R39376 vdd.n12714 vdd.n12663 23.783
R39377 vdd.n12714 vdd.n12669 23.783
R39378 vdd.n12715 vdd.n12655 23.783
R39379 vdd.n12715 vdd.n12661 23.783
R39380 vdd.n12716 vdd.n12647 23.783
R39381 vdd.n12716 vdd.n12653 23.783
R39382 vdd.n12717 vdd.n12639 23.783
R39383 vdd.n12717 vdd.n12645 23.783
R39384 vdd.n12718 vdd.n12631 23.783
R39385 vdd.n12718 vdd.n12637 23.783
R39386 vdd.n12719 vdd.n12623 23.783
R39387 vdd.n12719 vdd.n12627 23.783
R39388 vdd.n12720 vdd.n12615 23.783
R39389 vdd.n12720 vdd.n12621 23.783
R39390 vdd.n12721 vdd.n12607 23.783
R39391 vdd.n12721 vdd.n12613 23.783
R39392 vdd.n12722 vdd.n12599 23.783
R39393 vdd.n12722 vdd.n12605 23.783
R39394 vdd.n12723 vdd.n12591 23.783
R39395 vdd.n12723 vdd.n12597 23.783
R39396 vdd.n12724 vdd.n12583 23.783
R39397 vdd.n12724 vdd.n12589 23.783
R39398 vdd.n12725 vdd.n12575 23.783
R39399 vdd.n12725 vdd.n12581 23.783
R39400 vdd.n12726 vdd.n12567 23.783
R39401 vdd.n12726 vdd.n12573 23.783
R39402 vdd.n12727 vdd.n12559 23.783
R39403 vdd.n12727 vdd.n12565 23.783
R39404 vdd.n12738 vdd.n12737 23.783
R39405 vdd.n12738 vdd.n12732 23.783
R39406 vdd.n12529 vdd.n12528 23.783
R39407 vdd.n12529 vdd.n12526 23.783
R39408 vdd.n12530 vdd.n12515 23.783
R39409 vdd.n12530 vdd.n12521 23.783
R39410 vdd.n12531 vdd.n12507 23.783
R39411 vdd.n12531 vdd.n12513 23.783
R39412 vdd.n12532 vdd.n12499 23.783
R39413 vdd.n12532 vdd.n12505 23.783
R39414 vdd.n12533 vdd.n12491 23.783
R39415 vdd.n12533 vdd.n12497 23.783
R39416 vdd.n12534 vdd.n12483 23.783
R39417 vdd.n12534 vdd.n12489 23.783
R39418 vdd.n12535 vdd.n12475 23.783
R39419 vdd.n12535 vdd.n12481 23.783
R39420 vdd.n12536 vdd.n12467 23.783
R39421 vdd.n12536 vdd.n12473 23.783
R39422 vdd.n12537 vdd.n12459 23.783
R39423 vdd.n12537 vdd.n12465 23.783
R39424 vdd.n12538 vdd.n12451 23.783
R39425 vdd.n12538 vdd.n12457 23.783
R39426 vdd.n12539 vdd.n12443 23.783
R39427 vdd.n12539 vdd.n12447 23.783
R39428 vdd.n12540 vdd.n12435 23.783
R39429 vdd.n12540 vdd.n12441 23.783
R39430 vdd.n12541 vdd.n12427 23.783
R39431 vdd.n12541 vdd.n12433 23.783
R39432 vdd.n12542 vdd.n12419 23.783
R39433 vdd.n12542 vdd.n12425 23.783
R39434 vdd.n12543 vdd.n12411 23.783
R39435 vdd.n12543 vdd.n12417 23.783
R39436 vdd.n12544 vdd.n12403 23.783
R39437 vdd.n12544 vdd.n12409 23.783
R39438 vdd.n12545 vdd.n12395 23.783
R39439 vdd.n12545 vdd.n12401 23.783
R39440 vdd.n12546 vdd.n12387 23.783
R39441 vdd.n12546 vdd.n12393 23.783
R39442 vdd.n12547 vdd.n12379 23.783
R39443 vdd.n12547 vdd.n12385 23.783
R39444 vdd.n12558 vdd.n12557 23.783
R39445 vdd.n12558 vdd.n12552 23.783
R39446 vdd.n12349 vdd.n12348 23.783
R39447 vdd.n12349 vdd.n12346 23.783
R39448 vdd.n12350 vdd.n12335 23.783
R39449 vdd.n12350 vdd.n12341 23.783
R39450 vdd.n12351 vdd.n12327 23.783
R39451 vdd.n12351 vdd.n12333 23.783
R39452 vdd.n12352 vdd.n12319 23.783
R39453 vdd.n12352 vdd.n12325 23.783
R39454 vdd.n12353 vdd.n12311 23.783
R39455 vdd.n12353 vdd.n12317 23.783
R39456 vdd.n12354 vdd.n12303 23.783
R39457 vdd.n12354 vdd.n12309 23.783
R39458 vdd.n12355 vdd.n12295 23.783
R39459 vdd.n12355 vdd.n12301 23.783
R39460 vdd.n12356 vdd.n12287 23.783
R39461 vdd.n12356 vdd.n12293 23.783
R39462 vdd.n12357 vdd.n12279 23.783
R39463 vdd.n12357 vdd.n12285 23.783
R39464 vdd.n12358 vdd.n12271 23.783
R39465 vdd.n12358 vdd.n12277 23.783
R39466 vdd.n12359 vdd.n12263 23.783
R39467 vdd.n12359 vdd.n12267 23.783
R39468 vdd.n12360 vdd.n12255 23.783
R39469 vdd.n12360 vdd.n12261 23.783
R39470 vdd.n12361 vdd.n12247 23.783
R39471 vdd.n12361 vdd.n12253 23.783
R39472 vdd.n12362 vdd.n12239 23.783
R39473 vdd.n12362 vdd.n12245 23.783
R39474 vdd.n12363 vdd.n12231 23.783
R39475 vdd.n12363 vdd.n12237 23.783
R39476 vdd.n12364 vdd.n12223 23.783
R39477 vdd.n12364 vdd.n12229 23.783
R39478 vdd.n12365 vdd.n12215 23.783
R39479 vdd.n12365 vdd.n12221 23.783
R39480 vdd.n12366 vdd.n12207 23.783
R39481 vdd.n12366 vdd.n12213 23.783
R39482 vdd.n12367 vdd.n12199 23.783
R39483 vdd.n12367 vdd.n12205 23.783
R39484 vdd.n12378 vdd.n12377 23.783
R39485 vdd.n12378 vdd.n12372 23.783
R39486 vdd.n12169 vdd.n12168 23.783
R39487 vdd.n12169 vdd.n12166 23.783
R39488 vdd.n12170 vdd.n12155 23.783
R39489 vdd.n12170 vdd.n12161 23.783
R39490 vdd.n12171 vdd.n12147 23.783
R39491 vdd.n12171 vdd.n12153 23.783
R39492 vdd.n12172 vdd.n12139 23.783
R39493 vdd.n12172 vdd.n12145 23.783
R39494 vdd.n12173 vdd.n12131 23.783
R39495 vdd.n12173 vdd.n12137 23.783
R39496 vdd.n12174 vdd.n12123 23.783
R39497 vdd.n12174 vdd.n12129 23.783
R39498 vdd.n12175 vdd.n12115 23.783
R39499 vdd.n12175 vdd.n12121 23.783
R39500 vdd.n12176 vdd.n12107 23.783
R39501 vdd.n12176 vdd.n12113 23.783
R39502 vdd.n12177 vdd.n12099 23.783
R39503 vdd.n12177 vdd.n12105 23.783
R39504 vdd.n12178 vdd.n12091 23.783
R39505 vdd.n12178 vdd.n12097 23.783
R39506 vdd.n12179 vdd.n12083 23.783
R39507 vdd.n12179 vdd.n12087 23.783
R39508 vdd.n12180 vdd.n12075 23.783
R39509 vdd.n12180 vdd.n12081 23.783
R39510 vdd.n12181 vdd.n12067 23.783
R39511 vdd.n12181 vdd.n12073 23.783
R39512 vdd.n12182 vdd.n12059 23.783
R39513 vdd.n12182 vdd.n12065 23.783
R39514 vdd.n12183 vdd.n12051 23.783
R39515 vdd.n12183 vdd.n12057 23.783
R39516 vdd.n12184 vdd.n12043 23.783
R39517 vdd.n12184 vdd.n12049 23.783
R39518 vdd.n12185 vdd.n12035 23.783
R39519 vdd.n12185 vdd.n12041 23.783
R39520 vdd.n12186 vdd.n12027 23.783
R39521 vdd.n12186 vdd.n12033 23.783
R39522 vdd.n12187 vdd.n12019 23.783
R39523 vdd.n12187 vdd.n12025 23.783
R39524 vdd.n12198 vdd.n12197 23.783
R39525 vdd.n12198 vdd.n12192 23.783
R39526 vdd.n11989 vdd.n11988 23.783
R39527 vdd.n11989 vdd.n11986 23.783
R39528 vdd.n11990 vdd.n11975 23.783
R39529 vdd.n11990 vdd.n11981 23.783
R39530 vdd.n11991 vdd.n11967 23.783
R39531 vdd.n11991 vdd.n11973 23.783
R39532 vdd.n11992 vdd.n11959 23.783
R39533 vdd.n11992 vdd.n11965 23.783
R39534 vdd.n11993 vdd.n11951 23.783
R39535 vdd.n11993 vdd.n11957 23.783
R39536 vdd.n11994 vdd.n11943 23.783
R39537 vdd.n11994 vdd.n11949 23.783
R39538 vdd.n11995 vdd.n11935 23.783
R39539 vdd.n11995 vdd.n11941 23.783
R39540 vdd.n11996 vdd.n11927 23.783
R39541 vdd.n11996 vdd.n11933 23.783
R39542 vdd.n11997 vdd.n11919 23.783
R39543 vdd.n11997 vdd.n11925 23.783
R39544 vdd.n11998 vdd.n11911 23.783
R39545 vdd.n11998 vdd.n11917 23.783
R39546 vdd.n11999 vdd.n11903 23.783
R39547 vdd.n11999 vdd.n11907 23.783
R39548 vdd.n12000 vdd.n11895 23.783
R39549 vdd.n12000 vdd.n11901 23.783
R39550 vdd.n12001 vdd.n11887 23.783
R39551 vdd.n12001 vdd.n11893 23.783
R39552 vdd.n12002 vdd.n11879 23.783
R39553 vdd.n12002 vdd.n11885 23.783
R39554 vdd.n12003 vdd.n11871 23.783
R39555 vdd.n12003 vdd.n11877 23.783
R39556 vdd.n12004 vdd.n11863 23.783
R39557 vdd.n12004 vdd.n11869 23.783
R39558 vdd.n12005 vdd.n11855 23.783
R39559 vdd.n12005 vdd.n11861 23.783
R39560 vdd.n12006 vdd.n11847 23.783
R39561 vdd.n12006 vdd.n11853 23.783
R39562 vdd.n12007 vdd.n11839 23.783
R39563 vdd.n12007 vdd.n11845 23.783
R39564 vdd.n12018 vdd.n12017 23.783
R39565 vdd.n12018 vdd.n12012 23.783
R39566 vdd.n11809 vdd.n11808 23.783
R39567 vdd.n11809 vdd.n11806 23.783
R39568 vdd.n11810 vdd.n11795 23.783
R39569 vdd.n11810 vdd.n11801 23.783
R39570 vdd.n11811 vdd.n11787 23.783
R39571 vdd.n11811 vdd.n11793 23.783
R39572 vdd.n11812 vdd.n11779 23.783
R39573 vdd.n11812 vdd.n11785 23.783
R39574 vdd.n11813 vdd.n11771 23.783
R39575 vdd.n11813 vdd.n11777 23.783
R39576 vdd.n11814 vdd.n11763 23.783
R39577 vdd.n11814 vdd.n11769 23.783
R39578 vdd.n11815 vdd.n11755 23.783
R39579 vdd.n11815 vdd.n11761 23.783
R39580 vdd.n11816 vdd.n11747 23.783
R39581 vdd.n11816 vdd.n11753 23.783
R39582 vdd.n11817 vdd.n11739 23.783
R39583 vdd.n11817 vdd.n11745 23.783
R39584 vdd.n11818 vdd.n11731 23.783
R39585 vdd.n11818 vdd.n11737 23.783
R39586 vdd.n11819 vdd.n11723 23.783
R39587 vdd.n11819 vdd.n11727 23.783
R39588 vdd.n11820 vdd.n11715 23.783
R39589 vdd.n11820 vdd.n11721 23.783
R39590 vdd.n11821 vdd.n11707 23.783
R39591 vdd.n11821 vdd.n11713 23.783
R39592 vdd.n11822 vdd.n11699 23.783
R39593 vdd.n11822 vdd.n11705 23.783
R39594 vdd.n11823 vdd.n11691 23.783
R39595 vdd.n11823 vdd.n11697 23.783
R39596 vdd.n11824 vdd.n11683 23.783
R39597 vdd.n11824 vdd.n11689 23.783
R39598 vdd.n11825 vdd.n11675 23.783
R39599 vdd.n11825 vdd.n11681 23.783
R39600 vdd.n11826 vdd.n11667 23.783
R39601 vdd.n11826 vdd.n11673 23.783
R39602 vdd.n11827 vdd.n11659 23.783
R39603 vdd.n11827 vdd.n11665 23.783
R39604 vdd.n11838 vdd.n11837 23.783
R39605 vdd.n11838 vdd.n11832 23.783
R39606 vdd.n11629 vdd.n11628 23.783
R39607 vdd.n11629 vdd.n11626 23.783
R39608 vdd.n11630 vdd.n11615 23.783
R39609 vdd.n11630 vdd.n11621 23.783
R39610 vdd.n11631 vdd.n11607 23.783
R39611 vdd.n11631 vdd.n11613 23.783
R39612 vdd.n11632 vdd.n11599 23.783
R39613 vdd.n11632 vdd.n11605 23.783
R39614 vdd.n11633 vdd.n11591 23.783
R39615 vdd.n11633 vdd.n11597 23.783
R39616 vdd.n11634 vdd.n11583 23.783
R39617 vdd.n11634 vdd.n11589 23.783
R39618 vdd.n11635 vdd.n11575 23.783
R39619 vdd.n11635 vdd.n11581 23.783
R39620 vdd.n11636 vdd.n11567 23.783
R39621 vdd.n11636 vdd.n11573 23.783
R39622 vdd.n11637 vdd.n11559 23.783
R39623 vdd.n11637 vdd.n11565 23.783
R39624 vdd.n11638 vdd.n11551 23.783
R39625 vdd.n11638 vdd.n11557 23.783
R39626 vdd.n11639 vdd.n11543 23.783
R39627 vdd.n11639 vdd.n11547 23.783
R39628 vdd.n11640 vdd.n11535 23.783
R39629 vdd.n11640 vdd.n11541 23.783
R39630 vdd.n11641 vdd.n11527 23.783
R39631 vdd.n11641 vdd.n11533 23.783
R39632 vdd.n11642 vdd.n11519 23.783
R39633 vdd.n11642 vdd.n11525 23.783
R39634 vdd.n11643 vdd.n11511 23.783
R39635 vdd.n11643 vdd.n11517 23.783
R39636 vdd.n11644 vdd.n11503 23.783
R39637 vdd.n11644 vdd.n11509 23.783
R39638 vdd.n11645 vdd.n11495 23.783
R39639 vdd.n11645 vdd.n11501 23.783
R39640 vdd.n11646 vdd.n11487 23.783
R39641 vdd.n11646 vdd.n11493 23.783
R39642 vdd.n11647 vdd.n11479 23.783
R39643 vdd.n11647 vdd.n11485 23.783
R39644 vdd.n11658 vdd.n11657 23.783
R39645 vdd.n11658 vdd.n11652 23.783
R39646 vdd.n150 vdd.n149 23.783
R39647 vdd.n150 vdd.n147 23.783
R39648 vdd.n151 vdd.n136 23.783
R39649 vdd.n151 vdd.n142 23.783
R39650 vdd.n152 vdd.n128 23.783
R39651 vdd.n152 vdd.n134 23.783
R39652 vdd.n153 vdd.n120 23.783
R39653 vdd.n153 vdd.n126 23.783
R39654 vdd.n154 vdd.n112 23.783
R39655 vdd.n154 vdd.n118 23.783
R39656 vdd.n155 vdd.n104 23.783
R39657 vdd.n155 vdd.n110 23.783
R39658 vdd.n156 vdd.n96 23.783
R39659 vdd.n156 vdd.n102 23.783
R39660 vdd.n157 vdd.n88 23.783
R39661 vdd.n157 vdd.n94 23.783
R39662 vdd.n158 vdd.n80 23.783
R39663 vdd.n158 vdd.n86 23.783
R39664 vdd.n159 vdd.n72 23.783
R39665 vdd.n159 vdd.n78 23.783
R39666 vdd.n160 vdd.n64 23.783
R39667 vdd.n160 vdd.n68 23.783
R39668 vdd.n161 vdd.n56 23.783
R39669 vdd.n161 vdd.n62 23.783
R39670 vdd.n162 vdd.n48 23.783
R39671 vdd.n162 vdd.n54 23.783
R39672 vdd.n163 vdd.n40 23.783
R39673 vdd.n163 vdd.n46 23.783
R39674 vdd.n164 vdd.n32 23.783
R39675 vdd.n164 vdd.n38 23.783
R39676 vdd.n165 vdd.n24 23.783
R39677 vdd.n165 vdd.n30 23.783
R39678 vdd.n166 vdd.n16 23.783
R39679 vdd.n166 vdd.n22 23.783
R39680 vdd.n167 vdd.n8 23.783
R39681 vdd.n167 vdd.n14 23.783
R39682 vdd.n168 vdd.n0 23.783
R39683 vdd.n168 vdd.n6 23.783
R39684 vdd.n179 vdd.n178 23.783
R39685 vdd.n179 vdd.n173 23.783
R39686 vdd.n330 vdd.n329 23.783
R39687 vdd.n330 vdd.n327 23.783
R39688 vdd.n331 vdd.n316 23.783
R39689 vdd.n331 vdd.n322 23.783
R39690 vdd.n332 vdd.n308 23.783
R39691 vdd.n332 vdd.n314 23.783
R39692 vdd.n333 vdd.n300 23.783
R39693 vdd.n333 vdd.n306 23.783
R39694 vdd.n334 vdd.n292 23.783
R39695 vdd.n334 vdd.n298 23.783
R39696 vdd.n335 vdd.n284 23.783
R39697 vdd.n335 vdd.n290 23.783
R39698 vdd.n336 vdd.n276 23.783
R39699 vdd.n336 vdd.n282 23.783
R39700 vdd.n337 vdd.n268 23.783
R39701 vdd.n337 vdd.n274 23.783
R39702 vdd.n338 vdd.n260 23.783
R39703 vdd.n338 vdd.n266 23.783
R39704 vdd.n339 vdd.n252 23.783
R39705 vdd.n339 vdd.n258 23.783
R39706 vdd.n340 vdd.n244 23.783
R39707 vdd.n340 vdd.n248 23.783
R39708 vdd.n341 vdd.n236 23.783
R39709 vdd.n341 vdd.n242 23.783
R39710 vdd.n342 vdd.n228 23.783
R39711 vdd.n342 vdd.n234 23.783
R39712 vdd.n343 vdd.n220 23.783
R39713 vdd.n343 vdd.n226 23.783
R39714 vdd.n344 vdd.n212 23.783
R39715 vdd.n344 vdd.n218 23.783
R39716 vdd.n345 vdd.n204 23.783
R39717 vdd.n345 vdd.n210 23.783
R39718 vdd.n346 vdd.n196 23.783
R39719 vdd.n346 vdd.n202 23.783
R39720 vdd.n347 vdd.n188 23.783
R39721 vdd.n347 vdd.n194 23.783
R39722 vdd.n348 vdd.n180 23.783
R39723 vdd.n348 vdd.n186 23.783
R39724 vdd.n359 vdd.n358 23.783
R39725 vdd.n359 vdd.n353 23.783
R39726 vdd.n510 vdd.n509 23.783
R39727 vdd.n510 vdd.n507 23.783
R39728 vdd.n511 vdd.n496 23.783
R39729 vdd.n511 vdd.n502 23.783
R39730 vdd.n512 vdd.n488 23.783
R39731 vdd.n512 vdd.n494 23.783
R39732 vdd.n513 vdd.n480 23.783
R39733 vdd.n513 vdd.n486 23.783
R39734 vdd.n514 vdd.n472 23.783
R39735 vdd.n514 vdd.n478 23.783
R39736 vdd.n515 vdd.n464 23.783
R39737 vdd.n515 vdd.n470 23.783
R39738 vdd.n516 vdd.n456 23.783
R39739 vdd.n516 vdd.n462 23.783
R39740 vdd.n517 vdd.n448 23.783
R39741 vdd.n517 vdd.n454 23.783
R39742 vdd.n518 vdd.n440 23.783
R39743 vdd.n518 vdd.n446 23.783
R39744 vdd.n519 vdd.n432 23.783
R39745 vdd.n519 vdd.n438 23.783
R39746 vdd.n520 vdd.n424 23.783
R39747 vdd.n520 vdd.n428 23.783
R39748 vdd.n521 vdd.n416 23.783
R39749 vdd.n521 vdd.n422 23.783
R39750 vdd.n522 vdd.n408 23.783
R39751 vdd.n522 vdd.n414 23.783
R39752 vdd.n523 vdd.n400 23.783
R39753 vdd.n523 vdd.n406 23.783
R39754 vdd.n524 vdd.n392 23.783
R39755 vdd.n524 vdd.n398 23.783
R39756 vdd.n525 vdd.n384 23.783
R39757 vdd.n525 vdd.n390 23.783
R39758 vdd.n526 vdd.n376 23.783
R39759 vdd.n526 vdd.n382 23.783
R39760 vdd.n527 vdd.n368 23.783
R39761 vdd.n527 vdd.n374 23.783
R39762 vdd.n528 vdd.n360 23.783
R39763 vdd.n528 vdd.n366 23.783
R39764 vdd.n539 vdd.n538 23.783
R39765 vdd.n539 vdd.n533 23.783
R39766 vdd.n690 vdd.n689 23.783
R39767 vdd.n690 vdd.n687 23.783
R39768 vdd.n691 vdd.n676 23.783
R39769 vdd.n691 vdd.n682 23.783
R39770 vdd.n692 vdd.n668 23.783
R39771 vdd.n692 vdd.n674 23.783
R39772 vdd.n693 vdd.n660 23.783
R39773 vdd.n693 vdd.n666 23.783
R39774 vdd.n694 vdd.n652 23.783
R39775 vdd.n694 vdd.n658 23.783
R39776 vdd.n695 vdd.n644 23.783
R39777 vdd.n695 vdd.n650 23.783
R39778 vdd.n696 vdd.n636 23.783
R39779 vdd.n696 vdd.n642 23.783
R39780 vdd.n697 vdd.n628 23.783
R39781 vdd.n697 vdd.n634 23.783
R39782 vdd.n698 vdd.n620 23.783
R39783 vdd.n698 vdd.n626 23.783
R39784 vdd.n699 vdd.n612 23.783
R39785 vdd.n699 vdd.n618 23.783
R39786 vdd.n700 vdd.n604 23.783
R39787 vdd.n700 vdd.n608 23.783
R39788 vdd.n701 vdd.n596 23.783
R39789 vdd.n701 vdd.n602 23.783
R39790 vdd.n702 vdd.n588 23.783
R39791 vdd.n702 vdd.n594 23.783
R39792 vdd.n703 vdd.n580 23.783
R39793 vdd.n703 vdd.n586 23.783
R39794 vdd.n704 vdd.n572 23.783
R39795 vdd.n704 vdd.n578 23.783
R39796 vdd.n705 vdd.n564 23.783
R39797 vdd.n705 vdd.n570 23.783
R39798 vdd.n706 vdd.n556 23.783
R39799 vdd.n706 vdd.n562 23.783
R39800 vdd.n707 vdd.n548 23.783
R39801 vdd.n707 vdd.n554 23.783
R39802 vdd.n708 vdd.n540 23.783
R39803 vdd.n708 vdd.n546 23.783
R39804 vdd.n719 vdd.n718 23.783
R39805 vdd.n719 vdd.n713 23.783
R39806 vdd.n870 vdd.n869 23.783
R39807 vdd.n870 vdd.n867 23.783
R39808 vdd.n871 vdd.n856 23.783
R39809 vdd.n871 vdd.n862 23.783
R39810 vdd.n872 vdd.n848 23.783
R39811 vdd.n872 vdd.n854 23.783
R39812 vdd.n873 vdd.n840 23.783
R39813 vdd.n873 vdd.n846 23.783
R39814 vdd.n874 vdd.n832 23.783
R39815 vdd.n874 vdd.n838 23.783
R39816 vdd.n875 vdd.n824 23.783
R39817 vdd.n875 vdd.n830 23.783
R39818 vdd.n876 vdd.n816 23.783
R39819 vdd.n876 vdd.n822 23.783
R39820 vdd.n877 vdd.n808 23.783
R39821 vdd.n877 vdd.n814 23.783
R39822 vdd.n878 vdd.n800 23.783
R39823 vdd.n878 vdd.n806 23.783
R39824 vdd.n879 vdd.n792 23.783
R39825 vdd.n879 vdd.n798 23.783
R39826 vdd.n880 vdd.n784 23.783
R39827 vdd.n880 vdd.n788 23.783
R39828 vdd.n881 vdd.n776 23.783
R39829 vdd.n881 vdd.n782 23.783
R39830 vdd.n882 vdd.n768 23.783
R39831 vdd.n882 vdd.n774 23.783
R39832 vdd.n883 vdd.n760 23.783
R39833 vdd.n883 vdd.n766 23.783
R39834 vdd.n884 vdd.n752 23.783
R39835 vdd.n884 vdd.n758 23.783
R39836 vdd.n885 vdd.n744 23.783
R39837 vdd.n885 vdd.n750 23.783
R39838 vdd.n886 vdd.n736 23.783
R39839 vdd.n886 vdd.n742 23.783
R39840 vdd.n887 vdd.n728 23.783
R39841 vdd.n887 vdd.n734 23.783
R39842 vdd.n888 vdd.n720 23.783
R39843 vdd.n888 vdd.n726 23.783
R39844 vdd.n899 vdd.n898 23.783
R39845 vdd.n899 vdd.n893 23.783
R39846 vdd.n1050 vdd.n1049 23.783
R39847 vdd.n1050 vdd.n1047 23.783
R39848 vdd.n1051 vdd.n1036 23.783
R39849 vdd.n1051 vdd.n1042 23.783
R39850 vdd.n1052 vdd.n1028 23.783
R39851 vdd.n1052 vdd.n1034 23.783
R39852 vdd.n1053 vdd.n1020 23.783
R39853 vdd.n1053 vdd.n1026 23.783
R39854 vdd.n1054 vdd.n1012 23.783
R39855 vdd.n1054 vdd.n1018 23.783
R39856 vdd.n1055 vdd.n1004 23.783
R39857 vdd.n1055 vdd.n1010 23.783
R39858 vdd.n1056 vdd.n996 23.783
R39859 vdd.n1056 vdd.n1002 23.783
R39860 vdd.n1057 vdd.n988 23.783
R39861 vdd.n1057 vdd.n994 23.783
R39862 vdd.n1058 vdd.n980 23.783
R39863 vdd.n1058 vdd.n986 23.783
R39864 vdd.n1059 vdd.n972 23.783
R39865 vdd.n1059 vdd.n978 23.783
R39866 vdd.n1060 vdd.n964 23.783
R39867 vdd.n1060 vdd.n968 23.783
R39868 vdd.n1061 vdd.n956 23.783
R39869 vdd.n1061 vdd.n962 23.783
R39870 vdd.n1062 vdd.n948 23.783
R39871 vdd.n1062 vdd.n954 23.783
R39872 vdd.n1063 vdd.n940 23.783
R39873 vdd.n1063 vdd.n946 23.783
R39874 vdd.n1064 vdd.n932 23.783
R39875 vdd.n1064 vdd.n938 23.783
R39876 vdd.n1065 vdd.n924 23.783
R39877 vdd.n1065 vdd.n930 23.783
R39878 vdd.n1066 vdd.n916 23.783
R39879 vdd.n1066 vdd.n922 23.783
R39880 vdd.n1067 vdd.n908 23.783
R39881 vdd.n1067 vdd.n914 23.783
R39882 vdd.n1068 vdd.n900 23.783
R39883 vdd.n1068 vdd.n906 23.783
R39884 vdd.n1079 vdd.n1078 23.783
R39885 vdd.n1079 vdd.n1073 23.783
R39886 vdd.n1230 vdd.n1229 23.783
R39887 vdd.n1230 vdd.n1227 23.783
R39888 vdd.n1231 vdd.n1216 23.783
R39889 vdd.n1231 vdd.n1222 23.783
R39890 vdd.n1232 vdd.n1208 23.783
R39891 vdd.n1232 vdd.n1214 23.783
R39892 vdd.n1233 vdd.n1200 23.783
R39893 vdd.n1233 vdd.n1206 23.783
R39894 vdd.n1234 vdd.n1192 23.783
R39895 vdd.n1234 vdd.n1198 23.783
R39896 vdd.n1235 vdd.n1184 23.783
R39897 vdd.n1235 vdd.n1190 23.783
R39898 vdd.n1236 vdd.n1176 23.783
R39899 vdd.n1236 vdd.n1182 23.783
R39900 vdd.n1237 vdd.n1168 23.783
R39901 vdd.n1237 vdd.n1174 23.783
R39902 vdd.n1238 vdd.n1160 23.783
R39903 vdd.n1238 vdd.n1166 23.783
R39904 vdd.n1239 vdd.n1152 23.783
R39905 vdd.n1239 vdd.n1158 23.783
R39906 vdd.n1240 vdd.n1144 23.783
R39907 vdd.n1240 vdd.n1148 23.783
R39908 vdd.n1241 vdd.n1136 23.783
R39909 vdd.n1241 vdd.n1142 23.783
R39910 vdd.n1242 vdd.n1128 23.783
R39911 vdd.n1242 vdd.n1134 23.783
R39912 vdd.n1243 vdd.n1120 23.783
R39913 vdd.n1243 vdd.n1126 23.783
R39914 vdd.n1244 vdd.n1112 23.783
R39915 vdd.n1244 vdd.n1118 23.783
R39916 vdd.n1245 vdd.n1104 23.783
R39917 vdd.n1245 vdd.n1110 23.783
R39918 vdd.n1246 vdd.n1096 23.783
R39919 vdd.n1246 vdd.n1102 23.783
R39920 vdd.n1247 vdd.n1088 23.783
R39921 vdd.n1247 vdd.n1094 23.783
R39922 vdd.n1248 vdd.n1080 23.783
R39923 vdd.n1248 vdd.n1086 23.783
R39924 vdd.n1259 vdd.n1258 23.783
R39925 vdd.n1259 vdd.n1253 23.783
R39926 vdd.n1410 vdd.n1409 23.783
R39927 vdd.n1410 vdd.n1407 23.783
R39928 vdd.n1411 vdd.n1396 23.783
R39929 vdd.n1411 vdd.n1402 23.783
R39930 vdd.n1412 vdd.n1388 23.783
R39931 vdd.n1412 vdd.n1394 23.783
R39932 vdd.n1413 vdd.n1380 23.783
R39933 vdd.n1413 vdd.n1386 23.783
R39934 vdd.n1414 vdd.n1372 23.783
R39935 vdd.n1414 vdd.n1378 23.783
R39936 vdd.n1415 vdd.n1364 23.783
R39937 vdd.n1415 vdd.n1370 23.783
R39938 vdd.n1416 vdd.n1356 23.783
R39939 vdd.n1416 vdd.n1362 23.783
R39940 vdd.n1417 vdd.n1348 23.783
R39941 vdd.n1417 vdd.n1354 23.783
R39942 vdd.n1418 vdd.n1340 23.783
R39943 vdd.n1418 vdd.n1346 23.783
R39944 vdd.n1419 vdd.n1332 23.783
R39945 vdd.n1419 vdd.n1338 23.783
R39946 vdd.n1420 vdd.n1324 23.783
R39947 vdd.n1420 vdd.n1328 23.783
R39948 vdd.n1421 vdd.n1316 23.783
R39949 vdd.n1421 vdd.n1322 23.783
R39950 vdd.n1422 vdd.n1308 23.783
R39951 vdd.n1422 vdd.n1314 23.783
R39952 vdd.n1423 vdd.n1300 23.783
R39953 vdd.n1423 vdd.n1306 23.783
R39954 vdd.n1424 vdd.n1292 23.783
R39955 vdd.n1424 vdd.n1298 23.783
R39956 vdd.n1425 vdd.n1284 23.783
R39957 vdd.n1425 vdd.n1290 23.783
R39958 vdd.n1426 vdd.n1276 23.783
R39959 vdd.n1426 vdd.n1282 23.783
R39960 vdd.n1427 vdd.n1268 23.783
R39961 vdd.n1427 vdd.n1274 23.783
R39962 vdd.n1428 vdd.n1260 23.783
R39963 vdd.n1428 vdd.n1266 23.783
R39964 vdd.n1439 vdd.n1438 23.783
R39965 vdd.n1439 vdd.n1433 23.783
R39966 vdd.n1590 vdd.n1589 23.783
R39967 vdd.n1590 vdd.n1587 23.783
R39968 vdd.n1591 vdd.n1576 23.783
R39969 vdd.n1591 vdd.n1582 23.783
R39970 vdd.n1592 vdd.n1568 23.783
R39971 vdd.n1592 vdd.n1574 23.783
R39972 vdd.n1593 vdd.n1560 23.783
R39973 vdd.n1593 vdd.n1566 23.783
R39974 vdd.n1594 vdd.n1552 23.783
R39975 vdd.n1594 vdd.n1558 23.783
R39976 vdd.n1595 vdd.n1544 23.783
R39977 vdd.n1595 vdd.n1550 23.783
R39978 vdd.n1596 vdd.n1536 23.783
R39979 vdd.n1596 vdd.n1542 23.783
R39980 vdd.n1597 vdd.n1528 23.783
R39981 vdd.n1597 vdd.n1534 23.783
R39982 vdd.n1598 vdd.n1520 23.783
R39983 vdd.n1598 vdd.n1526 23.783
R39984 vdd.n1599 vdd.n1512 23.783
R39985 vdd.n1599 vdd.n1518 23.783
R39986 vdd.n1600 vdd.n1504 23.783
R39987 vdd.n1600 vdd.n1508 23.783
R39988 vdd.n1601 vdd.n1496 23.783
R39989 vdd.n1601 vdd.n1502 23.783
R39990 vdd.n1602 vdd.n1488 23.783
R39991 vdd.n1602 vdd.n1494 23.783
R39992 vdd.n1603 vdd.n1480 23.783
R39993 vdd.n1603 vdd.n1486 23.783
R39994 vdd.n1604 vdd.n1472 23.783
R39995 vdd.n1604 vdd.n1478 23.783
R39996 vdd.n1605 vdd.n1464 23.783
R39997 vdd.n1605 vdd.n1470 23.783
R39998 vdd.n1606 vdd.n1456 23.783
R39999 vdd.n1606 vdd.n1462 23.783
R40000 vdd.n1607 vdd.n1448 23.783
R40001 vdd.n1607 vdd.n1454 23.783
R40002 vdd.n1608 vdd.n1440 23.783
R40003 vdd.n1608 vdd.n1446 23.783
R40004 vdd.n1619 vdd.n1618 23.783
R40005 vdd.n1619 vdd.n1613 23.783
R40006 vdd.n1770 vdd.n1769 23.783
R40007 vdd.n1770 vdd.n1767 23.783
R40008 vdd.n1771 vdd.n1756 23.783
R40009 vdd.n1771 vdd.n1762 23.783
R40010 vdd.n1772 vdd.n1748 23.783
R40011 vdd.n1772 vdd.n1754 23.783
R40012 vdd.n1773 vdd.n1740 23.783
R40013 vdd.n1773 vdd.n1746 23.783
R40014 vdd.n1774 vdd.n1732 23.783
R40015 vdd.n1774 vdd.n1738 23.783
R40016 vdd.n1775 vdd.n1724 23.783
R40017 vdd.n1775 vdd.n1730 23.783
R40018 vdd.n1776 vdd.n1716 23.783
R40019 vdd.n1776 vdd.n1722 23.783
R40020 vdd.n1777 vdd.n1708 23.783
R40021 vdd.n1777 vdd.n1714 23.783
R40022 vdd.n1778 vdd.n1700 23.783
R40023 vdd.n1778 vdd.n1706 23.783
R40024 vdd.n1779 vdd.n1692 23.783
R40025 vdd.n1779 vdd.n1698 23.783
R40026 vdd.n1780 vdd.n1684 23.783
R40027 vdd.n1780 vdd.n1688 23.783
R40028 vdd.n1781 vdd.n1676 23.783
R40029 vdd.n1781 vdd.n1682 23.783
R40030 vdd.n1782 vdd.n1668 23.783
R40031 vdd.n1782 vdd.n1674 23.783
R40032 vdd.n1783 vdd.n1660 23.783
R40033 vdd.n1783 vdd.n1666 23.783
R40034 vdd.n1784 vdd.n1652 23.783
R40035 vdd.n1784 vdd.n1658 23.783
R40036 vdd.n1785 vdd.n1644 23.783
R40037 vdd.n1785 vdd.n1650 23.783
R40038 vdd.n1786 vdd.n1636 23.783
R40039 vdd.n1786 vdd.n1642 23.783
R40040 vdd.n1787 vdd.n1628 23.783
R40041 vdd.n1787 vdd.n1634 23.783
R40042 vdd.n1788 vdd.n1620 23.783
R40043 vdd.n1788 vdd.n1626 23.783
R40044 vdd.n1799 vdd.n1798 23.783
R40045 vdd.n1799 vdd.n1793 23.783
R40046 vdd.n1950 vdd.n1949 23.783
R40047 vdd.n1950 vdd.n1947 23.783
R40048 vdd.n1951 vdd.n1936 23.783
R40049 vdd.n1951 vdd.n1942 23.783
R40050 vdd.n1952 vdd.n1928 23.783
R40051 vdd.n1952 vdd.n1934 23.783
R40052 vdd.n1953 vdd.n1920 23.783
R40053 vdd.n1953 vdd.n1926 23.783
R40054 vdd.n1954 vdd.n1912 23.783
R40055 vdd.n1954 vdd.n1918 23.783
R40056 vdd.n1955 vdd.n1904 23.783
R40057 vdd.n1955 vdd.n1910 23.783
R40058 vdd.n1956 vdd.n1896 23.783
R40059 vdd.n1956 vdd.n1902 23.783
R40060 vdd.n1957 vdd.n1888 23.783
R40061 vdd.n1957 vdd.n1894 23.783
R40062 vdd.n1958 vdd.n1880 23.783
R40063 vdd.n1958 vdd.n1886 23.783
R40064 vdd.n1959 vdd.n1872 23.783
R40065 vdd.n1959 vdd.n1878 23.783
R40066 vdd.n1960 vdd.n1864 23.783
R40067 vdd.n1960 vdd.n1868 23.783
R40068 vdd.n1961 vdd.n1856 23.783
R40069 vdd.n1961 vdd.n1862 23.783
R40070 vdd.n1962 vdd.n1848 23.783
R40071 vdd.n1962 vdd.n1854 23.783
R40072 vdd.n1963 vdd.n1840 23.783
R40073 vdd.n1963 vdd.n1846 23.783
R40074 vdd.n1964 vdd.n1832 23.783
R40075 vdd.n1964 vdd.n1838 23.783
R40076 vdd.n1965 vdd.n1824 23.783
R40077 vdd.n1965 vdd.n1830 23.783
R40078 vdd.n1966 vdd.n1816 23.783
R40079 vdd.n1966 vdd.n1822 23.783
R40080 vdd.n1967 vdd.n1808 23.783
R40081 vdd.n1967 vdd.n1814 23.783
R40082 vdd.n1968 vdd.n1800 23.783
R40083 vdd.n1968 vdd.n1806 23.783
R40084 vdd.n1979 vdd.n1978 23.783
R40085 vdd.n1979 vdd.n1973 23.783
R40086 vdd.n2130 vdd.n2129 23.783
R40087 vdd.n2130 vdd.n2127 23.783
R40088 vdd.n2131 vdd.n2116 23.783
R40089 vdd.n2131 vdd.n2122 23.783
R40090 vdd.n2132 vdd.n2108 23.783
R40091 vdd.n2132 vdd.n2114 23.783
R40092 vdd.n2133 vdd.n2100 23.783
R40093 vdd.n2133 vdd.n2106 23.783
R40094 vdd.n2134 vdd.n2092 23.783
R40095 vdd.n2134 vdd.n2098 23.783
R40096 vdd.n2135 vdd.n2084 23.783
R40097 vdd.n2135 vdd.n2090 23.783
R40098 vdd.n2136 vdd.n2076 23.783
R40099 vdd.n2136 vdd.n2082 23.783
R40100 vdd.n2137 vdd.n2068 23.783
R40101 vdd.n2137 vdd.n2074 23.783
R40102 vdd.n2138 vdd.n2060 23.783
R40103 vdd.n2138 vdd.n2066 23.783
R40104 vdd.n2139 vdd.n2052 23.783
R40105 vdd.n2139 vdd.n2058 23.783
R40106 vdd.n2140 vdd.n2044 23.783
R40107 vdd.n2140 vdd.n2048 23.783
R40108 vdd.n2141 vdd.n2036 23.783
R40109 vdd.n2141 vdd.n2042 23.783
R40110 vdd.n2142 vdd.n2028 23.783
R40111 vdd.n2142 vdd.n2034 23.783
R40112 vdd.n2143 vdd.n2020 23.783
R40113 vdd.n2143 vdd.n2026 23.783
R40114 vdd.n2144 vdd.n2012 23.783
R40115 vdd.n2144 vdd.n2018 23.783
R40116 vdd.n2145 vdd.n2004 23.783
R40117 vdd.n2145 vdd.n2010 23.783
R40118 vdd.n2146 vdd.n1996 23.783
R40119 vdd.n2146 vdd.n2002 23.783
R40120 vdd.n2147 vdd.n1988 23.783
R40121 vdd.n2147 vdd.n1994 23.783
R40122 vdd.n2148 vdd.n1980 23.783
R40123 vdd.n2148 vdd.n1986 23.783
R40124 vdd.n2159 vdd.n2158 23.783
R40125 vdd.n2159 vdd.n2153 23.783
R40126 vdd.n2310 vdd.n2309 23.783
R40127 vdd.n2310 vdd.n2307 23.783
R40128 vdd.n2311 vdd.n2296 23.783
R40129 vdd.n2311 vdd.n2302 23.783
R40130 vdd.n2312 vdd.n2288 23.783
R40131 vdd.n2312 vdd.n2294 23.783
R40132 vdd.n2313 vdd.n2280 23.783
R40133 vdd.n2313 vdd.n2286 23.783
R40134 vdd.n2314 vdd.n2272 23.783
R40135 vdd.n2314 vdd.n2278 23.783
R40136 vdd.n2315 vdd.n2264 23.783
R40137 vdd.n2315 vdd.n2270 23.783
R40138 vdd.n2316 vdd.n2256 23.783
R40139 vdd.n2316 vdd.n2262 23.783
R40140 vdd.n2317 vdd.n2248 23.783
R40141 vdd.n2317 vdd.n2254 23.783
R40142 vdd.n2318 vdd.n2240 23.783
R40143 vdd.n2318 vdd.n2246 23.783
R40144 vdd.n2319 vdd.n2232 23.783
R40145 vdd.n2319 vdd.n2238 23.783
R40146 vdd.n2320 vdd.n2224 23.783
R40147 vdd.n2320 vdd.n2228 23.783
R40148 vdd.n2321 vdd.n2216 23.783
R40149 vdd.n2321 vdd.n2222 23.783
R40150 vdd.n2322 vdd.n2208 23.783
R40151 vdd.n2322 vdd.n2214 23.783
R40152 vdd.n2323 vdd.n2200 23.783
R40153 vdd.n2323 vdd.n2206 23.783
R40154 vdd.n2324 vdd.n2192 23.783
R40155 vdd.n2324 vdd.n2198 23.783
R40156 vdd.n2325 vdd.n2184 23.783
R40157 vdd.n2325 vdd.n2190 23.783
R40158 vdd.n2326 vdd.n2176 23.783
R40159 vdd.n2326 vdd.n2182 23.783
R40160 vdd.n2327 vdd.n2168 23.783
R40161 vdd.n2327 vdd.n2174 23.783
R40162 vdd.n2328 vdd.n2160 23.783
R40163 vdd.n2328 vdd.n2166 23.783
R40164 vdd.n2339 vdd.n2338 23.783
R40165 vdd.n2339 vdd.n2333 23.783
R40166 vdd.n2490 vdd.n2489 23.783
R40167 vdd.n2490 vdd.n2487 23.783
R40168 vdd.n2491 vdd.n2476 23.783
R40169 vdd.n2491 vdd.n2482 23.783
R40170 vdd.n2492 vdd.n2468 23.783
R40171 vdd.n2492 vdd.n2474 23.783
R40172 vdd.n2493 vdd.n2460 23.783
R40173 vdd.n2493 vdd.n2466 23.783
R40174 vdd.n2494 vdd.n2452 23.783
R40175 vdd.n2494 vdd.n2458 23.783
R40176 vdd.n2495 vdd.n2444 23.783
R40177 vdd.n2495 vdd.n2450 23.783
R40178 vdd.n2496 vdd.n2436 23.783
R40179 vdd.n2496 vdd.n2442 23.783
R40180 vdd.n2497 vdd.n2428 23.783
R40181 vdd.n2497 vdd.n2434 23.783
R40182 vdd.n2498 vdd.n2420 23.783
R40183 vdd.n2498 vdd.n2426 23.783
R40184 vdd.n2499 vdd.n2412 23.783
R40185 vdd.n2499 vdd.n2418 23.783
R40186 vdd.n2500 vdd.n2404 23.783
R40187 vdd.n2500 vdd.n2408 23.783
R40188 vdd.n2501 vdd.n2396 23.783
R40189 vdd.n2501 vdd.n2402 23.783
R40190 vdd.n2502 vdd.n2388 23.783
R40191 vdd.n2502 vdd.n2394 23.783
R40192 vdd.n2503 vdd.n2380 23.783
R40193 vdd.n2503 vdd.n2386 23.783
R40194 vdd.n2504 vdd.n2372 23.783
R40195 vdd.n2504 vdd.n2378 23.783
R40196 vdd.n2505 vdd.n2364 23.783
R40197 vdd.n2505 vdd.n2370 23.783
R40198 vdd.n2506 vdd.n2356 23.783
R40199 vdd.n2506 vdd.n2362 23.783
R40200 vdd.n2507 vdd.n2348 23.783
R40201 vdd.n2507 vdd.n2354 23.783
R40202 vdd.n2508 vdd.n2340 23.783
R40203 vdd.n2508 vdd.n2346 23.783
R40204 vdd.n2519 vdd.n2518 23.783
R40205 vdd.n2519 vdd.n2513 23.783
R40206 vdd.n2670 vdd.n2669 23.783
R40207 vdd.n2670 vdd.n2667 23.783
R40208 vdd.n2671 vdd.n2656 23.783
R40209 vdd.n2671 vdd.n2662 23.783
R40210 vdd.n2672 vdd.n2648 23.783
R40211 vdd.n2672 vdd.n2654 23.783
R40212 vdd.n2673 vdd.n2640 23.783
R40213 vdd.n2673 vdd.n2646 23.783
R40214 vdd.n2674 vdd.n2632 23.783
R40215 vdd.n2674 vdd.n2638 23.783
R40216 vdd.n2675 vdd.n2624 23.783
R40217 vdd.n2675 vdd.n2630 23.783
R40218 vdd.n2676 vdd.n2616 23.783
R40219 vdd.n2676 vdd.n2622 23.783
R40220 vdd.n2677 vdd.n2608 23.783
R40221 vdd.n2677 vdd.n2614 23.783
R40222 vdd.n2678 vdd.n2600 23.783
R40223 vdd.n2678 vdd.n2606 23.783
R40224 vdd.n2679 vdd.n2592 23.783
R40225 vdd.n2679 vdd.n2598 23.783
R40226 vdd.n2680 vdd.n2584 23.783
R40227 vdd.n2680 vdd.n2588 23.783
R40228 vdd.n2681 vdd.n2576 23.783
R40229 vdd.n2681 vdd.n2582 23.783
R40230 vdd.n2682 vdd.n2568 23.783
R40231 vdd.n2682 vdd.n2574 23.783
R40232 vdd.n2683 vdd.n2560 23.783
R40233 vdd.n2683 vdd.n2566 23.783
R40234 vdd.n2684 vdd.n2552 23.783
R40235 vdd.n2684 vdd.n2558 23.783
R40236 vdd.n2685 vdd.n2544 23.783
R40237 vdd.n2685 vdd.n2550 23.783
R40238 vdd.n2686 vdd.n2536 23.783
R40239 vdd.n2686 vdd.n2542 23.783
R40240 vdd.n2687 vdd.n2528 23.783
R40241 vdd.n2687 vdd.n2534 23.783
R40242 vdd.n2688 vdd.n2520 23.783
R40243 vdd.n2688 vdd.n2526 23.783
R40244 vdd.n2699 vdd.n2698 23.783
R40245 vdd.n2699 vdd.n2693 23.783
R40246 vdd.n2850 vdd.n2849 23.783
R40247 vdd.n2850 vdd.n2847 23.783
R40248 vdd.n2851 vdd.n2836 23.783
R40249 vdd.n2851 vdd.n2842 23.783
R40250 vdd.n2852 vdd.n2828 23.783
R40251 vdd.n2852 vdd.n2834 23.783
R40252 vdd.n2853 vdd.n2820 23.783
R40253 vdd.n2853 vdd.n2826 23.783
R40254 vdd.n2854 vdd.n2812 23.783
R40255 vdd.n2854 vdd.n2818 23.783
R40256 vdd.n2855 vdd.n2804 23.783
R40257 vdd.n2855 vdd.n2810 23.783
R40258 vdd.n2856 vdd.n2796 23.783
R40259 vdd.n2856 vdd.n2802 23.783
R40260 vdd.n2857 vdd.n2788 23.783
R40261 vdd.n2857 vdd.n2794 23.783
R40262 vdd.n2858 vdd.n2780 23.783
R40263 vdd.n2858 vdd.n2786 23.783
R40264 vdd.n2859 vdd.n2772 23.783
R40265 vdd.n2859 vdd.n2778 23.783
R40266 vdd.n2860 vdd.n2764 23.783
R40267 vdd.n2860 vdd.n2768 23.783
R40268 vdd.n2861 vdd.n2756 23.783
R40269 vdd.n2861 vdd.n2762 23.783
R40270 vdd.n2862 vdd.n2748 23.783
R40271 vdd.n2862 vdd.n2754 23.783
R40272 vdd.n2863 vdd.n2740 23.783
R40273 vdd.n2863 vdd.n2746 23.783
R40274 vdd.n2864 vdd.n2732 23.783
R40275 vdd.n2864 vdd.n2738 23.783
R40276 vdd.n2865 vdd.n2724 23.783
R40277 vdd.n2865 vdd.n2730 23.783
R40278 vdd.n2866 vdd.n2716 23.783
R40279 vdd.n2866 vdd.n2722 23.783
R40280 vdd.n2867 vdd.n2708 23.783
R40281 vdd.n2867 vdd.n2714 23.783
R40282 vdd.n2868 vdd.n2700 23.783
R40283 vdd.n2868 vdd.n2706 23.783
R40284 vdd.n2879 vdd.n2878 23.783
R40285 vdd.n2879 vdd.n2873 23.783
R40286 vdd.n3030 vdd.n3029 23.783
R40287 vdd.n3030 vdd.n3027 23.783
R40288 vdd.n3031 vdd.n3016 23.783
R40289 vdd.n3031 vdd.n3022 23.783
R40290 vdd.n3032 vdd.n3008 23.783
R40291 vdd.n3032 vdd.n3014 23.783
R40292 vdd.n3033 vdd.n3000 23.783
R40293 vdd.n3033 vdd.n3006 23.783
R40294 vdd.n3034 vdd.n2992 23.783
R40295 vdd.n3034 vdd.n2998 23.783
R40296 vdd.n3035 vdd.n2984 23.783
R40297 vdd.n3035 vdd.n2990 23.783
R40298 vdd.n3036 vdd.n2976 23.783
R40299 vdd.n3036 vdd.n2982 23.783
R40300 vdd.n3037 vdd.n2968 23.783
R40301 vdd.n3037 vdd.n2974 23.783
R40302 vdd.n3038 vdd.n2960 23.783
R40303 vdd.n3038 vdd.n2966 23.783
R40304 vdd.n3039 vdd.n2952 23.783
R40305 vdd.n3039 vdd.n2958 23.783
R40306 vdd.n3040 vdd.n2944 23.783
R40307 vdd.n3040 vdd.n2948 23.783
R40308 vdd.n3041 vdd.n2936 23.783
R40309 vdd.n3041 vdd.n2942 23.783
R40310 vdd.n3042 vdd.n2928 23.783
R40311 vdd.n3042 vdd.n2934 23.783
R40312 vdd.n3043 vdd.n2920 23.783
R40313 vdd.n3043 vdd.n2926 23.783
R40314 vdd.n3044 vdd.n2912 23.783
R40315 vdd.n3044 vdd.n2918 23.783
R40316 vdd.n3045 vdd.n2904 23.783
R40317 vdd.n3045 vdd.n2910 23.783
R40318 vdd.n3046 vdd.n2896 23.783
R40319 vdd.n3046 vdd.n2902 23.783
R40320 vdd.n3047 vdd.n2888 23.783
R40321 vdd.n3047 vdd.n2894 23.783
R40322 vdd.n3048 vdd.n2880 23.783
R40323 vdd.n3048 vdd.n2886 23.783
R40324 vdd.n3059 vdd.n3058 23.783
R40325 vdd.n3059 vdd.n3053 23.783
R40326 vdd.n3210 vdd.n3209 23.783
R40327 vdd.n3210 vdd.n3207 23.783
R40328 vdd.n3211 vdd.n3196 23.783
R40329 vdd.n3211 vdd.n3202 23.783
R40330 vdd.n3212 vdd.n3188 23.783
R40331 vdd.n3212 vdd.n3194 23.783
R40332 vdd.n3213 vdd.n3180 23.783
R40333 vdd.n3213 vdd.n3186 23.783
R40334 vdd.n3214 vdd.n3172 23.783
R40335 vdd.n3214 vdd.n3178 23.783
R40336 vdd.n3215 vdd.n3164 23.783
R40337 vdd.n3215 vdd.n3170 23.783
R40338 vdd.n3216 vdd.n3156 23.783
R40339 vdd.n3216 vdd.n3162 23.783
R40340 vdd.n3217 vdd.n3148 23.783
R40341 vdd.n3217 vdd.n3154 23.783
R40342 vdd.n3218 vdd.n3140 23.783
R40343 vdd.n3218 vdd.n3146 23.783
R40344 vdd.n3219 vdd.n3132 23.783
R40345 vdd.n3219 vdd.n3138 23.783
R40346 vdd.n3220 vdd.n3124 23.783
R40347 vdd.n3220 vdd.n3128 23.783
R40348 vdd.n3221 vdd.n3116 23.783
R40349 vdd.n3221 vdd.n3122 23.783
R40350 vdd.n3222 vdd.n3108 23.783
R40351 vdd.n3222 vdd.n3114 23.783
R40352 vdd.n3223 vdd.n3100 23.783
R40353 vdd.n3223 vdd.n3106 23.783
R40354 vdd.n3224 vdd.n3092 23.783
R40355 vdd.n3224 vdd.n3098 23.783
R40356 vdd.n3225 vdd.n3084 23.783
R40357 vdd.n3225 vdd.n3090 23.783
R40358 vdd.n3226 vdd.n3076 23.783
R40359 vdd.n3226 vdd.n3082 23.783
R40360 vdd.n3227 vdd.n3068 23.783
R40361 vdd.n3227 vdd.n3074 23.783
R40362 vdd.n3228 vdd.n3060 23.783
R40363 vdd.n3228 vdd.n3066 23.783
R40364 vdd.n3239 vdd.n3238 23.783
R40365 vdd.n3239 vdd.n3233 23.783
R40366 vdd.n3390 vdd.n3389 23.783
R40367 vdd.n3390 vdd.n3387 23.783
R40368 vdd.n3391 vdd.n3376 23.783
R40369 vdd.n3391 vdd.n3382 23.783
R40370 vdd.n3392 vdd.n3368 23.783
R40371 vdd.n3392 vdd.n3374 23.783
R40372 vdd.n3393 vdd.n3360 23.783
R40373 vdd.n3393 vdd.n3366 23.783
R40374 vdd.n3394 vdd.n3352 23.783
R40375 vdd.n3394 vdd.n3358 23.783
R40376 vdd.n3395 vdd.n3344 23.783
R40377 vdd.n3395 vdd.n3350 23.783
R40378 vdd.n3396 vdd.n3336 23.783
R40379 vdd.n3396 vdd.n3342 23.783
R40380 vdd.n3397 vdd.n3328 23.783
R40381 vdd.n3397 vdd.n3334 23.783
R40382 vdd.n3398 vdd.n3320 23.783
R40383 vdd.n3398 vdd.n3326 23.783
R40384 vdd.n3399 vdd.n3312 23.783
R40385 vdd.n3399 vdd.n3318 23.783
R40386 vdd.n3400 vdd.n3304 23.783
R40387 vdd.n3400 vdd.n3308 23.783
R40388 vdd.n3401 vdd.n3296 23.783
R40389 vdd.n3401 vdd.n3302 23.783
R40390 vdd.n3402 vdd.n3288 23.783
R40391 vdd.n3402 vdd.n3294 23.783
R40392 vdd.n3403 vdd.n3280 23.783
R40393 vdd.n3403 vdd.n3286 23.783
R40394 vdd.n3404 vdd.n3272 23.783
R40395 vdd.n3404 vdd.n3278 23.783
R40396 vdd.n3405 vdd.n3264 23.783
R40397 vdd.n3405 vdd.n3270 23.783
R40398 vdd.n3406 vdd.n3256 23.783
R40399 vdd.n3406 vdd.n3262 23.783
R40400 vdd.n3407 vdd.n3248 23.783
R40401 vdd.n3407 vdd.n3254 23.783
R40402 vdd.n3408 vdd.n3240 23.783
R40403 vdd.n3408 vdd.n3246 23.783
R40404 vdd.n3419 vdd.n3418 23.783
R40405 vdd.n3419 vdd.n3413 23.783
R40406 vdd.n3570 vdd.n3569 23.783
R40407 vdd.n3570 vdd.n3567 23.783
R40408 vdd.n3571 vdd.n3556 23.783
R40409 vdd.n3571 vdd.n3562 23.783
R40410 vdd.n3572 vdd.n3548 23.783
R40411 vdd.n3572 vdd.n3554 23.783
R40412 vdd.n3573 vdd.n3540 23.783
R40413 vdd.n3573 vdd.n3546 23.783
R40414 vdd.n3574 vdd.n3532 23.783
R40415 vdd.n3574 vdd.n3538 23.783
R40416 vdd.n3575 vdd.n3524 23.783
R40417 vdd.n3575 vdd.n3530 23.783
R40418 vdd.n3576 vdd.n3516 23.783
R40419 vdd.n3576 vdd.n3522 23.783
R40420 vdd.n3577 vdd.n3508 23.783
R40421 vdd.n3577 vdd.n3514 23.783
R40422 vdd.n3578 vdd.n3500 23.783
R40423 vdd.n3578 vdd.n3506 23.783
R40424 vdd.n3579 vdd.n3492 23.783
R40425 vdd.n3579 vdd.n3498 23.783
R40426 vdd.n3580 vdd.n3484 23.783
R40427 vdd.n3580 vdd.n3488 23.783
R40428 vdd.n3581 vdd.n3476 23.783
R40429 vdd.n3581 vdd.n3482 23.783
R40430 vdd.n3582 vdd.n3468 23.783
R40431 vdd.n3582 vdd.n3474 23.783
R40432 vdd.n3583 vdd.n3460 23.783
R40433 vdd.n3583 vdd.n3466 23.783
R40434 vdd.n3584 vdd.n3452 23.783
R40435 vdd.n3584 vdd.n3458 23.783
R40436 vdd.n3585 vdd.n3444 23.783
R40437 vdd.n3585 vdd.n3450 23.783
R40438 vdd.n3586 vdd.n3436 23.783
R40439 vdd.n3586 vdd.n3442 23.783
R40440 vdd.n3587 vdd.n3428 23.783
R40441 vdd.n3587 vdd.n3434 23.783
R40442 vdd.n3588 vdd.n3420 23.783
R40443 vdd.n3588 vdd.n3426 23.783
R40444 vdd.n3599 vdd.n3598 23.783
R40445 vdd.n3599 vdd.n3593 23.783
R40446 vdd.n3750 vdd.n3749 23.783
R40447 vdd.n3750 vdd.n3747 23.783
R40448 vdd.n3751 vdd.n3736 23.783
R40449 vdd.n3751 vdd.n3742 23.783
R40450 vdd.n3752 vdd.n3728 23.783
R40451 vdd.n3752 vdd.n3734 23.783
R40452 vdd.n3753 vdd.n3720 23.783
R40453 vdd.n3753 vdd.n3726 23.783
R40454 vdd.n3754 vdd.n3712 23.783
R40455 vdd.n3754 vdd.n3718 23.783
R40456 vdd.n3755 vdd.n3704 23.783
R40457 vdd.n3755 vdd.n3710 23.783
R40458 vdd.n3756 vdd.n3696 23.783
R40459 vdd.n3756 vdd.n3702 23.783
R40460 vdd.n3757 vdd.n3688 23.783
R40461 vdd.n3757 vdd.n3694 23.783
R40462 vdd.n3758 vdd.n3680 23.783
R40463 vdd.n3758 vdd.n3686 23.783
R40464 vdd.n3759 vdd.n3672 23.783
R40465 vdd.n3759 vdd.n3678 23.783
R40466 vdd.n3760 vdd.n3664 23.783
R40467 vdd.n3760 vdd.n3668 23.783
R40468 vdd.n3761 vdd.n3656 23.783
R40469 vdd.n3761 vdd.n3662 23.783
R40470 vdd.n3762 vdd.n3648 23.783
R40471 vdd.n3762 vdd.n3654 23.783
R40472 vdd.n3763 vdd.n3640 23.783
R40473 vdd.n3763 vdd.n3646 23.783
R40474 vdd.n3764 vdd.n3632 23.783
R40475 vdd.n3764 vdd.n3638 23.783
R40476 vdd.n3765 vdd.n3624 23.783
R40477 vdd.n3765 vdd.n3630 23.783
R40478 vdd.n3766 vdd.n3616 23.783
R40479 vdd.n3766 vdd.n3622 23.783
R40480 vdd.n3767 vdd.n3608 23.783
R40481 vdd.n3767 vdd.n3614 23.783
R40482 vdd.n3768 vdd.n3600 23.783
R40483 vdd.n3768 vdd.n3606 23.783
R40484 vdd.n3779 vdd.n3778 23.783
R40485 vdd.n3779 vdd.n3773 23.783
R40486 vdd.n3930 vdd.n3929 23.783
R40487 vdd.n3930 vdd.n3927 23.783
R40488 vdd.n3931 vdd.n3916 23.783
R40489 vdd.n3931 vdd.n3922 23.783
R40490 vdd.n3932 vdd.n3908 23.783
R40491 vdd.n3932 vdd.n3914 23.783
R40492 vdd.n3933 vdd.n3900 23.783
R40493 vdd.n3933 vdd.n3906 23.783
R40494 vdd.n3934 vdd.n3892 23.783
R40495 vdd.n3934 vdd.n3898 23.783
R40496 vdd.n3935 vdd.n3884 23.783
R40497 vdd.n3935 vdd.n3890 23.783
R40498 vdd.n3936 vdd.n3876 23.783
R40499 vdd.n3936 vdd.n3882 23.783
R40500 vdd.n3937 vdd.n3868 23.783
R40501 vdd.n3937 vdd.n3874 23.783
R40502 vdd.n3938 vdd.n3860 23.783
R40503 vdd.n3938 vdd.n3866 23.783
R40504 vdd.n3939 vdd.n3852 23.783
R40505 vdd.n3939 vdd.n3858 23.783
R40506 vdd.n3940 vdd.n3844 23.783
R40507 vdd.n3940 vdd.n3848 23.783
R40508 vdd.n3941 vdd.n3836 23.783
R40509 vdd.n3941 vdd.n3842 23.783
R40510 vdd.n3942 vdd.n3828 23.783
R40511 vdd.n3942 vdd.n3834 23.783
R40512 vdd.n3943 vdd.n3820 23.783
R40513 vdd.n3943 vdd.n3826 23.783
R40514 vdd.n3944 vdd.n3812 23.783
R40515 vdd.n3944 vdd.n3818 23.783
R40516 vdd.n3945 vdd.n3804 23.783
R40517 vdd.n3945 vdd.n3810 23.783
R40518 vdd.n3946 vdd.n3796 23.783
R40519 vdd.n3946 vdd.n3802 23.783
R40520 vdd.n3947 vdd.n3788 23.783
R40521 vdd.n3947 vdd.n3794 23.783
R40522 vdd.n3948 vdd.n3780 23.783
R40523 vdd.n3948 vdd.n3786 23.783
R40524 vdd.n3959 vdd.n3958 23.783
R40525 vdd.n3959 vdd.n3953 23.783
R40526 vdd.n4110 vdd.n4109 23.783
R40527 vdd.n4110 vdd.n4107 23.783
R40528 vdd.n4111 vdd.n4096 23.783
R40529 vdd.n4111 vdd.n4102 23.783
R40530 vdd.n4112 vdd.n4088 23.783
R40531 vdd.n4112 vdd.n4094 23.783
R40532 vdd.n4113 vdd.n4080 23.783
R40533 vdd.n4113 vdd.n4086 23.783
R40534 vdd.n4114 vdd.n4072 23.783
R40535 vdd.n4114 vdd.n4078 23.783
R40536 vdd.n4115 vdd.n4064 23.783
R40537 vdd.n4115 vdd.n4070 23.783
R40538 vdd.n4116 vdd.n4056 23.783
R40539 vdd.n4116 vdd.n4062 23.783
R40540 vdd.n4117 vdd.n4048 23.783
R40541 vdd.n4117 vdd.n4054 23.783
R40542 vdd.n4118 vdd.n4040 23.783
R40543 vdd.n4118 vdd.n4046 23.783
R40544 vdd.n4119 vdd.n4032 23.783
R40545 vdd.n4119 vdd.n4038 23.783
R40546 vdd.n4120 vdd.n4024 23.783
R40547 vdd.n4120 vdd.n4028 23.783
R40548 vdd.n4121 vdd.n4016 23.783
R40549 vdd.n4121 vdd.n4022 23.783
R40550 vdd.n4122 vdd.n4008 23.783
R40551 vdd.n4122 vdd.n4014 23.783
R40552 vdd.n4123 vdd.n4000 23.783
R40553 vdd.n4123 vdd.n4006 23.783
R40554 vdd.n4124 vdd.n3992 23.783
R40555 vdd.n4124 vdd.n3998 23.783
R40556 vdd.n4125 vdd.n3984 23.783
R40557 vdd.n4125 vdd.n3990 23.783
R40558 vdd.n4126 vdd.n3976 23.783
R40559 vdd.n4126 vdd.n3982 23.783
R40560 vdd.n4127 vdd.n3968 23.783
R40561 vdd.n4127 vdd.n3974 23.783
R40562 vdd.n4128 vdd.n3960 23.783
R40563 vdd.n4128 vdd.n3966 23.783
R40564 vdd.n4139 vdd.n4138 23.783
R40565 vdd.n4139 vdd.n4133 23.783
R40566 vdd.n4290 vdd.n4289 23.783
R40567 vdd.n4290 vdd.n4287 23.783
R40568 vdd.n4291 vdd.n4276 23.783
R40569 vdd.n4291 vdd.n4282 23.783
R40570 vdd.n4292 vdd.n4268 23.783
R40571 vdd.n4292 vdd.n4274 23.783
R40572 vdd.n4293 vdd.n4260 23.783
R40573 vdd.n4293 vdd.n4266 23.783
R40574 vdd.n4294 vdd.n4252 23.783
R40575 vdd.n4294 vdd.n4258 23.783
R40576 vdd.n4295 vdd.n4244 23.783
R40577 vdd.n4295 vdd.n4250 23.783
R40578 vdd.n4296 vdd.n4236 23.783
R40579 vdd.n4296 vdd.n4242 23.783
R40580 vdd.n4297 vdd.n4228 23.783
R40581 vdd.n4297 vdd.n4234 23.783
R40582 vdd.n4298 vdd.n4220 23.783
R40583 vdd.n4298 vdd.n4226 23.783
R40584 vdd.n4299 vdd.n4212 23.783
R40585 vdd.n4299 vdd.n4218 23.783
R40586 vdd.n4300 vdd.n4204 23.783
R40587 vdd.n4300 vdd.n4208 23.783
R40588 vdd.n4301 vdd.n4196 23.783
R40589 vdd.n4301 vdd.n4202 23.783
R40590 vdd.n4302 vdd.n4188 23.783
R40591 vdd.n4302 vdd.n4194 23.783
R40592 vdd.n4303 vdd.n4180 23.783
R40593 vdd.n4303 vdd.n4186 23.783
R40594 vdd.n4304 vdd.n4172 23.783
R40595 vdd.n4304 vdd.n4178 23.783
R40596 vdd.n4305 vdd.n4164 23.783
R40597 vdd.n4305 vdd.n4170 23.783
R40598 vdd.n4306 vdd.n4156 23.783
R40599 vdd.n4306 vdd.n4162 23.783
R40600 vdd.n4307 vdd.n4148 23.783
R40601 vdd.n4307 vdd.n4154 23.783
R40602 vdd.n4308 vdd.n4140 23.783
R40603 vdd.n4308 vdd.n4146 23.783
R40604 vdd.n4319 vdd.n4318 23.783
R40605 vdd.n4319 vdd.n4313 23.783
R40606 vdd.n4470 vdd.n4469 23.783
R40607 vdd.n4470 vdd.n4467 23.783
R40608 vdd.n4471 vdd.n4456 23.783
R40609 vdd.n4471 vdd.n4462 23.783
R40610 vdd.n4472 vdd.n4448 23.783
R40611 vdd.n4472 vdd.n4454 23.783
R40612 vdd.n4473 vdd.n4440 23.783
R40613 vdd.n4473 vdd.n4446 23.783
R40614 vdd.n4474 vdd.n4432 23.783
R40615 vdd.n4474 vdd.n4438 23.783
R40616 vdd.n4475 vdd.n4424 23.783
R40617 vdd.n4475 vdd.n4430 23.783
R40618 vdd.n4476 vdd.n4416 23.783
R40619 vdd.n4476 vdd.n4422 23.783
R40620 vdd.n4477 vdd.n4408 23.783
R40621 vdd.n4477 vdd.n4414 23.783
R40622 vdd.n4478 vdd.n4400 23.783
R40623 vdd.n4478 vdd.n4406 23.783
R40624 vdd.n4479 vdd.n4392 23.783
R40625 vdd.n4479 vdd.n4398 23.783
R40626 vdd.n4480 vdd.n4384 23.783
R40627 vdd.n4480 vdd.n4388 23.783
R40628 vdd.n4481 vdd.n4376 23.783
R40629 vdd.n4481 vdd.n4382 23.783
R40630 vdd.n4482 vdd.n4368 23.783
R40631 vdd.n4482 vdd.n4374 23.783
R40632 vdd.n4483 vdd.n4360 23.783
R40633 vdd.n4483 vdd.n4366 23.783
R40634 vdd.n4484 vdd.n4352 23.783
R40635 vdd.n4484 vdd.n4358 23.783
R40636 vdd.n4485 vdd.n4344 23.783
R40637 vdd.n4485 vdd.n4350 23.783
R40638 vdd.n4486 vdd.n4336 23.783
R40639 vdd.n4486 vdd.n4342 23.783
R40640 vdd.n4487 vdd.n4328 23.783
R40641 vdd.n4487 vdd.n4334 23.783
R40642 vdd.n4488 vdd.n4320 23.783
R40643 vdd.n4488 vdd.n4326 23.783
R40644 vdd.n4499 vdd.n4498 23.783
R40645 vdd.n4499 vdd.n4493 23.783
R40646 vdd.n4650 vdd.n4649 23.783
R40647 vdd.n4650 vdd.n4647 23.783
R40648 vdd.n4651 vdd.n4636 23.783
R40649 vdd.n4651 vdd.n4642 23.783
R40650 vdd.n4652 vdd.n4628 23.783
R40651 vdd.n4652 vdd.n4634 23.783
R40652 vdd.n4653 vdd.n4620 23.783
R40653 vdd.n4653 vdd.n4626 23.783
R40654 vdd.n4654 vdd.n4612 23.783
R40655 vdd.n4654 vdd.n4618 23.783
R40656 vdd.n4655 vdd.n4604 23.783
R40657 vdd.n4655 vdd.n4610 23.783
R40658 vdd.n4656 vdd.n4596 23.783
R40659 vdd.n4656 vdd.n4602 23.783
R40660 vdd.n4657 vdd.n4588 23.783
R40661 vdd.n4657 vdd.n4594 23.783
R40662 vdd.n4658 vdd.n4580 23.783
R40663 vdd.n4658 vdd.n4586 23.783
R40664 vdd.n4659 vdd.n4572 23.783
R40665 vdd.n4659 vdd.n4578 23.783
R40666 vdd.n4660 vdd.n4564 23.783
R40667 vdd.n4660 vdd.n4568 23.783
R40668 vdd.n4661 vdd.n4556 23.783
R40669 vdd.n4661 vdd.n4562 23.783
R40670 vdd.n4662 vdd.n4548 23.783
R40671 vdd.n4662 vdd.n4554 23.783
R40672 vdd.n4663 vdd.n4540 23.783
R40673 vdd.n4663 vdd.n4546 23.783
R40674 vdd.n4664 vdd.n4532 23.783
R40675 vdd.n4664 vdd.n4538 23.783
R40676 vdd.n4665 vdd.n4524 23.783
R40677 vdd.n4665 vdd.n4530 23.783
R40678 vdd.n4666 vdd.n4516 23.783
R40679 vdd.n4666 vdd.n4522 23.783
R40680 vdd.n4667 vdd.n4508 23.783
R40681 vdd.n4667 vdd.n4514 23.783
R40682 vdd.n4668 vdd.n4500 23.783
R40683 vdd.n4668 vdd.n4506 23.783
R40684 vdd.n4679 vdd.n4678 23.783
R40685 vdd.n4679 vdd.n4673 23.783
R40686 vdd.n4830 vdd.n4829 23.783
R40687 vdd.n4830 vdd.n4827 23.783
R40688 vdd.n4831 vdd.n4816 23.783
R40689 vdd.n4831 vdd.n4822 23.783
R40690 vdd.n4832 vdd.n4808 23.783
R40691 vdd.n4832 vdd.n4814 23.783
R40692 vdd.n4833 vdd.n4800 23.783
R40693 vdd.n4833 vdd.n4806 23.783
R40694 vdd.n4834 vdd.n4792 23.783
R40695 vdd.n4834 vdd.n4798 23.783
R40696 vdd.n4835 vdd.n4784 23.783
R40697 vdd.n4835 vdd.n4790 23.783
R40698 vdd.n4836 vdd.n4776 23.783
R40699 vdd.n4836 vdd.n4782 23.783
R40700 vdd.n4837 vdd.n4768 23.783
R40701 vdd.n4837 vdd.n4774 23.783
R40702 vdd.n4838 vdd.n4760 23.783
R40703 vdd.n4838 vdd.n4766 23.783
R40704 vdd.n4839 vdd.n4752 23.783
R40705 vdd.n4839 vdd.n4758 23.783
R40706 vdd.n4840 vdd.n4744 23.783
R40707 vdd.n4840 vdd.n4748 23.783
R40708 vdd.n4841 vdd.n4736 23.783
R40709 vdd.n4841 vdd.n4742 23.783
R40710 vdd.n4842 vdd.n4728 23.783
R40711 vdd.n4842 vdd.n4734 23.783
R40712 vdd.n4843 vdd.n4720 23.783
R40713 vdd.n4843 vdd.n4726 23.783
R40714 vdd.n4844 vdd.n4712 23.783
R40715 vdd.n4844 vdd.n4718 23.783
R40716 vdd.n4845 vdd.n4704 23.783
R40717 vdd.n4845 vdd.n4710 23.783
R40718 vdd.n4846 vdd.n4696 23.783
R40719 vdd.n4846 vdd.n4702 23.783
R40720 vdd.n4847 vdd.n4688 23.783
R40721 vdd.n4847 vdd.n4694 23.783
R40722 vdd.n4848 vdd.n4680 23.783
R40723 vdd.n4848 vdd.n4686 23.783
R40724 vdd.n4859 vdd.n4858 23.783
R40725 vdd.n4859 vdd.n4853 23.783
R40726 vdd.n5010 vdd.n5009 23.783
R40727 vdd.n5010 vdd.n5007 23.783
R40728 vdd.n5011 vdd.n4996 23.783
R40729 vdd.n5011 vdd.n5002 23.783
R40730 vdd.n5012 vdd.n4988 23.783
R40731 vdd.n5012 vdd.n4994 23.783
R40732 vdd.n5013 vdd.n4980 23.783
R40733 vdd.n5013 vdd.n4986 23.783
R40734 vdd.n5014 vdd.n4972 23.783
R40735 vdd.n5014 vdd.n4978 23.783
R40736 vdd.n5015 vdd.n4964 23.783
R40737 vdd.n5015 vdd.n4970 23.783
R40738 vdd.n5016 vdd.n4956 23.783
R40739 vdd.n5016 vdd.n4962 23.783
R40740 vdd.n5017 vdd.n4948 23.783
R40741 vdd.n5017 vdd.n4954 23.783
R40742 vdd.n5018 vdd.n4940 23.783
R40743 vdd.n5018 vdd.n4946 23.783
R40744 vdd.n5019 vdd.n4932 23.783
R40745 vdd.n5019 vdd.n4938 23.783
R40746 vdd.n5020 vdd.n4924 23.783
R40747 vdd.n5020 vdd.n4928 23.783
R40748 vdd.n5021 vdd.n4916 23.783
R40749 vdd.n5021 vdd.n4922 23.783
R40750 vdd.n5022 vdd.n4908 23.783
R40751 vdd.n5022 vdd.n4914 23.783
R40752 vdd.n5023 vdd.n4900 23.783
R40753 vdd.n5023 vdd.n4906 23.783
R40754 vdd.n5024 vdd.n4892 23.783
R40755 vdd.n5024 vdd.n4898 23.783
R40756 vdd.n5025 vdd.n4884 23.783
R40757 vdd.n5025 vdd.n4890 23.783
R40758 vdd.n5026 vdd.n4876 23.783
R40759 vdd.n5026 vdd.n4882 23.783
R40760 vdd.n5027 vdd.n4868 23.783
R40761 vdd.n5027 vdd.n4874 23.783
R40762 vdd.n5028 vdd.n4860 23.783
R40763 vdd.n5028 vdd.n4866 23.783
R40764 vdd.n5039 vdd.n5038 23.783
R40765 vdd.n5039 vdd.n5033 23.783
R40766 vdd.n5190 vdd.n5189 23.783
R40767 vdd.n5190 vdd.n5187 23.783
R40768 vdd.n5191 vdd.n5176 23.783
R40769 vdd.n5191 vdd.n5182 23.783
R40770 vdd.n5192 vdd.n5168 23.783
R40771 vdd.n5192 vdd.n5174 23.783
R40772 vdd.n5193 vdd.n5160 23.783
R40773 vdd.n5193 vdd.n5166 23.783
R40774 vdd.n5194 vdd.n5152 23.783
R40775 vdd.n5194 vdd.n5158 23.783
R40776 vdd.n5195 vdd.n5144 23.783
R40777 vdd.n5195 vdd.n5150 23.783
R40778 vdd.n5196 vdd.n5136 23.783
R40779 vdd.n5196 vdd.n5142 23.783
R40780 vdd.n5197 vdd.n5128 23.783
R40781 vdd.n5197 vdd.n5134 23.783
R40782 vdd.n5198 vdd.n5120 23.783
R40783 vdd.n5198 vdd.n5126 23.783
R40784 vdd.n5199 vdd.n5112 23.783
R40785 vdd.n5199 vdd.n5118 23.783
R40786 vdd.n5200 vdd.n5104 23.783
R40787 vdd.n5200 vdd.n5108 23.783
R40788 vdd.n5201 vdd.n5096 23.783
R40789 vdd.n5201 vdd.n5102 23.783
R40790 vdd.n5202 vdd.n5088 23.783
R40791 vdd.n5202 vdd.n5094 23.783
R40792 vdd.n5203 vdd.n5080 23.783
R40793 vdd.n5203 vdd.n5086 23.783
R40794 vdd.n5204 vdd.n5072 23.783
R40795 vdd.n5204 vdd.n5078 23.783
R40796 vdd.n5205 vdd.n5064 23.783
R40797 vdd.n5205 vdd.n5070 23.783
R40798 vdd.n5206 vdd.n5056 23.783
R40799 vdd.n5206 vdd.n5062 23.783
R40800 vdd.n5207 vdd.n5048 23.783
R40801 vdd.n5207 vdd.n5054 23.783
R40802 vdd.n5208 vdd.n5040 23.783
R40803 vdd.n5208 vdd.n5046 23.783
R40804 vdd.n5219 vdd.n5218 23.783
R40805 vdd.n5219 vdd.n5213 23.783
R40806 vdd.n5370 vdd.n5369 23.783
R40807 vdd.n5370 vdd.n5367 23.783
R40808 vdd.n5371 vdd.n5356 23.783
R40809 vdd.n5371 vdd.n5362 23.783
R40810 vdd.n5372 vdd.n5348 23.783
R40811 vdd.n5372 vdd.n5354 23.783
R40812 vdd.n5373 vdd.n5340 23.783
R40813 vdd.n5373 vdd.n5346 23.783
R40814 vdd.n5374 vdd.n5332 23.783
R40815 vdd.n5374 vdd.n5338 23.783
R40816 vdd.n5375 vdd.n5324 23.783
R40817 vdd.n5375 vdd.n5330 23.783
R40818 vdd.n5376 vdd.n5316 23.783
R40819 vdd.n5376 vdd.n5322 23.783
R40820 vdd.n5377 vdd.n5308 23.783
R40821 vdd.n5377 vdd.n5314 23.783
R40822 vdd.n5378 vdd.n5300 23.783
R40823 vdd.n5378 vdd.n5306 23.783
R40824 vdd.n5379 vdd.n5292 23.783
R40825 vdd.n5379 vdd.n5298 23.783
R40826 vdd.n5380 vdd.n5284 23.783
R40827 vdd.n5380 vdd.n5288 23.783
R40828 vdd.n5381 vdd.n5276 23.783
R40829 vdd.n5381 vdd.n5282 23.783
R40830 vdd.n5382 vdd.n5268 23.783
R40831 vdd.n5382 vdd.n5274 23.783
R40832 vdd.n5383 vdd.n5260 23.783
R40833 vdd.n5383 vdd.n5266 23.783
R40834 vdd.n5384 vdd.n5252 23.783
R40835 vdd.n5384 vdd.n5258 23.783
R40836 vdd.n5385 vdd.n5244 23.783
R40837 vdd.n5385 vdd.n5250 23.783
R40838 vdd.n5386 vdd.n5236 23.783
R40839 vdd.n5386 vdd.n5242 23.783
R40840 vdd.n5387 vdd.n5228 23.783
R40841 vdd.n5387 vdd.n5234 23.783
R40842 vdd.n5388 vdd.n5220 23.783
R40843 vdd.n5388 vdd.n5226 23.783
R40844 vdd.n5399 vdd.n5398 23.783
R40845 vdd.n5399 vdd.n5393 23.783
R40846 vdd.n5550 vdd.n5549 23.783
R40847 vdd.n5550 vdd.n5547 23.783
R40848 vdd.n5551 vdd.n5536 23.783
R40849 vdd.n5551 vdd.n5542 23.783
R40850 vdd.n5552 vdd.n5528 23.783
R40851 vdd.n5552 vdd.n5534 23.783
R40852 vdd.n5553 vdd.n5520 23.783
R40853 vdd.n5553 vdd.n5526 23.783
R40854 vdd.n5554 vdd.n5512 23.783
R40855 vdd.n5554 vdd.n5518 23.783
R40856 vdd.n5555 vdd.n5504 23.783
R40857 vdd.n5555 vdd.n5510 23.783
R40858 vdd.n5556 vdd.n5496 23.783
R40859 vdd.n5556 vdd.n5502 23.783
R40860 vdd.n5557 vdd.n5488 23.783
R40861 vdd.n5557 vdd.n5494 23.783
R40862 vdd.n5558 vdd.n5480 23.783
R40863 vdd.n5558 vdd.n5486 23.783
R40864 vdd.n5559 vdd.n5472 23.783
R40865 vdd.n5559 vdd.n5478 23.783
R40866 vdd.n5560 vdd.n5464 23.783
R40867 vdd.n5560 vdd.n5468 23.783
R40868 vdd.n5561 vdd.n5456 23.783
R40869 vdd.n5561 vdd.n5462 23.783
R40870 vdd.n5562 vdd.n5448 23.783
R40871 vdd.n5562 vdd.n5454 23.783
R40872 vdd.n5563 vdd.n5440 23.783
R40873 vdd.n5563 vdd.n5446 23.783
R40874 vdd.n5564 vdd.n5432 23.783
R40875 vdd.n5564 vdd.n5438 23.783
R40876 vdd.n5565 vdd.n5424 23.783
R40877 vdd.n5565 vdd.n5430 23.783
R40878 vdd.n5566 vdd.n5416 23.783
R40879 vdd.n5566 vdd.n5422 23.783
R40880 vdd.n5567 vdd.n5408 23.783
R40881 vdd.n5567 vdd.n5414 23.783
R40882 vdd.n5568 vdd.n5400 23.783
R40883 vdd.n5568 vdd.n5406 23.783
R40884 vdd.n5579 vdd.n5578 23.783
R40885 vdd.n5579 vdd.n5573 23.783
R40886 vdd.n5730 vdd.n5729 23.783
R40887 vdd.n5730 vdd.n5727 23.783
R40888 vdd.n5731 vdd.n5716 23.783
R40889 vdd.n5731 vdd.n5722 23.783
R40890 vdd.n5732 vdd.n5708 23.783
R40891 vdd.n5732 vdd.n5714 23.783
R40892 vdd.n5733 vdd.n5700 23.783
R40893 vdd.n5733 vdd.n5706 23.783
R40894 vdd.n5734 vdd.n5692 23.783
R40895 vdd.n5734 vdd.n5698 23.783
R40896 vdd.n5735 vdd.n5684 23.783
R40897 vdd.n5735 vdd.n5690 23.783
R40898 vdd.n5736 vdd.n5676 23.783
R40899 vdd.n5736 vdd.n5682 23.783
R40900 vdd.n5737 vdd.n5668 23.783
R40901 vdd.n5737 vdd.n5674 23.783
R40902 vdd.n5738 vdd.n5660 23.783
R40903 vdd.n5738 vdd.n5666 23.783
R40904 vdd.n5739 vdd.n5652 23.783
R40905 vdd.n5739 vdd.n5658 23.783
R40906 vdd.n5740 vdd.n5644 23.783
R40907 vdd.n5740 vdd.n5648 23.783
R40908 vdd.n5741 vdd.n5636 23.783
R40909 vdd.n5741 vdd.n5642 23.783
R40910 vdd.n5742 vdd.n5628 23.783
R40911 vdd.n5742 vdd.n5634 23.783
R40912 vdd.n5743 vdd.n5620 23.783
R40913 vdd.n5743 vdd.n5626 23.783
R40914 vdd.n5744 vdd.n5612 23.783
R40915 vdd.n5744 vdd.n5618 23.783
R40916 vdd.n5745 vdd.n5604 23.783
R40917 vdd.n5745 vdd.n5610 23.783
R40918 vdd.n5746 vdd.n5596 23.783
R40919 vdd.n5746 vdd.n5602 23.783
R40920 vdd.n5747 vdd.n5588 23.783
R40921 vdd.n5747 vdd.n5594 23.783
R40922 vdd.n5748 vdd.n5580 23.783
R40923 vdd.n5748 vdd.n5586 23.783
R40924 vdd.n5759 vdd.n5758 23.783
R40925 vdd.n5759 vdd.n5753 23.783
R40926 vdd.n5910 vdd.n5909 23.783
R40927 vdd.n5910 vdd.n5907 23.783
R40928 vdd.n5911 vdd.n5896 23.783
R40929 vdd.n5911 vdd.n5902 23.783
R40930 vdd.n5912 vdd.n5888 23.783
R40931 vdd.n5912 vdd.n5894 23.783
R40932 vdd.n5913 vdd.n5880 23.783
R40933 vdd.n5913 vdd.n5886 23.783
R40934 vdd.n5914 vdd.n5872 23.783
R40935 vdd.n5914 vdd.n5878 23.783
R40936 vdd.n5915 vdd.n5864 23.783
R40937 vdd.n5915 vdd.n5870 23.783
R40938 vdd.n5916 vdd.n5856 23.783
R40939 vdd.n5916 vdd.n5862 23.783
R40940 vdd.n5917 vdd.n5848 23.783
R40941 vdd.n5917 vdd.n5854 23.783
R40942 vdd.n5918 vdd.n5840 23.783
R40943 vdd.n5918 vdd.n5846 23.783
R40944 vdd.n5919 vdd.n5832 23.783
R40945 vdd.n5919 vdd.n5838 23.783
R40946 vdd.n5920 vdd.n5824 23.783
R40947 vdd.n5920 vdd.n5828 23.783
R40948 vdd.n5921 vdd.n5816 23.783
R40949 vdd.n5921 vdd.n5822 23.783
R40950 vdd.n5922 vdd.n5808 23.783
R40951 vdd.n5922 vdd.n5814 23.783
R40952 vdd.n5923 vdd.n5800 23.783
R40953 vdd.n5923 vdd.n5806 23.783
R40954 vdd.n5924 vdd.n5792 23.783
R40955 vdd.n5924 vdd.n5798 23.783
R40956 vdd.n5925 vdd.n5784 23.783
R40957 vdd.n5925 vdd.n5790 23.783
R40958 vdd.n5926 vdd.n5776 23.783
R40959 vdd.n5926 vdd.n5782 23.783
R40960 vdd.n5927 vdd.n5768 23.783
R40961 vdd.n5927 vdd.n5774 23.783
R40962 vdd.n5928 vdd.n5760 23.783
R40963 vdd.n5928 vdd.n5766 23.783
R40964 vdd.n5939 vdd.n5938 23.783
R40965 vdd.n5939 vdd.n5933 23.783
R40966 vdd.n6090 vdd.n6089 23.783
R40967 vdd.n6090 vdd.n6087 23.783
R40968 vdd.n6091 vdd.n6076 23.783
R40969 vdd.n6091 vdd.n6082 23.783
R40970 vdd.n6092 vdd.n6068 23.783
R40971 vdd.n6092 vdd.n6074 23.783
R40972 vdd.n6093 vdd.n6060 23.783
R40973 vdd.n6093 vdd.n6066 23.783
R40974 vdd.n6094 vdd.n6052 23.783
R40975 vdd.n6094 vdd.n6058 23.783
R40976 vdd.n6095 vdd.n6044 23.783
R40977 vdd.n6095 vdd.n6050 23.783
R40978 vdd.n6096 vdd.n6036 23.783
R40979 vdd.n6096 vdd.n6042 23.783
R40980 vdd.n6097 vdd.n6028 23.783
R40981 vdd.n6097 vdd.n6034 23.783
R40982 vdd.n6098 vdd.n6020 23.783
R40983 vdd.n6098 vdd.n6026 23.783
R40984 vdd.n6099 vdd.n6012 23.783
R40985 vdd.n6099 vdd.n6018 23.783
R40986 vdd.n6100 vdd.n6004 23.783
R40987 vdd.n6100 vdd.n6008 23.783
R40988 vdd.n6101 vdd.n5996 23.783
R40989 vdd.n6101 vdd.n6002 23.783
R40990 vdd.n6102 vdd.n5988 23.783
R40991 vdd.n6102 vdd.n5994 23.783
R40992 vdd.n6103 vdd.n5980 23.783
R40993 vdd.n6103 vdd.n5986 23.783
R40994 vdd.n6104 vdd.n5972 23.783
R40995 vdd.n6104 vdd.n5978 23.783
R40996 vdd.n6105 vdd.n5964 23.783
R40997 vdd.n6105 vdd.n5970 23.783
R40998 vdd.n6106 vdd.n5956 23.783
R40999 vdd.n6106 vdd.n5962 23.783
R41000 vdd.n6107 vdd.n5948 23.783
R41001 vdd.n6107 vdd.n5954 23.783
R41002 vdd.n6108 vdd.n5940 23.783
R41003 vdd.n6108 vdd.n5946 23.783
R41004 vdd.n6119 vdd.n6118 23.783
R41005 vdd.n6119 vdd.n6113 23.783
R41006 vdd.n6270 vdd.n6269 23.783
R41007 vdd.n6270 vdd.n6267 23.783
R41008 vdd.n6271 vdd.n6256 23.783
R41009 vdd.n6271 vdd.n6262 23.783
R41010 vdd.n6272 vdd.n6248 23.783
R41011 vdd.n6272 vdd.n6254 23.783
R41012 vdd.n6273 vdd.n6240 23.783
R41013 vdd.n6273 vdd.n6246 23.783
R41014 vdd.n6274 vdd.n6232 23.783
R41015 vdd.n6274 vdd.n6238 23.783
R41016 vdd.n6275 vdd.n6224 23.783
R41017 vdd.n6275 vdd.n6230 23.783
R41018 vdd.n6276 vdd.n6216 23.783
R41019 vdd.n6276 vdd.n6222 23.783
R41020 vdd.n6277 vdd.n6208 23.783
R41021 vdd.n6277 vdd.n6214 23.783
R41022 vdd.n6278 vdd.n6200 23.783
R41023 vdd.n6278 vdd.n6206 23.783
R41024 vdd.n6279 vdd.n6192 23.783
R41025 vdd.n6279 vdd.n6198 23.783
R41026 vdd.n6280 vdd.n6184 23.783
R41027 vdd.n6280 vdd.n6188 23.783
R41028 vdd.n6281 vdd.n6176 23.783
R41029 vdd.n6281 vdd.n6182 23.783
R41030 vdd.n6282 vdd.n6168 23.783
R41031 vdd.n6282 vdd.n6174 23.783
R41032 vdd.n6283 vdd.n6160 23.783
R41033 vdd.n6283 vdd.n6166 23.783
R41034 vdd.n6284 vdd.n6152 23.783
R41035 vdd.n6284 vdd.n6158 23.783
R41036 vdd.n6285 vdd.n6144 23.783
R41037 vdd.n6285 vdd.n6150 23.783
R41038 vdd.n6286 vdd.n6136 23.783
R41039 vdd.n6286 vdd.n6142 23.783
R41040 vdd.n6287 vdd.n6128 23.783
R41041 vdd.n6287 vdd.n6134 23.783
R41042 vdd.n6288 vdd.n6120 23.783
R41043 vdd.n6288 vdd.n6126 23.783
R41044 vdd.n6299 vdd.n6298 23.783
R41045 vdd.n6299 vdd.n6293 23.783
R41046 vdd.n6450 vdd.n6449 23.783
R41047 vdd.n6450 vdd.n6447 23.783
R41048 vdd.n6451 vdd.n6436 23.783
R41049 vdd.n6451 vdd.n6442 23.783
R41050 vdd.n6452 vdd.n6428 23.783
R41051 vdd.n6452 vdd.n6434 23.783
R41052 vdd.n6453 vdd.n6420 23.783
R41053 vdd.n6453 vdd.n6426 23.783
R41054 vdd.n6454 vdd.n6412 23.783
R41055 vdd.n6454 vdd.n6418 23.783
R41056 vdd.n6455 vdd.n6404 23.783
R41057 vdd.n6455 vdd.n6410 23.783
R41058 vdd.n6456 vdd.n6396 23.783
R41059 vdd.n6456 vdd.n6402 23.783
R41060 vdd.n6457 vdd.n6388 23.783
R41061 vdd.n6457 vdd.n6394 23.783
R41062 vdd.n6458 vdd.n6380 23.783
R41063 vdd.n6458 vdd.n6386 23.783
R41064 vdd.n6459 vdd.n6372 23.783
R41065 vdd.n6459 vdd.n6378 23.783
R41066 vdd.n6460 vdd.n6364 23.783
R41067 vdd.n6460 vdd.n6368 23.783
R41068 vdd.n6461 vdd.n6356 23.783
R41069 vdd.n6461 vdd.n6362 23.783
R41070 vdd.n6462 vdd.n6348 23.783
R41071 vdd.n6462 vdd.n6354 23.783
R41072 vdd.n6463 vdd.n6340 23.783
R41073 vdd.n6463 vdd.n6346 23.783
R41074 vdd.n6464 vdd.n6332 23.783
R41075 vdd.n6464 vdd.n6338 23.783
R41076 vdd.n6465 vdd.n6324 23.783
R41077 vdd.n6465 vdd.n6330 23.783
R41078 vdd.n6466 vdd.n6316 23.783
R41079 vdd.n6466 vdd.n6322 23.783
R41080 vdd.n6467 vdd.n6308 23.783
R41081 vdd.n6467 vdd.n6314 23.783
R41082 vdd.n6468 vdd.n6300 23.783
R41083 vdd.n6468 vdd.n6306 23.783
R41084 vdd.n6479 vdd.n6478 23.783
R41085 vdd.n6479 vdd.n6473 23.783
R41086 vdd.n6630 vdd.n6629 23.783
R41087 vdd.n6630 vdd.n6627 23.783
R41088 vdd.n6631 vdd.n6616 23.783
R41089 vdd.n6631 vdd.n6622 23.783
R41090 vdd.n6632 vdd.n6608 23.783
R41091 vdd.n6632 vdd.n6614 23.783
R41092 vdd.n6633 vdd.n6600 23.783
R41093 vdd.n6633 vdd.n6606 23.783
R41094 vdd.n6634 vdd.n6592 23.783
R41095 vdd.n6634 vdd.n6598 23.783
R41096 vdd.n6635 vdd.n6584 23.783
R41097 vdd.n6635 vdd.n6590 23.783
R41098 vdd.n6636 vdd.n6576 23.783
R41099 vdd.n6636 vdd.n6582 23.783
R41100 vdd.n6637 vdd.n6568 23.783
R41101 vdd.n6637 vdd.n6574 23.783
R41102 vdd.n6638 vdd.n6560 23.783
R41103 vdd.n6638 vdd.n6566 23.783
R41104 vdd.n6639 vdd.n6552 23.783
R41105 vdd.n6639 vdd.n6558 23.783
R41106 vdd.n6640 vdd.n6544 23.783
R41107 vdd.n6640 vdd.n6548 23.783
R41108 vdd.n6641 vdd.n6536 23.783
R41109 vdd.n6641 vdd.n6542 23.783
R41110 vdd.n6642 vdd.n6528 23.783
R41111 vdd.n6642 vdd.n6534 23.783
R41112 vdd.n6643 vdd.n6520 23.783
R41113 vdd.n6643 vdd.n6526 23.783
R41114 vdd.n6644 vdd.n6512 23.783
R41115 vdd.n6644 vdd.n6518 23.783
R41116 vdd.n6645 vdd.n6504 23.783
R41117 vdd.n6645 vdd.n6510 23.783
R41118 vdd.n6646 vdd.n6496 23.783
R41119 vdd.n6646 vdd.n6502 23.783
R41120 vdd.n6647 vdd.n6488 23.783
R41121 vdd.n6647 vdd.n6494 23.783
R41122 vdd.n6648 vdd.n6480 23.783
R41123 vdd.n6648 vdd.n6486 23.783
R41124 vdd.n6659 vdd.n6658 23.783
R41125 vdd.n6659 vdd.n6653 23.783
R41126 vdd.n6810 vdd.n6809 23.783
R41127 vdd.n6810 vdd.n6807 23.783
R41128 vdd.n6811 vdd.n6796 23.783
R41129 vdd.n6811 vdd.n6802 23.783
R41130 vdd.n6812 vdd.n6788 23.783
R41131 vdd.n6812 vdd.n6794 23.783
R41132 vdd.n6813 vdd.n6780 23.783
R41133 vdd.n6813 vdd.n6786 23.783
R41134 vdd.n6814 vdd.n6772 23.783
R41135 vdd.n6814 vdd.n6778 23.783
R41136 vdd.n6815 vdd.n6764 23.783
R41137 vdd.n6815 vdd.n6770 23.783
R41138 vdd.n6816 vdd.n6756 23.783
R41139 vdd.n6816 vdd.n6762 23.783
R41140 vdd.n6817 vdd.n6748 23.783
R41141 vdd.n6817 vdd.n6754 23.783
R41142 vdd.n6818 vdd.n6740 23.783
R41143 vdd.n6818 vdd.n6746 23.783
R41144 vdd.n6819 vdd.n6732 23.783
R41145 vdd.n6819 vdd.n6738 23.783
R41146 vdd.n6820 vdd.n6724 23.783
R41147 vdd.n6820 vdd.n6728 23.783
R41148 vdd.n6821 vdd.n6716 23.783
R41149 vdd.n6821 vdd.n6722 23.783
R41150 vdd.n6822 vdd.n6708 23.783
R41151 vdd.n6822 vdd.n6714 23.783
R41152 vdd.n6823 vdd.n6700 23.783
R41153 vdd.n6823 vdd.n6706 23.783
R41154 vdd.n6824 vdd.n6692 23.783
R41155 vdd.n6824 vdd.n6698 23.783
R41156 vdd.n6825 vdd.n6684 23.783
R41157 vdd.n6825 vdd.n6690 23.783
R41158 vdd.n6826 vdd.n6676 23.783
R41159 vdd.n6826 vdd.n6682 23.783
R41160 vdd.n6827 vdd.n6668 23.783
R41161 vdd.n6827 vdd.n6674 23.783
R41162 vdd.n6828 vdd.n6660 23.783
R41163 vdd.n6828 vdd.n6666 23.783
R41164 vdd.n6839 vdd.n6838 23.783
R41165 vdd.n6839 vdd.n6833 23.783
R41166 vdd.n6990 vdd.n6989 23.783
R41167 vdd.n6990 vdd.n6987 23.783
R41168 vdd.n6991 vdd.n6976 23.783
R41169 vdd.n6991 vdd.n6982 23.783
R41170 vdd.n6992 vdd.n6968 23.783
R41171 vdd.n6992 vdd.n6974 23.783
R41172 vdd.n6993 vdd.n6960 23.783
R41173 vdd.n6993 vdd.n6966 23.783
R41174 vdd.n6994 vdd.n6952 23.783
R41175 vdd.n6994 vdd.n6958 23.783
R41176 vdd.n6995 vdd.n6944 23.783
R41177 vdd.n6995 vdd.n6950 23.783
R41178 vdd.n6996 vdd.n6936 23.783
R41179 vdd.n6996 vdd.n6942 23.783
R41180 vdd.n6997 vdd.n6928 23.783
R41181 vdd.n6997 vdd.n6934 23.783
R41182 vdd.n6998 vdd.n6920 23.783
R41183 vdd.n6998 vdd.n6926 23.783
R41184 vdd.n6999 vdd.n6912 23.783
R41185 vdd.n6999 vdd.n6918 23.783
R41186 vdd.n7000 vdd.n6904 23.783
R41187 vdd.n7000 vdd.n6908 23.783
R41188 vdd.n7001 vdd.n6896 23.783
R41189 vdd.n7001 vdd.n6902 23.783
R41190 vdd.n7002 vdd.n6888 23.783
R41191 vdd.n7002 vdd.n6894 23.783
R41192 vdd.n7003 vdd.n6880 23.783
R41193 vdd.n7003 vdd.n6886 23.783
R41194 vdd.n7004 vdd.n6872 23.783
R41195 vdd.n7004 vdd.n6878 23.783
R41196 vdd.n7005 vdd.n6864 23.783
R41197 vdd.n7005 vdd.n6870 23.783
R41198 vdd.n7006 vdd.n6856 23.783
R41199 vdd.n7006 vdd.n6862 23.783
R41200 vdd.n7007 vdd.n6848 23.783
R41201 vdd.n7007 vdd.n6854 23.783
R41202 vdd.n7008 vdd.n6840 23.783
R41203 vdd.n7008 vdd.n6846 23.783
R41204 vdd.n7019 vdd.n7018 23.783
R41205 vdd.n7019 vdd.n7013 23.783
R41206 vdd.n7170 vdd.n7169 23.783
R41207 vdd.n7170 vdd.n7167 23.783
R41208 vdd.n7171 vdd.n7156 23.783
R41209 vdd.n7171 vdd.n7162 23.783
R41210 vdd.n7172 vdd.n7148 23.783
R41211 vdd.n7172 vdd.n7154 23.783
R41212 vdd.n7173 vdd.n7140 23.783
R41213 vdd.n7173 vdd.n7146 23.783
R41214 vdd.n7174 vdd.n7132 23.783
R41215 vdd.n7174 vdd.n7138 23.783
R41216 vdd.n7175 vdd.n7124 23.783
R41217 vdd.n7175 vdd.n7130 23.783
R41218 vdd.n7176 vdd.n7116 23.783
R41219 vdd.n7176 vdd.n7122 23.783
R41220 vdd.n7177 vdd.n7108 23.783
R41221 vdd.n7177 vdd.n7114 23.783
R41222 vdd.n7178 vdd.n7100 23.783
R41223 vdd.n7178 vdd.n7106 23.783
R41224 vdd.n7179 vdd.n7092 23.783
R41225 vdd.n7179 vdd.n7098 23.783
R41226 vdd.n7180 vdd.n7084 23.783
R41227 vdd.n7180 vdd.n7088 23.783
R41228 vdd.n7181 vdd.n7076 23.783
R41229 vdd.n7181 vdd.n7082 23.783
R41230 vdd.n7182 vdd.n7068 23.783
R41231 vdd.n7182 vdd.n7074 23.783
R41232 vdd.n7183 vdd.n7060 23.783
R41233 vdd.n7183 vdd.n7066 23.783
R41234 vdd.n7184 vdd.n7052 23.783
R41235 vdd.n7184 vdd.n7058 23.783
R41236 vdd.n7185 vdd.n7044 23.783
R41237 vdd.n7185 vdd.n7050 23.783
R41238 vdd.n7186 vdd.n7036 23.783
R41239 vdd.n7186 vdd.n7042 23.783
R41240 vdd.n7187 vdd.n7028 23.783
R41241 vdd.n7187 vdd.n7034 23.783
R41242 vdd.n7188 vdd.n7020 23.783
R41243 vdd.n7188 vdd.n7026 23.783
R41244 vdd.n7199 vdd.n7198 23.783
R41245 vdd.n7199 vdd.n7193 23.783
R41246 vdd.n7350 vdd.n7349 23.783
R41247 vdd.n7350 vdd.n7347 23.783
R41248 vdd.n7351 vdd.n7336 23.783
R41249 vdd.n7351 vdd.n7342 23.783
R41250 vdd.n7352 vdd.n7328 23.783
R41251 vdd.n7352 vdd.n7334 23.783
R41252 vdd.n7353 vdd.n7320 23.783
R41253 vdd.n7353 vdd.n7326 23.783
R41254 vdd.n7354 vdd.n7312 23.783
R41255 vdd.n7354 vdd.n7318 23.783
R41256 vdd.n7355 vdd.n7304 23.783
R41257 vdd.n7355 vdd.n7310 23.783
R41258 vdd.n7356 vdd.n7296 23.783
R41259 vdd.n7356 vdd.n7302 23.783
R41260 vdd.n7357 vdd.n7288 23.783
R41261 vdd.n7357 vdd.n7294 23.783
R41262 vdd.n7358 vdd.n7280 23.783
R41263 vdd.n7358 vdd.n7286 23.783
R41264 vdd.n7359 vdd.n7272 23.783
R41265 vdd.n7359 vdd.n7278 23.783
R41266 vdd.n7360 vdd.n7264 23.783
R41267 vdd.n7360 vdd.n7268 23.783
R41268 vdd.n7361 vdd.n7256 23.783
R41269 vdd.n7361 vdd.n7262 23.783
R41270 vdd.n7362 vdd.n7248 23.783
R41271 vdd.n7362 vdd.n7254 23.783
R41272 vdd.n7363 vdd.n7240 23.783
R41273 vdd.n7363 vdd.n7246 23.783
R41274 vdd.n7364 vdd.n7232 23.783
R41275 vdd.n7364 vdd.n7238 23.783
R41276 vdd.n7365 vdd.n7224 23.783
R41277 vdd.n7365 vdd.n7230 23.783
R41278 vdd.n7366 vdd.n7216 23.783
R41279 vdd.n7366 vdd.n7222 23.783
R41280 vdd.n7367 vdd.n7208 23.783
R41281 vdd.n7367 vdd.n7214 23.783
R41282 vdd.n7368 vdd.n7200 23.783
R41283 vdd.n7368 vdd.n7206 23.783
R41284 vdd.n7379 vdd.n7378 23.783
R41285 vdd.n7379 vdd.n7373 23.783
R41286 vdd.n7530 vdd.n7529 23.783
R41287 vdd.n7530 vdd.n7527 23.783
R41288 vdd.n7531 vdd.n7516 23.783
R41289 vdd.n7531 vdd.n7522 23.783
R41290 vdd.n7532 vdd.n7508 23.783
R41291 vdd.n7532 vdd.n7514 23.783
R41292 vdd.n7533 vdd.n7500 23.783
R41293 vdd.n7533 vdd.n7506 23.783
R41294 vdd.n7534 vdd.n7492 23.783
R41295 vdd.n7534 vdd.n7498 23.783
R41296 vdd.n7535 vdd.n7484 23.783
R41297 vdd.n7535 vdd.n7490 23.783
R41298 vdd.n7536 vdd.n7476 23.783
R41299 vdd.n7536 vdd.n7482 23.783
R41300 vdd.n7537 vdd.n7468 23.783
R41301 vdd.n7537 vdd.n7474 23.783
R41302 vdd.n7538 vdd.n7460 23.783
R41303 vdd.n7538 vdd.n7466 23.783
R41304 vdd.n7539 vdd.n7452 23.783
R41305 vdd.n7539 vdd.n7458 23.783
R41306 vdd.n7540 vdd.n7444 23.783
R41307 vdd.n7540 vdd.n7448 23.783
R41308 vdd.n7541 vdd.n7436 23.783
R41309 vdd.n7541 vdd.n7442 23.783
R41310 vdd.n7542 vdd.n7428 23.783
R41311 vdd.n7542 vdd.n7434 23.783
R41312 vdd.n7543 vdd.n7420 23.783
R41313 vdd.n7543 vdd.n7426 23.783
R41314 vdd.n7544 vdd.n7412 23.783
R41315 vdd.n7544 vdd.n7418 23.783
R41316 vdd.n7545 vdd.n7404 23.783
R41317 vdd.n7545 vdd.n7410 23.783
R41318 vdd.n7546 vdd.n7396 23.783
R41319 vdd.n7546 vdd.n7402 23.783
R41320 vdd.n7547 vdd.n7388 23.783
R41321 vdd.n7547 vdd.n7394 23.783
R41322 vdd.n7548 vdd.n7380 23.783
R41323 vdd.n7548 vdd.n7386 23.783
R41324 vdd.n7559 vdd.n7558 23.783
R41325 vdd.n7559 vdd.n7553 23.783
R41326 vdd.n7710 vdd.n7709 23.783
R41327 vdd.n7710 vdd.n7707 23.783
R41328 vdd.n7711 vdd.n7696 23.783
R41329 vdd.n7711 vdd.n7702 23.783
R41330 vdd.n7712 vdd.n7688 23.783
R41331 vdd.n7712 vdd.n7694 23.783
R41332 vdd.n7713 vdd.n7680 23.783
R41333 vdd.n7713 vdd.n7686 23.783
R41334 vdd.n7714 vdd.n7672 23.783
R41335 vdd.n7714 vdd.n7678 23.783
R41336 vdd.n7715 vdd.n7664 23.783
R41337 vdd.n7715 vdd.n7670 23.783
R41338 vdd.n7716 vdd.n7656 23.783
R41339 vdd.n7716 vdd.n7662 23.783
R41340 vdd.n7717 vdd.n7648 23.783
R41341 vdd.n7717 vdd.n7654 23.783
R41342 vdd.n7718 vdd.n7640 23.783
R41343 vdd.n7718 vdd.n7646 23.783
R41344 vdd.n7719 vdd.n7632 23.783
R41345 vdd.n7719 vdd.n7638 23.783
R41346 vdd.n7720 vdd.n7624 23.783
R41347 vdd.n7720 vdd.n7628 23.783
R41348 vdd.n7721 vdd.n7616 23.783
R41349 vdd.n7721 vdd.n7622 23.783
R41350 vdd.n7722 vdd.n7608 23.783
R41351 vdd.n7722 vdd.n7614 23.783
R41352 vdd.n7723 vdd.n7600 23.783
R41353 vdd.n7723 vdd.n7606 23.783
R41354 vdd.n7724 vdd.n7592 23.783
R41355 vdd.n7724 vdd.n7598 23.783
R41356 vdd.n7725 vdd.n7584 23.783
R41357 vdd.n7725 vdd.n7590 23.783
R41358 vdd.n7726 vdd.n7576 23.783
R41359 vdd.n7726 vdd.n7582 23.783
R41360 vdd.n7727 vdd.n7568 23.783
R41361 vdd.n7727 vdd.n7574 23.783
R41362 vdd.n7728 vdd.n7560 23.783
R41363 vdd.n7728 vdd.n7566 23.783
R41364 vdd.n7739 vdd.n7738 23.783
R41365 vdd.n7739 vdd.n7733 23.783
R41366 vdd.n7890 vdd.n7889 23.783
R41367 vdd.n7890 vdd.n7887 23.783
R41368 vdd.n7891 vdd.n7876 23.783
R41369 vdd.n7891 vdd.n7882 23.783
R41370 vdd.n7892 vdd.n7868 23.783
R41371 vdd.n7892 vdd.n7874 23.783
R41372 vdd.n7893 vdd.n7860 23.783
R41373 vdd.n7893 vdd.n7866 23.783
R41374 vdd.n7894 vdd.n7852 23.783
R41375 vdd.n7894 vdd.n7858 23.783
R41376 vdd.n7895 vdd.n7844 23.783
R41377 vdd.n7895 vdd.n7850 23.783
R41378 vdd.n7896 vdd.n7836 23.783
R41379 vdd.n7896 vdd.n7842 23.783
R41380 vdd.n7897 vdd.n7828 23.783
R41381 vdd.n7897 vdd.n7834 23.783
R41382 vdd.n7898 vdd.n7820 23.783
R41383 vdd.n7898 vdd.n7826 23.783
R41384 vdd.n7899 vdd.n7812 23.783
R41385 vdd.n7899 vdd.n7818 23.783
R41386 vdd.n7900 vdd.n7804 23.783
R41387 vdd.n7900 vdd.n7808 23.783
R41388 vdd.n7901 vdd.n7796 23.783
R41389 vdd.n7901 vdd.n7802 23.783
R41390 vdd.n7902 vdd.n7788 23.783
R41391 vdd.n7902 vdd.n7794 23.783
R41392 vdd.n7903 vdd.n7780 23.783
R41393 vdd.n7903 vdd.n7786 23.783
R41394 vdd.n7904 vdd.n7772 23.783
R41395 vdd.n7904 vdd.n7778 23.783
R41396 vdd.n7905 vdd.n7764 23.783
R41397 vdd.n7905 vdd.n7770 23.783
R41398 vdd.n7906 vdd.n7756 23.783
R41399 vdd.n7906 vdd.n7762 23.783
R41400 vdd.n7907 vdd.n7748 23.783
R41401 vdd.n7907 vdd.n7754 23.783
R41402 vdd.n7908 vdd.n7740 23.783
R41403 vdd.n7908 vdd.n7746 23.783
R41404 vdd.n7919 vdd.n7918 23.783
R41405 vdd.n7919 vdd.n7913 23.783
R41406 vdd.n8070 vdd.n8069 23.783
R41407 vdd.n8070 vdd.n8067 23.783
R41408 vdd.n8071 vdd.n8056 23.783
R41409 vdd.n8071 vdd.n8062 23.783
R41410 vdd.n8072 vdd.n8048 23.783
R41411 vdd.n8072 vdd.n8054 23.783
R41412 vdd.n8073 vdd.n8040 23.783
R41413 vdd.n8073 vdd.n8046 23.783
R41414 vdd.n8074 vdd.n8032 23.783
R41415 vdd.n8074 vdd.n8038 23.783
R41416 vdd.n8075 vdd.n8024 23.783
R41417 vdd.n8075 vdd.n8030 23.783
R41418 vdd.n8076 vdd.n8016 23.783
R41419 vdd.n8076 vdd.n8022 23.783
R41420 vdd.n8077 vdd.n8008 23.783
R41421 vdd.n8077 vdd.n8014 23.783
R41422 vdd.n8078 vdd.n8000 23.783
R41423 vdd.n8078 vdd.n8006 23.783
R41424 vdd.n8079 vdd.n7992 23.783
R41425 vdd.n8079 vdd.n7998 23.783
R41426 vdd.n8080 vdd.n7984 23.783
R41427 vdd.n8080 vdd.n7988 23.783
R41428 vdd.n8081 vdd.n7976 23.783
R41429 vdd.n8081 vdd.n7982 23.783
R41430 vdd.n8082 vdd.n7968 23.783
R41431 vdd.n8082 vdd.n7974 23.783
R41432 vdd.n8083 vdd.n7960 23.783
R41433 vdd.n8083 vdd.n7966 23.783
R41434 vdd.n8084 vdd.n7952 23.783
R41435 vdd.n8084 vdd.n7958 23.783
R41436 vdd.n8085 vdd.n7944 23.783
R41437 vdd.n8085 vdd.n7950 23.783
R41438 vdd.n8086 vdd.n7936 23.783
R41439 vdd.n8086 vdd.n7942 23.783
R41440 vdd.n8087 vdd.n7928 23.783
R41441 vdd.n8087 vdd.n7934 23.783
R41442 vdd.n8088 vdd.n7920 23.783
R41443 vdd.n8088 vdd.n7926 23.783
R41444 vdd.n8099 vdd.n8098 23.783
R41445 vdd.n8099 vdd.n8093 23.783
R41446 vdd.n8250 vdd.n8249 23.783
R41447 vdd.n8250 vdd.n8247 23.783
R41448 vdd.n8251 vdd.n8236 23.783
R41449 vdd.n8251 vdd.n8242 23.783
R41450 vdd.n8252 vdd.n8228 23.783
R41451 vdd.n8252 vdd.n8234 23.783
R41452 vdd.n8253 vdd.n8220 23.783
R41453 vdd.n8253 vdd.n8226 23.783
R41454 vdd.n8254 vdd.n8212 23.783
R41455 vdd.n8254 vdd.n8218 23.783
R41456 vdd.n8255 vdd.n8204 23.783
R41457 vdd.n8255 vdd.n8210 23.783
R41458 vdd.n8256 vdd.n8196 23.783
R41459 vdd.n8256 vdd.n8202 23.783
R41460 vdd.n8257 vdd.n8188 23.783
R41461 vdd.n8257 vdd.n8194 23.783
R41462 vdd.n8258 vdd.n8180 23.783
R41463 vdd.n8258 vdd.n8186 23.783
R41464 vdd.n8259 vdd.n8172 23.783
R41465 vdd.n8259 vdd.n8178 23.783
R41466 vdd.n8260 vdd.n8164 23.783
R41467 vdd.n8260 vdd.n8168 23.783
R41468 vdd.n8261 vdd.n8156 23.783
R41469 vdd.n8261 vdd.n8162 23.783
R41470 vdd.n8262 vdd.n8148 23.783
R41471 vdd.n8262 vdd.n8154 23.783
R41472 vdd.n8263 vdd.n8140 23.783
R41473 vdd.n8263 vdd.n8146 23.783
R41474 vdd.n8264 vdd.n8132 23.783
R41475 vdd.n8264 vdd.n8138 23.783
R41476 vdd.n8265 vdd.n8124 23.783
R41477 vdd.n8265 vdd.n8130 23.783
R41478 vdd.n8266 vdd.n8116 23.783
R41479 vdd.n8266 vdd.n8122 23.783
R41480 vdd.n8267 vdd.n8108 23.783
R41481 vdd.n8267 vdd.n8114 23.783
R41482 vdd.n8268 vdd.n8100 23.783
R41483 vdd.n8268 vdd.n8106 23.783
R41484 vdd.n8279 vdd.n8278 23.783
R41485 vdd.n8279 vdd.n8273 23.783
R41486 vdd.n8430 vdd.n8429 23.783
R41487 vdd.n8430 vdd.n8427 23.783
R41488 vdd.n8431 vdd.n8416 23.783
R41489 vdd.n8431 vdd.n8422 23.783
R41490 vdd.n8432 vdd.n8408 23.783
R41491 vdd.n8432 vdd.n8414 23.783
R41492 vdd.n8433 vdd.n8400 23.783
R41493 vdd.n8433 vdd.n8406 23.783
R41494 vdd.n8434 vdd.n8392 23.783
R41495 vdd.n8434 vdd.n8398 23.783
R41496 vdd.n8435 vdd.n8384 23.783
R41497 vdd.n8435 vdd.n8390 23.783
R41498 vdd.n8436 vdd.n8376 23.783
R41499 vdd.n8436 vdd.n8382 23.783
R41500 vdd.n8437 vdd.n8368 23.783
R41501 vdd.n8437 vdd.n8374 23.783
R41502 vdd.n8438 vdd.n8360 23.783
R41503 vdd.n8438 vdd.n8366 23.783
R41504 vdd.n8439 vdd.n8352 23.783
R41505 vdd.n8439 vdd.n8358 23.783
R41506 vdd.n8440 vdd.n8344 23.783
R41507 vdd.n8440 vdd.n8348 23.783
R41508 vdd.n8441 vdd.n8336 23.783
R41509 vdd.n8441 vdd.n8342 23.783
R41510 vdd.n8442 vdd.n8328 23.783
R41511 vdd.n8442 vdd.n8334 23.783
R41512 vdd.n8443 vdd.n8320 23.783
R41513 vdd.n8443 vdd.n8326 23.783
R41514 vdd.n8444 vdd.n8312 23.783
R41515 vdd.n8444 vdd.n8318 23.783
R41516 vdd.n8445 vdd.n8304 23.783
R41517 vdd.n8445 vdd.n8310 23.783
R41518 vdd.n8446 vdd.n8296 23.783
R41519 vdd.n8446 vdd.n8302 23.783
R41520 vdd.n8447 vdd.n8288 23.783
R41521 vdd.n8447 vdd.n8294 23.783
R41522 vdd.n8448 vdd.n8280 23.783
R41523 vdd.n8448 vdd.n8286 23.783
R41524 vdd.n8459 vdd.n8458 23.783
R41525 vdd.n8459 vdd.n8453 23.783
R41526 vdd.n8610 vdd.n8609 23.783
R41527 vdd.n8610 vdd.n8607 23.783
R41528 vdd.n8611 vdd.n8596 23.783
R41529 vdd.n8611 vdd.n8602 23.783
R41530 vdd.n8612 vdd.n8588 23.783
R41531 vdd.n8612 vdd.n8594 23.783
R41532 vdd.n8613 vdd.n8580 23.783
R41533 vdd.n8613 vdd.n8586 23.783
R41534 vdd.n8614 vdd.n8572 23.783
R41535 vdd.n8614 vdd.n8578 23.783
R41536 vdd.n8615 vdd.n8564 23.783
R41537 vdd.n8615 vdd.n8570 23.783
R41538 vdd.n8616 vdd.n8556 23.783
R41539 vdd.n8616 vdd.n8562 23.783
R41540 vdd.n8617 vdd.n8548 23.783
R41541 vdd.n8617 vdd.n8554 23.783
R41542 vdd.n8618 vdd.n8540 23.783
R41543 vdd.n8618 vdd.n8546 23.783
R41544 vdd.n8619 vdd.n8532 23.783
R41545 vdd.n8619 vdd.n8538 23.783
R41546 vdd.n8620 vdd.n8524 23.783
R41547 vdd.n8620 vdd.n8528 23.783
R41548 vdd.n8621 vdd.n8516 23.783
R41549 vdd.n8621 vdd.n8522 23.783
R41550 vdd.n8622 vdd.n8508 23.783
R41551 vdd.n8622 vdd.n8514 23.783
R41552 vdd.n8623 vdd.n8500 23.783
R41553 vdd.n8623 vdd.n8506 23.783
R41554 vdd.n8624 vdd.n8492 23.783
R41555 vdd.n8624 vdd.n8498 23.783
R41556 vdd.n8625 vdd.n8484 23.783
R41557 vdd.n8625 vdd.n8490 23.783
R41558 vdd.n8626 vdd.n8476 23.783
R41559 vdd.n8626 vdd.n8482 23.783
R41560 vdd.n8627 vdd.n8468 23.783
R41561 vdd.n8627 vdd.n8474 23.783
R41562 vdd.n8628 vdd.n8460 23.783
R41563 vdd.n8628 vdd.n8466 23.783
R41564 vdd.n8639 vdd.n8638 23.783
R41565 vdd.n8639 vdd.n8633 23.783
R41566 vdd.n8790 vdd.n8789 23.783
R41567 vdd.n8790 vdd.n8787 23.783
R41568 vdd.n8791 vdd.n8776 23.783
R41569 vdd.n8791 vdd.n8782 23.783
R41570 vdd.n8792 vdd.n8768 23.783
R41571 vdd.n8792 vdd.n8774 23.783
R41572 vdd.n8793 vdd.n8760 23.783
R41573 vdd.n8793 vdd.n8766 23.783
R41574 vdd.n8794 vdd.n8752 23.783
R41575 vdd.n8794 vdd.n8758 23.783
R41576 vdd.n8795 vdd.n8744 23.783
R41577 vdd.n8795 vdd.n8750 23.783
R41578 vdd.n8796 vdd.n8736 23.783
R41579 vdd.n8796 vdd.n8742 23.783
R41580 vdd.n8797 vdd.n8728 23.783
R41581 vdd.n8797 vdd.n8734 23.783
R41582 vdd.n8798 vdd.n8720 23.783
R41583 vdd.n8798 vdd.n8726 23.783
R41584 vdd.n8799 vdd.n8712 23.783
R41585 vdd.n8799 vdd.n8718 23.783
R41586 vdd.n8800 vdd.n8704 23.783
R41587 vdd.n8800 vdd.n8708 23.783
R41588 vdd.n8801 vdd.n8696 23.783
R41589 vdd.n8801 vdd.n8702 23.783
R41590 vdd.n8802 vdd.n8688 23.783
R41591 vdd.n8802 vdd.n8694 23.783
R41592 vdd.n8803 vdd.n8680 23.783
R41593 vdd.n8803 vdd.n8686 23.783
R41594 vdd.n8804 vdd.n8672 23.783
R41595 vdd.n8804 vdd.n8678 23.783
R41596 vdd.n8805 vdd.n8664 23.783
R41597 vdd.n8805 vdd.n8670 23.783
R41598 vdd.n8806 vdd.n8656 23.783
R41599 vdd.n8806 vdd.n8662 23.783
R41600 vdd.n8807 vdd.n8648 23.783
R41601 vdd.n8807 vdd.n8654 23.783
R41602 vdd.n8808 vdd.n8640 23.783
R41603 vdd.n8808 vdd.n8646 23.783
R41604 vdd.n8819 vdd.n8818 23.783
R41605 vdd.n8819 vdd.n8813 23.783
R41606 vdd.n8970 vdd.n8969 23.783
R41607 vdd.n8970 vdd.n8967 23.783
R41608 vdd.n8971 vdd.n8956 23.783
R41609 vdd.n8971 vdd.n8962 23.783
R41610 vdd.n8972 vdd.n8948 23.783
R41611 vdd.n8972 vdd.n8954 23.783
R41612 vdd.n8973 vdd.n8940 23.783
R41613 vdd.n8973 vdd.n8946 23.783
R41614 vdd.n8974 vdd.n8932 23.783
R41615 vdd.n8974 vdd.n8938 23.783
R41616 vdd.n8975 vdd.n8924 23.783
R41617 vdd.n8975 vdd.n8930 23.783
R41618 vdd.n8976 vdd.n8916 23.783
R41619 vdd.n8976 vdd.n8922 23.783
R41620 vdd.n8977 vdd.n8908 23.783
R41621 vdd.n8977 vdd.n8914 23.783
R41622 vdd.n8978 vdd.n8900 23.783
R41623 vdd.n8978 vdd.n8906 23.783
R41624 vdd.n8979 vdd.n8892 23.783
R41625 vdd.n8979 vdd.n8898 23.783
R41626 vdd.n8980 vdd.n8884 23.783
R41627 vdd.n8980 vdd.n8888 23.783
R41628 vdd.n8981 vdd.n8876 23.783
R41629 vdd.n8981 vdd.n8882 23.783
R41630 vdd.n8982 vdd.n8868 23.783
R41631 vdd.n8982 vdd.n8874 23.783
R41632 vdd.n8983 vdd.n8860 23.783
R41633 vdd.n8983 vdd.n8866 23.783
R41634 vdd.n8984 vdd.n8852 23.783
R41635 vdd.n8984 vdd.n8858 23.783
R41636 vdd.n8985 vdd.n8844 23.783
R41637 vdd.n8985 vdd.n8850 23.783
R41638 vdd.n8986 vdd.n8836 23.783
R41639 vdd.n8986 vdd.n8842 23.783
R41640 vdd.n8987 vdd.n8828 23.783
R41641 vdd.n8987 vdd.n8834 23.783
R41642 vdd.n8988 vdd.n8820 23.783
R41643 vdd.n8988 vdd.n8826 23.783
R41644 vdd.n8999 vdd.n8998 23.783
R41645 vdd.n8999 vdd.n8993 23.783
R41646 vdd.n9150 vdd.n9149 23.783
R41647 vdd.n9150 vdd.n9147 23.783
R41648 vdd.n9151 vdd.n9136 23.783
R41649 vdd.n9151 vdd.n9142 23.783
R41650 vdd.n9152 vdd.n9128 23.783
R41651 vdd.n9152 vdd.n9134 23.783
R41652 vdd.n9153 vdd.n9120 23.783
R41653 vdd.n9153 vdd.n9126 23.783
R41654 vdd.n9154 vdd.n9112 23.783
R41655 vdd.n9154 vdd.n9118 23.783
R41656 vdd.n9155 vdd.n9104 23.783
R41657 vdd.n9155 vdd.n9110 23.783
R41658 vdd.n9156 vdd.n9096 23.783
R41659 vdd.n9156 vdd.n9102 23.783
R41660 vdd.n9157 vdd.n9088 23.783
R41661 vdd.n9157 vdd.n9094 23.783
R41662 vdd.n9158 vdd.n9080 23.783
R41663 vdd.n9158 vdd.n9086 23.783
R41664 vdd.n9159 vdd.n9072 23.783
R41665 vdd.n9159 vdd.n9078 23.783
R41666 vdd.n9160 vdd.n9064 23.783
R41667 vdd.n9160 vdd.n9068 23.783
R41668 vdd.n9161 vdd.n9056 23.783
R41669 vdd.n9161 vdd.n9062 23.783
R41670 vdd.n9162 vdd.n9048 23.783
R41671 vdd.n9162 vdd.n9054 23.783
R41672 vdd.n9163 vdd.n9040 23.783
R41673 vdd.n9163 vdd.n9046 23.783
R41674 vdd.n9164 vdd.n9032 23.783
R41675 vdd.n9164 vdd.n9038 23.783
R41676 vdd.n9165 vdd.n9024 23.783
R41677 vdd.n9165 vdd.n9030 23.783
R41678 vdd.n9166 vdd.n9016 23.783
R41679 vdd.n9166 vdd.n9022 23.783
R41680 vdd.n9167 vdd.n9008 23.783
R41681 vdd.n9167 vdd.n9014 23.783
R41682 vdd.n9168 vdd.n9000 23.783
R41683 vdd.n9168 vdd.n9006 23.783
R41684 vdd.n9179 vdd.n9178 23.783
R41685 vdd.n9179 vdd.n9173 23.783
R41686 vdd.n9330 vdd.n9329 23.783
R41687 vdd.n9330 vdd.n9327 23.783
R41688 vdd.n9331 vdd.n9316 23.783
R41689 vdd.n9331 vdd.n9322 23.783
R41690 vdd.n9332 vdd.n9308 23.783
R41691 vdd.n9332 vdd.n9314 23.783
R41692 vdd.n9333 vdd.n9300 23.783
R41693 vdd.n9333 vdd.n9306 23.783
R41694 vdd.n9334 vdd.n9292 23.783
R41695 vdd.n9334 vdd.n9298 23.783
R41696 vdd.n9335 vdd.n9284 23.783
R41697 vdd.n9335 vdd.n9290 23.783
R41698 vdd.n9336 vdd.n9276 23.783
R41699 vdd.n9336 vdd.n9282 23.783
R41700 vdd.n9337 vdd.n9268 23.783
R41701 vdd.n9337 vdd.n9274 23.783
R41702 vdd.n9338 vdd.n9260 23.783
R41703 vdd.n9338 vdd.n9266 23.783
R41704 vdd.n9339 vdd.n9252 23.783
R41705 vdd.n9339 vdd.n9258 23.783
R41706 vdd.n9340 vdd.n9244 23.783
R41707 vdd.n9340 vdd.n9248 23.783
R41708 vdd.n9341 vdd.n9236 23.783
R41709 vdd.n9341 vdd.n9242 23.783
R41710 vdd.n9342 vdd.n9228 23.783
R41711 vdd.n9342 vdd.n9234 23.783
R41712 vdd.n9343 vdd.n9220 23.783
R41713 vdd.n9343 vdd.n9226 23.783
R41714 vdd.n9344 vdd.n9212 23.783
R41715 vdd.n9344 vdd.n9218 23.783
R41716 vdd.n9345 vdd.n9204 23.783
R41717 vdd.n9345 vdd.n9210 23.783
R41718 vdd.n9346 vdd.n9196 23.783
R41719 vdd.n9346 vdd.n9202 23.783
R41720 vdd.n9347 vdd.n9188 23.783
R41721 vdd.n9347 vdd.n9194 23.783
R41722 vdd.n9348 vdd.n9180 23.783
R41723 vdd.n9348 vdd.n9186 23.783
R41724 vdd.n9359 vdd.n9358 23.783
R41725 vdd.n9359 vdd.n9353 23.783
R41726 vdd.n9510 vdd.n9509 23.783
R41727 vdd.n9510 vdd.n9507 23.783
R41728 vdd.n9511 vdd.n9496 23.783
R41729 vdd.n9511 vdd.n9502 23.783
R41730 vdd.n9512 vdd.n9488 23.783
R41731 vdd.n9512 vdd.n9494 23.783
R41732 vdd.n9513 vdd.n9480 23.783
R41733 vdd.n9513 vdd.n9486 23.783
R41734 vdd.n9514 vdd.n9472 23.783
R41735 vdd.n9514 vdd.n9478 23.783
R41736 vdd.n9515 vdd.n9464 23.783
R41737 vdd.n9515 vdd.n9470 23.783
R41738 vdd.n9516 vdd.n9456 23.783
R41739 vdd.n9516 vdd.n9462 23.783
R41740 vdd.n9517 vdd.n9448 23.783
R41741 vdd.n9517 vdd.n9454 23.783
R41742 vdd.n9518 vdd.n9440 23.783
R41743 vdd.n9518 vdd.n9446 23.783
R41744 vdd.n9519 vdd.n9432 23.783
R41745 vdd.n9519 vdd.n9438 23.783
R41746 vdd.n9520 vdd.n9424 23.783
R41747 vdd.n9520 vdd.n9428 23.783
R41748 vdd.n9521 vdd.n9416 23.783
R41749 vdd.n9521 vdd.n9422 23.783
R41750 vdd.n9522 vdd.n9408 23.783
R41751 vdd.n9522 vdd.n9414 23.783
R41752 vdd.n9523 vdd.n9400 23.783
R41753 vdd.n9523 vdd.n9406 23.783
R41754 vdd.n9524 vdd.n9392 23.783
R41755 vdd.n9524 vdd.n9398 23.783
R41756 vdd.n9525 vdd.n9384 23.783
R41757 vdd.n9525 vdd.n9390 23.783
R41758 vdd.n9526 vdd.n9376 23.783
R41759 vdd.n9526 vdd.n9382 23.783
R41760 vdd.n9527 vdd.n9368 23.783
R41761 vdd.n9527 vdd.n9374 23.783
R41762 vdd.n9528 vdd.n9360 23.783
R41763 vdd.n9528 vdd.n9366 23.783
R41764 vdd.n9539 vdd.n9538 23.783
R41765 vdd.n9539 vdd.n9533 23.783
R41766 vdd.n9690 vdd.n9689 23.783
R41767 vdd.n9690 vdd.n9687 23.783
R41768 vdd.n9691 vdd.n9676 23.783
R41769 vdd.n9691 vdd.n9682 23.783
R41770 vdd.n9692 vdd.n9668 23.783
R41771 vdd.n9692 vdd.n9674 23.783
R41772 vdd.n9693 vdd.n9660 23.783
R41773 vdd.n9693 vdd.n9666 23.783
R41774 vdd.n9694 vdd.n9652 23.783
R41775 vdd.n9694 vdd.n9658 23.783
R41776 vdd.n9695 vdd.n9644 23.783
R41777 vdd.n9695 vdd.n9650 23.783
R41778 vdd.n9696 vdd.n9636 23.783
R41779 vdd.n9696 vdd.n9642 23.783
R41780 vdd.n9697 vdd.n9628 23.783
R41781 vdd.n9697 vdd.n9634 23.783
R41782 vdd.n9698 vdd.n9620 23.783
R41783 vdd.n9698 vdd.n9626 23.783
R41784 vdd.n9699 vdd.n9612 23.783
R41785 vdd.n9699 vdd.n9618 23.783
R41786 vdd.n9700 vdd.n9604 23.783
R41787 vdd.n9700 vdd.n9608 23.783
R41788 vdd.n9701 vdd.n9596 23.783
R41789 vdd.n9701 vdd.n9602 23.783
R41790 vdd.n9702 vdd.n9588 23.783
R41791 vdd.n9702 vdd.n9594 23.783
R41792 vdd.n9703 vdd.n9580 23.783
R41793 vdd.n9703 vdd.n9586 23.783
R41794 vdd.n9704 vdd.n9572 23.783
R41795 vdd.n9704 vdd.n9578 23.783
R41796 vdd.n9705 vdd.n9564 23.783
R41797 vdd.n9705 vdd.n9570 23.783
R41798 vdd.n9706 vdd.n9556 23.783
R41799 vdd.n9706 vdd.n9562 23.783
R41800 vdd.n9707 vdd.n9548 23.783
R41801 vdd.n9707 vdd.n9554 23.783
R41802 vdd.n9708 vdd.n9540 23.783
R41803 vdd.n9708 vdd.n9546 23.783
R41804 vdd.n9719 vdd.n9718 23.783
R41805 vdd.n9719 vdd.n9713 23.783
R41806 vdd.n9870 vdd.n9869 23.783
R41807 vdd.n9870 vdd.n9867 23.783
R41808 vdd.n9871 vdd.n9856 23.783
R41809 vdd.n9871 vdd.n9862 23.783
R41810 vdd.n9872 vdd.n9848 23.783
R41811 vdd.n9872 vdd.n9854 23.783
R41812 vdd.n9873 vdd.n9840 23.783
R41813 vdd.n9873 vdd.n9846 23.783
R41814 vdd.n9874 vdd.n9832 23.783
R41815 vdd.n9874 vdd.n9838 23.783
R41816 vdd.n9875 vdd.n9824 23.783
R41817 vdd.n9875 vdd.n9830 23.783
R41818 vdd.n9876 vdd.n9816 23.783
R41819 vdd.n9876 vdd.n9822 23.783
R41820 vdd.n9877 vdd.n9808 23.783
R41821 vdd.n9877 vdd.n9814 23.783
R41822 vdd.n9878 vdd.n9800 23.783
R41823 vdd.n9878 vdd.n9806 23.783
R41824 vdd.n9879 vdd.n9792 23.783
R41825 vdd.n9879 vdd.n9798 23.783
R41826 vdd.n9880 vdd.n9784 23.783
R41827 vdd.n9880 vdd.n9788 23.783
R41828 vdd.n9881 vdd.n9776 23.783
R41829 vdd.n9881 vdd.n9782 23.783
R41830 vdd.n9882 vdd.n9768 23.783
R41831 vdd.n9882 vdd.n9774 23.783
R41832 vdd.n9883 vdd.n9760 23.783
R41833 vdd.n9883 vdd.n9766 23.783
R41834 vdd.n9884 vdd.n9752 23.783
R41835 vdd.n9884 vdd.n9758 23.783
R41836 vdd.n9885 vdd.n9744 23.783
R41837 vdd.n9885 vdd.n9750 23.783
R41838 vdd.n9886 vdd.n9736 23.783
R41839 vdd.n9886 vdd.n9742 23.783
R41840 vdd.n9887 vdd.n9728 23.783
R41841 vdd.n9887 vdd.n9734 23.783
R41842 vdd.n9888 vdd.n9720 23.783
R41843 vdd.n9888 vdd.n9726 23.783
R41844 vdd.n9899 vdd.n9898 23.783
R41845 vdd.n9899 vdd.n9893 23.783
R41846 vdd.n10050 vdd.n10049 23.783
R41847 vdd.n10050 vdd.n10047 23.783
R41848 vdd.n10051 vdd.n10036 23.783
R41849 vdd.n10051 vdd.n10042 23.783
R41850 vdd.n10052 vdd.n10028 23.783
R41851 vdd.n10052 vdd.n10034 23.783
R41852 vdd.n10053 vdd.n10020 23.783
R41853 vdd.n10053 vdd.n10026 23.783
R41854 vdd.n10054 vdd.n10012 23.783
R41855 vdd.n10054 vdd.n10018 23.783
R41856 vdd.n10055 vdd.n10004 23.783
R41857 vdd.n10055 vdd.n10010 23.783
R41858 vdd.n10056 vdd.n9996 23.783
R41859 vdd.n10056 vdd.n10002 23.783
R41860 vdd.n10057 vdd.n9988 23.783
R41861 vdd.n10057 vdd.n9994 23.783
R41862 vdd.n10058 vdd.n9980 23.783
R41863 vdd.n10058 vdd.n9986 23.783
R41864 vdd.n10059 vdd.n9972 23.783
R41865 vdd.n10059 vdd.n9978 23.783
R41866 vdd.n10060 vdd.n9964 23.783
R41867 vdd.n10060 vdd.n9968 23.783
R41868 vdd.n10061 vdd.n9956 23.783
R41869 vdd.n10061 vdd.n9962 23.783
R41870 vdd.n10062 vdd.n9948 23.783
R41871 vdd.n10062 vdd.n9954 23.783
R41872 vdd.n10063 vdd.n9940 23.783
R41873 vdd.n10063 vdd.n9946 23.783
R41874 vdd.n10064 vdd.n9932 23.783
R41875 vdd.n10064 vdd.n9938 23.783
R41876 vdd.n10065 vdd.n9924 23.783
R41877 vdd.n10065 vdd.n9930 23.783
R41878 vdd.n10066 vdd.n9916 23.783
R41879 vdd.n10066 vdd.n9922 23.783
R41880 vdd.n10067 vdd.n9908 23.783
R41881 vdd.n10067 vdd.n9914 23.783
R41882 vdd.n10068 vdd.n9900 23.783
R41883 vdd.n10068 vdd.n9906 23.783
R41884 vdd.n10079 vdd.n10078 23.783
R41885 vdd.n10079 vdd.n10073 23.783
R41886 vdd.n10230 vdd.n10229 23.783
R41887 vdd.n10230 vdd.n10227 23.783
R41888 vdd.n10231 vdd.n10216 23.783
R41889 vdd.n10231 vdd.n10222 23.783
R41890 vdd.n10232 vdd.n10208 23.783
R41891 vdd.n10232 vdd.n10214 23.783
R41892 vdd.n10233 vdd.n10200 23.783
R41893 vdd.n10233 vdd.n10206 23.783
R41894 vdd.n10234 vdd.n10192 23.783
R41895 vdd.n10234 vdd.n10198 23.783
R41896 vdd.n10235 vdd.n10184 23.783
R41897 vdd.n10235 vdd.n10190 23.783
R41898 vdd.n10236 vdd.n10176 23.783
R41899 vdd.n10236 vdd.n10182 23.783
R41900 vdd.n10237 vdd.n10168 23.783
R41901 vdd.n10237 vdd.n10174 23.783
R41902 vdd.n10238 vdd.n10160 23.783
R41903 vdd.n10238 vdd.n10166 23.783
R41904 vdd.n10239 vdd.n10152 23.783
R41905 vdd.n10239 vdd.n10158 23.783
R41906 vdd.n10240 vdd.n10144 23.783
R41907 vdd.n10240 vdd.n10148 23.783
R41908 vdd.n10241 vdd.n10136 23.783
R41909 vdd.n10241 vdd.n10142 23.783
R41910 vdd.n10242 vdd.n10128 23.783
R41911 vdd.n10242 vdd.n10134 23.783
R41912 vdd.n10243 vdd.n10120 23.783
R41913 vdd.n10243 vdd.n10126 23.783
R41914 vdd.n10244 vdd.n10112 23.783
R41915 vdd.n10244 vdd.n10118 23.783
R41916 vdd.n10245 vdd.n10104 23.783
R41917 vdd.n10245 vdd.n10110 23.783
R41918 vdd.n10246 vdd.n10096 23.783
R41919 vdd.n10246 vdd.n10102 23.783
R41920 vdd.n10247 vdd.n10088 23.783
R41921 vdd.n10247 vdd.n10094 23.783
R41922 vdd.n10248 vdd.n10080 23.783
R41923 vdd.n10248 vdd.n10086 23.783
R41924 vdd.n10259 vdd.n10258 23.783
R41925 vdd.n10259 vdd.n10253 23.783
R41926 vdd.n10410 vdd.n10409 23.783
R41927 vdd.n10410 vdd.n10407 23.783
R41928 vdd.n10411 vdd.n10396 23.783
R41929 vdd.n10411 vdd.n10402 23.783
R41930 vdd.n10412 vdd.n10388 23.783
R41931 vdd.n10412 vdd.n10394 23.783
R41932 vdd.n10413 vdd.n10380 23.783
R41933 vdd.n10413 vdd.n10386 23.783
R41934 vdd.n10414 vdd.n10372 23.783
R41935 vdd.n10414 vdd.n10378 23.783
R41936 vdd.n10415 vdd.n10364 23.783
R41937 vdd.n10415 vdd.n10370 23.783
R41938 vdd.n10416 vdd.n10356 23.783
R41939 vdd.n10416 vdd.n10362 23.783
R41940 vdd.n10417 vdd.n10348 23.783
R41941 vdd.n10417 vdd.n10354 23.783
R41942 vdd.n10418 vdd.n10340 23.783
R41943 vdd.n10418 vdd.n10346 23.783
R41944 vdd.n10419 vdd.n10332 23.783
R41945 vdd.n10419 vdd.n10338 23.783
R41946 vdd.n10420 vdd.n10324 23.783
R41947 vdd.n10420 vdd.n10328 23.783
R41948 vdd.n10421 vdd.n10316 23.783
R41949 vdd.n10421 vdd.n10322 23.783
R41950 vdd.n10422 vdd.n10308 23.783
R41951 vdd.n10422 vdd.n10314 23.783
R41952 vdd.n10423 vdd.n10300 23.783
R41953 vdd.n10423 vdd.n10306 23.783
R41954 vdd.n10424 vdd.n10292 23.783
R41955 vdd.n10424 vdd.n10298 23.783
R41956 vdd.n10425 vdd.n10284 23.783
R41957 vdd.n10425 vdd.n10290 23.783
R41958 vdd.n10426 vdd.n10276 23.783
R41959 vdd.n10426 vdd.n10282 23.783
R41960 vdd.n10427 vdd.n10268 23.783
R41961 vdd.n10427 vdd.n10274 23.783
R41962 vdd.n10428 vdd.n10260 23.783
R41963 vdd.n10428 vdd.n10266 23.783
R41964 vdd.n10439 vdd.n10438 23.783
R41965 vdd.n10439 vdd.n10433 23.783
R41966 vdd.n10590 vdd.n10589 23.783
R41967 vdd.n10590 vdd.n10587 23.783
R41968 vdd.n10591 vdd.n10576 23.783
R41969 vdd.n10591 vdd.n10582 23.783
R41970 vdd.n10592 vdd.n10568 23.783
R41971 vdd.n10592 vdd.n10574 23.783
R41972 vdd.n10593 vdd.n10560 23.783
R41973 vdd.n10593 vdd.n10566 23.783
R41974 vdd.n10594 vdd.n10552 23.783
R41975 vdd.n10594 vdd.n10558 23.783
R41976 vdd.n10595 vdd.n10544 23.783
R41977 vdd.n10595 vdd.n10550 23.783
R41978 vdd.n10596 vdd.n10536 23.783
R41979 vdd.n10596 vdd.n10542 23.783
R41980 vdd.n10597 vdd.n10528 23.783
R41981 vdd.n10597 vdd.n10534 23.783
R41982 vdd.n10598 vdd.n10520 23.783
R41983 vdd.n10598 vdd.n10526 23.783
R41984 vdd.n10599 vdd.n10512 23.783
R41985 vdd.n10599 vdd.n10518 23.783
R41986 vdd.n10600 vdd.n10504 23.783
R41987 vdd.n10600 vdd.n10508 23.783
R41988 vdd.n10601 vdd.n10496 23.783
R41989 vdd.n10601 vdd.n10502 23.783
R41990 vdd.n10602 vdd.n10488 23.783
R41991 vdd.n10602 vdd.n10494 23.783
R41992 vdd.n10603 vdd.n10480 23.783
R41993 vdd.n10603 vdd.n10486 23.783
R41994 vdd.n10604 vdd.n10472 23.783
R41995 vdd.n10604 vdd.n10478 23.783
R41996 vdd.n10605 vdd.n10464 23.783
R41997 vdd.n10605 vdd.n10470 23.783
R41998 vdd.n10606 vdd.n10456 23.783
R41999 vdd.n10606 vdd.n10462 23.783
R42000 vdd.n10607 vdd.n10448 23.783
R42001 vdd.n10607 vdd.n10454 23.783
R42002 vdd.n10608 vdd.n10440 23.783
R42003 vdd.n10608 vdd.n10446 23.783
R42004 vdd.n10619 vdd.n10618 23.783
R42005 vdd.n10619 vdd.n10613 23.783
R42006 vdd.n10770 vdd.n10769 23.783
R42007 vdd.n10770 vdd.n10767 23.783
R42008 vdd.n10771 vdd.n10756 23.783
R42009 vdd.n10771 vdd.n10762 23.783
R42010 vdd.n10772 vdd.n10748 23.783
R42011 vdd.n10772 vdd.n10754 23.783
R42012 vdd.n10773 vdd.n10740 23.783
R42013 vdd.n10773 vdd.n10746 23.783
R42014 vdd.n10774 vdd.n10732 23.783
R42015 vdd.n10774 vdd.n10738 23.783
R42016 vdd.n10775 vdd.n10724 23.783
R42017 vdd.n10775 vdd.n10730 23.783
R42018 vdd.n10776 vdd.n10716 23.783
R42019 vdd.n10776 vdd.n10722 23.783
R42020 vdd.n10777 vdd.n10708 23.783
R42021 vdd.n10777 vdd.n10714 23.783
R42022 vdd.n10778 vdd.n10700 23.783
R42023 vdd.n10778 vdd.n10706 23.783
R42024 vdd.n10779 vdd.n10692 23.783
R42025 vdd.n10779 vdd.n10698 23.783
R42026 vdd.n10780 vdd.n10684 23.783
R42027 vdd.n10780 vdd.n10688 23.783
R42028 vdd.n10781 vdd.n10676 23.783
R42029 vdd.n10781 vdd.n10682 23.783
R42030 vdd.n10782 vdd.n10668 23.783
R42031 vdd.n10782 vdd.n10674 23.783
R42032 vdd.n10783 vdd.n10660 23.783
R42033 vdd.n10783 vdd.n10666 23.783
R42034 vdd.n10784 vdd.n10652 23.783
R42035 vdd.n10784 vdd.n10658 23.783
R42036 vdd.n10785 vdd.n10644 23.783
R42037 vdd.n10785 vdd.n10650 23.783
R42038 vdd.n10786 vdd.n10636 23.783
R42039 vdd.n10786 vdd.n10642 23.783
R42040 vdd.n10787 vdd.n10628 23.783
R42041 vdd.n10787 vdd.n10634 23.783
R42042 vdd.n10788 vdd.n10620 23.783
R42043 vdd.n10788 vdd.n10626 23.783
R42044 vdd.n10799 vdd.n10798 23.783
R42045 vdd.n10799 vdd.n10793 23.783
R42046 vdd.n10950 vdd.n10949 23.783
R42047 vdd.n10950 vdd.n10947 23.783
R42048 vdd.n10951 vdd.n10936 23.783
R42049 vdd.n10951 vdd.n10942 23.783
R42050 vdd.n10952 vdd.n10928 23.783
R42051 vdd.n10952 vdd.n10934 23.783
R42052 vdd.n10953 vdd.n10920 23.783
R42053 vdd.n10953 vdd.n10926 23.783
R42054 vdd.n10954 vdd.n10912 23.783
R42055 vdd.n10954 vdd.n10918 23.783
R42056 vdd.n10955 vdd.n10904 23.783
R42057 vdd.n10955 vdd.n10910 23.783
R42058 vdd.n10956 vdd.n10896 23.783
R42059 vdd.n10956 vdd.n10902 23.783
R42060 vdd.n10957 vdd.n10888 23.783
R42061 vdd.n10957 vdd.n10894 23.783
R42062 vdd.n10958 vdd.n10880 23.783
R42063 vdd.n10958 vdd.n10886 23.783
R42064 vdd.n10959 vdd.n10872 23.783
R42065 vdd.n10959 vdd.n10878 23.783
R42066 vdd.n10960 vdd.n10864 23.783
R42067 vdd.n10960 vdd.n10868 23.783
R42068 vdd.n10961 vdd.n10856 23.783
R42069 vdd.n10961 vdd.n10862 23.783
R42070 vdd.n10962 vdd.n10848 23.783
R42071 vdd.n10962 vdd.n10854 23.783
R42072 vdd.n10963 vdd.n10840 23.783
R42073 vdd.n10963 vdd.n10846 23.783
R42074 vdd.n10964 vdd.n10832 23.783
R42075 vdd.n10964 vdd.n10838 23.783
R42076 vdd.n10965 vdd.n10824 23.783
R42077 vdd.n10965 vdd.n10830 23.783
R42078 vdd.n10966 vdd.n10816 23.783
R42079 vdd.n10966 vdd.n10822 23.783
R42080 vdd.n10967 vdd.n10808 23.783
R42081 vdd.n10967 vdd.n10814 23.783
R42082 vdd.n10968 vdd.n10800 23.783
R42083 vdd.n10968 vdd.n10806 23.783
R42084 vdd.n10979 vdd.n10978 23.783
R42085 vdd.n10979 vdd.n10973 23.783
R42086 vdd.n11130 vdd.n11129 23.783
R42087 vdd.n11130 vdd.n11127 23.783
R42088 vdd.n11131 vdd.n11116 23.783
R42089 vdd.n11131 vdd.n11122 23.783
R42090 vdd.n11132 vdd.n11108 23.783
R42091 vdd.n11132 vdd.n11114 23.783
R42092 vdd.n11133 vdd.n11100 23.783
R42093 vdd.n11133 vdd.n11106 23.783
R42094 vdd.n11134 vdd.n11092 23.783
R42095 vdd.n11134 vdd.n11098 23.783
R42096 vdd.n11135 vdd.n11084 23.783
R42097 vdd.n11135 vdd.n11090 23.783
R42098 vdd.n11136 vdd.n11076 23.783
R42099 vdd.n11136 vdd.n11082 23.783
R42100 vdd.n11137 vdd.n11068 23.783
R42101 vdd.n11137 vdd.n11074 23.783
R42102 vdd.n11138 vdd.n11060 23.783
R42103 vdd.n11138 vdd.n11066 23.783
R42104 vdd.n11139 vdd.n11052 23.783
R42105 vdd.n11139 vdd.n11058 23.783
R42106 vdd.n11140 vdd.n11044 23.783
R42107 vdd.n11140 vdd.n11048 23.783
R42108 vdd.n11141 vdd.n11036 23.783
R42109 vdd.n11141 vdd.n11042 23.783
R42110 vdd.n11142 vdd.n11028 23.783
R42111 vdd.n11142 vdd.n11034 23.783
R42112 vdd.n11143 vdd.n11020 23.783
R42113 vdd.n11143 vdd.n11026 23.783
R42114 vdd.n11144 vdd.n11012 23.783
R42115 vdd.n11144 vdd.n11018 23.783
R42116 vdd.n11145 vdd.n11004 23.783
R42117 vdd.n11145 vdd.n11010 23.783
R42118 vdd.n11146 vdd.n10996 23.783
R42119 vdd.n11146 vdd.n11002 23.783
R42120 vdd.n11147 vdd.n10988 23.783
R42121 vdd.n11147 vdd.n10994 23.783
R42122 vdd.n11148 vdd.n10980 23.783
R42123 vdd.n11148 vdd.n10986 23.783
R42124 vdd.n11159 vdd.n11158 23.783
R42125 vdd.n11159 vdd.n11153 23.783
R42126 vdd.n11310 vdd.n11309 23.783
R42127 vdd.n11310 vdd.n11307 23.783
R42128 vdd.n11311 vdd.n11296 23.783
R42129 vdd.n11311 vdd.n11302 23.783
R42130 vdd.n11312 vdd.n11288 23.783
R42131 vdd.n11312 vdd.n11294 23.783
R42132 vdd.n11313 vdd.n11280 23.783
R42133 vdd.n11313 vdd.n11286 23.783
R42134 vdd.n11314 vdd.n11272 23.783
R42135 vdd.n11314 vdd.n11278 23.783
R42136 vdd.n11315 vdd.n11264 23.783
R42137 vdd.n11315 vdd.n11270 23.783
R42138 vdd.n11316 vdd.n11256 23.783
R42139 vdd.n11316 vdd.n11262 23.783
R42140 vdd.n11317 vdd.n11248 23.783
R42141 vdd.n11317 vdd.n11254 23.783
R42142 vdd.n11318 vdd.n11240 23.783
R42143 vdd.n11318 vdd.n11246 23.783
R42144 vdd.n11319 vdd.n11232 23.783
R42145 vdd.n11319 vdd.n11238 23.783
R42146 vdd.n11320 vdd.n11224 23.783
R42147 vdd.n11320 vdd.n11228 23.783
R42148 vdd.n11321 vdd.n11216 23.783
R42149 vdd.n11321 vdd.n11222 23.783
R42150 vdd.n11322 vdd.n11208 23.783
R42151 vdd.n11322 vdd.n11214 23.783
R42152 vdd.n11323 vdd.n11200 23.783
R42153 vdd.n11323 vdd.n11206 23.783
R42154 vdd.n11324 vdd.n11192 23.783
R42155 vdd.n11324 vdd.n11198 23.783
R42156 vdd.n11325 vdd.n11184 23.783
R42157 vdd.n11325 vdd.n11190 23.783
R42158 vdd.n11326 vdd.n11176 23.783
R42159 vdd.n11326 vdd.n11182 23.783
R42160 vdd.n11327 vdd.n11168 23.783
R42161 vdd.n11327 vdd.n11174 23.783
R42162 vdd.n11328 vdd.n11160 23.783
R42163 vdd.n11328 vdd.n11166 23.783
R42164 vdd.n11339 vdd.n11338 23.783
R42165 vdd.n11339 vdd.n11333 23.783
R42166 vdd.n13481 vdd.t1083 7.146
R42167 vdd.n13478 vdd.t677 7.146
R42168 vdd.n13534 vdd.t2430 7.146
R42169 vdd.n13530 vdd.t2697 7.146
R42170 vdd.n13527 vdd.t884 7.146
R42171 vdd.n13524 vdd.t1123 7.146
R42172 vdd.n13521 vdd.t2269 7.146
R42173 vdd.n13518 vdd.t2695 7.146
R42174 vdd.n13515 vdd.t2926 7.146
R42175 vdd.n13512 vdd.t1060 7.146
R42176 vdd.n13509 vdd.t603 7.146
R42177 vdd.n13506 vdd.t1723 7.146
R42178 vdd.n13505 vdd.t2135 7.146
R42179 vdd.n13502 vdd.t2997 7.146
R42180 vdd.n13499 vdd.t1030 7.146
R42181 vdd.n13496 vdd.t1253 7.146
R42182 vdd.n13493 vdd.t138 7.146
R42183 vdd.n13490 vdd.t1980 7.146
R42184 vdd.n13487 vdd.t2455 7.146
R42185 vdd.n13484 vdd.t1315 7.146
R42186 vdd.n13458 vdd.t510 7.146
R42187 vdd.n13458 vdd.t2634 7.146
R42188 vdd.n13447 vdd.t762 7.146
R42189 vdd.n13447 vdd.t2880 7.146
R42190 vdd.n13446 vdd.t2976 7.146
R42191 vdd.n13446 vdd.t313 7.146
R42192 vdd.n13445 vdd.t247 7.146
R42193 vdd.n13445 vdd.t560 7.146
R42194 vdd.n13444 vdd.t1362 7.146
R42195 vdd.n13444 vdd.t1675 7.146
R42196 vdd.n13443 vdd.t1774 7.146
R42197 vdd.n13443 vdd.t2100 7.146
R42198 vdd.n13442 vdd.t2028 7.146
R42199 vdd.n13442 vdd.t2329 7.146
R42200 vdd.n13441 vdd.t174 7.146
R42201 vdd.n13441 vdd.t481 7.146
R42202 vdd.n13440 vdd.t2689 7.146
R42203 vdd.n13440 vdd.t2999 7.146
R42204 vdd.n13439 vdd.t824 7.146
R42205 vdd.n13439 vdd.t1129 7.146
R42206 vdd.n13438 vdd.t1228 7.146
R42207 vdd.n13438 vdd.t1551 7.146
R42208 vdd.n13437 vdd.t1467 7.146
R42209 vdd.n13437 vdd.t746 7.146
R42210 vdd.n13436 vdd.t150 7.146
R42211 vdd.n13436 vdd.t464 7.146
R42212 vdd.n13435 vdd.t2311 7.146
R42213 vdd.n13435 vdd.t1438 7.146
R42214 vdd.n13434 vdd.t1173 7.146
R42215 vdd.n13434 vdd.t323 7.146
R42216 vdd.n13433 vdd.t48 7.146
R42217 vdd.n13433 vdd.t2180 7.146
R42218 vdd.n13432 vdd.t526 7.146
R42219 vdd.n13432 vdd.t2653 7.146
R42220 vdd.n13431 vdd.t2372 7.146
R42221 vdd.n13431 vdd.t1507 7.146
R42222 vdd.n13430 vdd.t2137 7.146
R42223 vdd.n13430 vdd.t1265 7.146
R42224 vdd.n13429 vdd.t1724 7.146
R42225 vdd.n13429 vdd.t855 7.146
R42226 vdd.n13278 vdd.t2305 7.146
R42227 vdd.n13278 vdd.t2117 7.146
R42228 vdd.n13267 vdd.t2557 7.146
R42229 vdd.n13267 vdd.t2358 7.146
R42230 vdd.n13266 vdd.t1280 7.146
R42231 vdd.n13266 vdd.t1877 7.146
R42232 vdd.n13265 vdd.t1537 7.146
R42233 vdd.n13265 vdd.t2120 7.146
R42234 vdd.n13264 vdd.t2687 7.146
R42235 vdd.n13264 vdd.t281 7.146
R42236 vdd.n13263 vdd.t108 7.146
R42237 vdd.n13263 vdd.t694 7.146
R42238 vdd.n13262 vdd.t348 7.146
R42239 vdd.n13262 vdd.t913 7.146
R42240 vdd.n13261 vdd.t1461 7.146
R42241 vdd.n13261 vdd.t2067 7.146
R42242 vdd.n13260 vdd.t983 7.146
R42243 vdd.n13260 vdd.t1580 7.146
R42244 vdd.n13259 vdd.t2126 7.146
R42245 vdd.n13259 vdd.t2734 7.146
R42246 vdd.n13258 vdd.t2550 7.146
R42247 vdd.n13258 vdd.t155 7.146
R42248 vdd.n13257 vdd.t95 7.146
R42249 vdd.n13257 vdd.t2341 7.146
R42250 vdd.n13256 vdd.t1437 7.146
R42251 vdd.n13256 vdd.t2042 7.146
R42252 vdd.n13255 vdd.t1122 7.146
R42253 vdd.n13255 vdd.t929 7.146
R42254 vdd.n13254 vdd.t2992 7.146
R42255 vdd.n13254 vdd.t2797 7.146
R42256 vdd.n13253 vdd.t1846 7.146
R42257 vdd.n13253 vdd.t1656 7.146
R42258 vdd.n13252 vdd.t2320 7.146
R42259 vdd.n13252 vdd.t2140 7.146
R42260 vdd.n13251 vdd.t1188 7.146
R42261 vdd.n13251 vdd.t994 7.146
R42262 vdd.n13250 vdd.t941 7.146
R42263 vdd.n13250 vdd.t780 7.146
R42264 vdd.n13249 vdd.t550 7.146
R42265 vdd.n13249 vdd.t357 7.146
R42266 vdd.n13098 vdd.t2139 7.146
R42267 vdd.n13098 vdd.t924 7.146
R42268 vdd.n13087 vdd.t2376 7.146
R42269 vdd.n13087 vdd.t1171 7.146
R42270 vdd.n13086 vdd.t1851 7.146
R42271 vdd.n13086 vdd.t213 7.146
R42272 vdd.n13085 vdd.t2104 7.146
R42273 vdd.n13085 vdd.t457 7.146
R42274 vdd.n13084 vdd.t261 7.146
R42275 vdd.n13084 vdd.t1575 7.146
R42276 vdd.n13083 vdd.t662 7.146
R42277 vdd.n13083 vdd.t1994 7.146
R42278 vdd.n13082 vdd.t896 7.146
R42279 vdd.n13082 vdd.t2246 7.146
R42280 vdd.n13081 vdd.t2047 7.146
R42281 vdd.n13081 vdd.t393 7.146
R42282 vdd.n13080 vdd.t1560 7.146
R42283 vdd.n13080 vdd.t2904 7.146
R42284 vdd.n13079 vdd.t2713 7.146
R42285 vdd.n13079 vdd.t1023 7.146
R42286 vdd.n13078 vdd.t127 7.146
R42287 vdd.n13078 vdd.t1440 7.146
R42288 vdd.n13077 vdd.t2449 7.146
R42289 vdd.n13077 vdd.t938 7.146
R42290 vdd.n13076 vdd.t2013 7.146
R42291 vdd.n13076 vdd.t360 7.146
R42292 vdd.n13075 vdd.t947 7.146
R42293 vdd.n13075 vdd.t2761 7.146
R42294 vdd.n13074 vdd.t2819 7.146
R42295 vdd.n13074 vdd.t1605 7.146
R42296 vdd.n13073 vdd.t1679 7.146
R42297 vdd.n13073 vdd.t480 7.146
R42298 vdd.n13072 vdd.t2161 7.146
R42299 vdd.n13072 vdd.t943 7.146
R42300 vdd.n13071 vdd.t1016 7.146
R42301 vdd.n13071 vdd.t2816 7.146
R42302 vdd.n13070 vdd.t797 7.146
R42303 vdd.n13070 vdd.t2586 7.146
R42304 vdd.n13069 vdd.t383 7.146
R42305 vdd.n13069 vdd.t2157 7.146
R42306 vdd.n12918 vdd.t942 7.146
R42307 vdd.n12918 vdd.t1993 7.146
R42308 vdd.n12907 vdd.t1192 7.146
R42309 vdd.n12907 vdd.t2245 7.146
R42310 vdd.n12906 vdd.t191 7.146
R42311 vdd.n12906 vdd.t2288 7.146
R42312 vdd.n12905 vdd.t435 7.146
R42313 vdd.n12905 vdd.t2532 7.146
R42314 vdd.n12904 vdd.t1555 7.146
R42315 vdd.n12904 vdd.t685 7.146
R42316 vdd.n12903 vdd.t1964 7.146
R42317 vdd.n12903 vdd.t1091 7.146
R42318 vdd.n12902 vdd.t2224 7.146
R42319 vdd.n12902 vdd.t1322 7.146
R42320 vdd.n12901 vdd.t367 7.146
R42321 vdd.n12901 vdd.t2461 7.146
R42322 vdd.n12900 vdd.t2879 7.146
R42323 vdd.n12900 vdd.t1987 7.146
R42324 vdd.n12899 vdd.t998 7.146
R42325 vdd.n12899 vdd.t147 7.146
R42326 vdd.n12898 vdd.t1420 7.146
R42327 vdd.n12898 vdd.t556 7.146
R42328 vdd.n12897 vdd.t1054 7.146
R42329 vdd.n12897 vdd.t2420 7.146
R42330 vdd.n12896 vdd.t337 7.146
R42331 vdd.n12896 vdd.t2433 7.146
R42332 vdd.n12895 vdd.t2774 7.146
R42333 vdd.n12895 vdd.t817 7.146
R42334 vdd.n12894 vdd.t1630 7.146
R42335 vdd.n12894 vdd.t2682 7.146
R42336 vdd.n12893 vdd.t505 7.146
R42337 vdd.n12893 vdd.t1530 7.146
R42338 vdd.n12892 vdd.t959 7.146
R42339 vdd.n12892 vdd.t2019 7.146
R42340 vdd.n12891 vdd.t2836 7.146
R42341 vdd.n12891 vdd.t876 7.146
R42342 vdd.n12890 vdd.t2603 7.146
R42343 vdd.n12890 vdd.t639 7.146
R42344 vdd.n12889 vdd.t2184 7.146
R42345 vdd.n12889 vdd.t239 7.146
R42346 vdd.n12738 vdd.t2414 7.146
R42347 vdd.n12738 vdd.t1814 7.146
R42348 vdd.n12727 vdd.t2681 7.146
R42349 vdd.n12727 vdd.t2074 7.146
R42350 vdd.n12726 vdd.t2498 7.146
R42351 vdd.n12726 vdd.t2856 7.146
R42352 vdd.n12725 vdd.t2760 7.146
R42353 vdd.n12725 vdd.t114 7.146
R42354 vdd.n12724 vdd.t885 7.146
R42355 vdd.n12724 vdd.t1232 7.146
R42356 vdd.n12723 vdd.t1288 7.146
R42357 vdd.n12723 vdd.t1642 7.146
R42358 vdd.n12722 vdd.t1548 7.146
R42359 vdd.n12722 vdd.t1895 7.146
R42360 vdd.n12721 vdd.t2701 7.146
R42361 vdd.n12721 vdd.t35 7.146
R42362 vdd.n12720 vdd.t2217 7.146
R42363 vdd.n12720 vdd.t2554 7.146
R42364 vdd.n12719 vdd.t356 7.146
R42365 vdd.n12719 vdd.t708 7.146
R42366 vdd.n12718 vdd.t778 7.146
R42367 vdd.n12718 vdd.t1104 7.146
R42368 vdd.n12717 vdd.t1903 7.146
R42369 vdd.n12717 vdd.t1796 7.146
R42370 vdd.n12716 vdd.t2661 7.146
R42371 vdd.n12716 vdd.t5 7.146
R42372 vdd.n12715 vdd.t1244 7.146
R42373 vdd.n12715 vdd.t646 7.146
R42374 vdd.n12714 vdd.t123 7.146
R42375 vdd.n12714 vdd.t2494 7.146
R42376 vdd.n12713 vdd.t1960 7.146
R42377 vdd.n12713 vdd.t1365 7.146
R42378 vdd.n12712 vdd.t2439 7.146
R42379 vdd.n12712 vdd.t1831 7.146
R42380 vdd.n12711 vdd.t1301 7.146
R42381 vdd.n12711 vdd.t727 7.146
R42382 vdd.n12710 vdd.t1071 7.146
R42383 vdd.n12710 vdd.t471 7.146
R42384 vdd.n12709 vdd.t659 7.146
R42385 vdd.n12709 vdd.t53 7.146
R42386 vdd.n12558 vdd.t1498 7.146
R42387 vdd.n12558 vdd.t641 7.146
R42388 vdd.n12547 vdd.t1748 7.146
R42389 vdd.n12547 vdd.t875 7.146
R42390 vdd.n12546 vdd.t847 7.146
R42391 vdd.n12546 vdd.t1158 7.146
R42392 vdd.n12545 vdd.t1097 7.146
R42393 vdd.n12545 vdd.t1405 7.146
R42394 vdd.n12544 vdd.t2240 7.146
R42395 vdd.n12544 vdd.t2551 7.146
R42396 vdd.n12543 vdd.t2648 7.146
R42397 vdd.n12543 vdd.t2964 7.146
R42398 vdd.n12542 vdd.t2899 7.146
R42399 vdd.n12542 vdd.t227 7.146
R42400 vdd.n12541 vdd.t1015 7.146
R42401 vdd.n12541 vdd.t1338 7.146
R42402 vdd.n12540 vdd.t565 7.146
R42403 vdd.n12540 vdd.t869 7.146
R42404 vdd.n12539 vdd.t1678 7.146
R42405 vdd.n12539 vdd.t2008 7.146
R42406 vdd.n12538 vdd.t2103 7.146
R42407 vdd.n12538 vdd.t2411 7.146
R42408 vdd.n12537 vdd.t1145 7.146
R42409 vdd.n12537 vdd.t425 7.146
R42410 vdd.n12536 vdd.t987 7.146
R42411 vdd.n12536 vdd.t1312 7.146
R42412 vdd.n12535 vdd.t331 7.146
R42413 vdd.n12535 vdd.t2444 7.146
R42414 vdd.n12534 vdd.t2190 7.146
R42415 vdd.n12534 vdd.t1306 7.146
R42416 vdd.n12533 vdd.t1045 7.146
R42417 vdd.n12533 vdd.t193 7.146
R42418 vdd.n12532 vdd.t1516 7.146
R42419 vdd.n12532 vdd.t661 7.146
R42420 vdd.n12531 vdd.t407 7.146
R42421 vdd.n12531 vdd.t2510 7.146
R42422 vdd.n12530 vdd.t165 7.146
R42423 vdd.n12530 vdd.t2277 7.146
R42424 vdd.n12529 vdd.t2740 7.146
R42425 vdd.n12529 vdd.t1850 7.146
R42426 vdd.n12378 vdd.t326 7.146
R42427 vdd.n12378 vdd.t2438 7.146
R42428 vdd.n12367 vdd.t577 7.146
R42429 vdd.n12367 vdd.t2706 7.146
R42430 vdd.n12366 vdd.t2163 7.146
R42431 vdd.n12366 vdd.t2475 7.146
R42432 vdd.n12365 vdd.t2398 7.146
R42433 vdd.n12365 vdd.t2742 7.146
R42434 vdd.n12364 vdd.t559 7.146
R42435 vdd.n12364 vdd.t862 7.146
R42436 vdd.n12363 vdd.t950 7.146
R42437 vdd.n12363 vdd.t1271 7.146
R42438 vdd.n12362 vdd.t1200 7.146
R42439 vdd.n12362 vdd.t1519 7.146
R42440 vdd.n12361 vdd.t2328 7.146
R42441 vdd.n12361 vdd.t2667 7.146
R42442 vdd.n12360 vdd.t1859 7.146
R42443 vdd.n12360 vdd.t2193 7.146
R42444 vdd.n12359 vdd.t1 7.146
R42445 vdd.n12359 vdd.t333 7.146
R42446 vdd.n12358 vdd.t434 7.146
R42447 vdd.n12358 vdd.t758 7.146
R42448 vdd.n12357 vdd.t2765 7.146
R42449 vdd.n12357 vdd.t2007 7.146
R42450 vdd.n12356 vdd.t2310 7.146
R42451 vdd.n12356 vdd.t2639 7.146
R42452 vdd.n12355 vdd.t2129 7.146
R42453 vdd.n12355 vdd.t1260 7.146
R42454 vdd.n12354 vdd.t982 7.146
R42455 vdd.n12354 vdd.t146 7.146
R42456 vdd.n12353 vdd.t2862 7.146
R42457 vdd.n12353 vdd.t1986 7.146
R42458 vdd.n12352 vdd.t347 7.146
R42459 vdd.n12352 vdd.t2460 7.146
R42460 vdd.n12351 vdd.t2207 7.146
R42461 vdd.n12351 vdd.t1321 7.146
R42462 vdd.n12350 vdd.t1950 7.146
R42463 vdd.n12350 vdd.t1090 7.146
R42464 vdd.n12349 vdd.t1536 7.146
R42465 vdd.n12349 vdd.t684 7.146
R42466 vdd.n12198 vdd.t2123 7.146
R42467 vdd.n12198 vdd.t2278 7.146
R42468 vdd.n12187 vdd.t2365 7.146
R42469 vdd.n12187 vdd.t2512 7.146
R42470 vdd.n12186 vdd.t484 7.146
R42471 vdd.n12186 vdd.t57 7.146
R42472 vdd.n12185 vdd.t745 7.146
R42473 vdd.n12185 vdd.t307 7.146
R42474 vdd.n12184 vdd.t1853 7.146
R42475 vdd.n12184 vdd.t1422 7.146
R42476 vdd.n12183 vdd.t2280 7.146
R42477 vdd.n12183 vdd.t1833 7.146
R42478 vdd.n12182 vdd.t2514 7.146
R42479 vdd.n12182 vdd.t2096 7.146
R42480 vdd.n12181 vdd.t665 7.146
R42481 vdd.n12181 vdd.t249 7.146
R42482 vdd.n12180 vdd.t198 7.146
R42483 vdd.n12180 vdd.t2756 7.146
R42484 vdd.n12179 vdd.t1308 7.146
R42485 vdd.n12179 vdd.t881 7.146
R42486 vdd.n12178 vdd.t1733 7.146
R42487 vdd.n12178 vdd.t1282 7.146
R42488 vdd.n12177 vdd.t1355 7.146
R42489 vdd.n12177 vdd.t1380 7.146
R42490 vdd.n12176 vdd.t638 7.146
R42491 vdd.n12176 vdd.t217 7.146
R42492 vdd.n12175 vdd.t932 7.146
R42493 vdd.n12175 vdd.t1096 7.146
R42494 vdd.n12174 vdd.t2803 7.146
R42495 vdd.n12174 vdd.t2958 7.146
R42496 vdd.n12173 vdd.t1664 7.146
R42497 vdd.n12173 vdd.t1811 7.146
R42498 vdd.n12172 vdd.t2148 7.146
R42499 vdd.n12172 vdd.t2295 7.146
R42500 vdd.n12171 vdd.t1002 7.146
R42501 vdd.n12171 vdd.t1149 7.146
R42502 vdd.n12170 vdd.t789 7.146
R42503 vdd.n12170 vdd.t909 7.146
R42504 vdd.n12169 vdd.t366 7.146
R42505 vdd.n12169 vdd.t509 7.146
R42506 vdd.n12018 vdd.t689 7.146
R42507 vdd.n12018 vdd.t2996 7.146
R42508 vdd.n12007 vdd.t908 7.146
R42509 vdd.n12007 vdd.t262 7.146
R42510 vdd.n12006 vdd.t1384 7.146
R42511 vdd.n12006 vdd.t177 7.146
R42512 vdd.n12005 vdd.t1623 7.146
R42513 vdd.n12005 vdd.t423 7.146
R42514 vdd.n12004 vdd.t2771 7.146
R42515 vdd.n12004 vdd.t1535 7.146
R42516 vdd.n12003 vdd.t195 7.146
R42517 vdd.n12003 vdd.t1949 7.146
R42518 vdd.n12002 vdd.t440 7.146
R42519 vdd.n12002 vdd.t2206 7.146
R42520 vdd.n12001 vdd.t1559 7.146
R42521 vdd.n12001 vdd.t349 7.146
R42522 vdd.n12000 vdd.t1085 7.146
R42523 vdd.n12000 vdd.t2861 7.146
R42524 vdd.n11999 vdd.t2230 7.146
R42525 vdd.n11999 vdd.t981 7.146
R42526 vdd.n11998 vdd.t2637 7.146
R42527 vdd.n11998 vdd.t1404 7.146
R42528 vdd.n11997 vdd.t2728 7.146
R42529 vdd.n11997 vdd.t2108 7.146
R42530 vdd.n11996 vdd.t1528 7.146
R42531 vdd.n11996 vdd.t325 7.146
R42532 vdd.n11995 vdd.t2482 7.146
R42533 vdd.n11995 vdd.t1803 7.146
R42534 vdd.n11994 vdd.t1351 7.146
R42535 vdd.n11994 vdd.t693 7.146
R42536 vdd.n11993 vdd.t238 7.146
R42537 vdd.n11993 vdd.t2539 7.146
R42538 vdd.n11992 vdd.t714 7.146
R42539 vdd.n11992 vdd.t20 7.146
R42540 vdd.n11991 vdd.t2566 7.146
R42541 vdd.n11991 vdd.t1876 7.146
R42542 vdd.n11990 vdd.t2308 7.146
R42543 vdd.n11990 vdd.t1632 7.146
R42544 vdd.n11989 vdd.t1900 7.146
R42545 vdd.n11989 vdd.t1216 7.146
R42546 vdd.n11838 vdd.t2474 7.146
R42547 vdd.n11838 vdd.t536 7.146
R42548 vdd.n11827 vdd.t2741 7.146
R42549 vdd.n11827 vdd.t793 7.146
R42550 vdd.n11826 vdd.t2714 7.146
R42551 vdd.n11826 vdd.t1805 7.146
R42552 vdd.n11825 vdd.t2940 7.146
R42553 vdd.n11825 vdd.t2066 7.146
R42554 vdd.n11824 vdd.t1080 7.146
R42555 vdd.n11824 vdd.t211 7.146
R42556 vdd.n11823 vdd.t1484 7.146
R42557 vdd.n11823 vdd.t620 7.146
R42558 vdd.n11822 vdd.t1742 7.146
R42559 vdd.n11822 vdd.t854 7.146
R42560 vdd.n11821 vdd.t2884 7.146
R42561 vdd.n11821 vdd.t1985 7.146
R42562 vdd.n11820 vdd.t2389 7.146
R42563 vdd.n11820 vdd.t1506 7.146
R42564 vdd.n11819 vdd.t548 7.146
R42565 vdd.n11819 vdd.t2652 7.146
R42566 vdd.n11818 vdd.t940 7.146
R42567 vdd.n11818 vdd.t76 7.146
R42568 vdd.n11817 vdd.t1305 7.146
R42569 vdd.n11817 vdd.t2705 7.146
R42570 vdd.n11816 vdd.t2851 7.146
R42571 vdd.n11816 vdd.t1956 7.146
R42572 vdd.n11815 vdd.t1287 7.146
R42573 vdd.n11815 vdd.t2332 7.146
R42574 vdd.n11814 vdd.t184 7.146
R42575 vdd.n11814 vdd.t1202 7.146
R42576 vdd.n11813 vdd.t2039 7.146
R42577 vdd.n11813 vdd.t80 7.146
R42578 vdd.n11812 vdd.t2497 7.146
R42579 vdd.n11812 vdd.t563 7.146
R42580 vdd.n11811 vdd.t1371 7.146
R42581 vdd.n11811 vdd.t2401 7.146
R42582 vdd.n11810 vdd.t1119 7.146
R42583 vdd.n11810 vdd.t2165 7.146
R42584 vdd.n11809 vdd.t730 7.146
R42585 vdd.n11809 vdd.t1752 7.146
R42586 vdd.n11658 vdd.t558 7.146
R42587 vdd.n11658 vdd.t370 7.146
R42588 vdd.n11647 vdd.t803 7.146
R42589 vdd.n11647 vdd.t614 7.146
R42590 vdd.n11646 vdd.t1787 7.146
R42591 vdd.n11646 vdd.t2368 7.146
R42592 vdd.n11645 vdd.t2046 7.146
R42593 vdd.n11645 vdd.t2620 7.146
R42594 vdd.n11644 vdd.t189 7.146
R42595 vdd.n11644 vdd.t776 7.146
R42596 vdd.n11643 vdd.t606 7.146
R42597 vdd.n11643 vdd.t1164 7.146
R42598 vdd.n11642 vdd.t835 7.146
R42599 vdd.n11642 vdd.t1408 7.146
R42600 vdd.n11641 vdd.t1958 7.146
R42601 vdd.n11641 vdd.t2553 7.146
R42602 vdd.n11640 vdd.t1481 7.146
R42603 vdd.n11640 vdd.t2085 7.146
R42604 vdd.n11639 vdd.t2629 7.146
R42605 vdd.n11639 vdd.t231 7.146
R42606 vdd.n11638 vdd.t49 7.146
R42607 vdd.n11638 vdd.t634 7.146
R42608 vdd.n11637 vdd.t2790 7.146
R42609 vdd.n11637 vdd.t2077 7.146
R42610 vdd.n11636 vdd.t1941 7.146
R42611 vdd.n11636 vdd.t2524 7.146
R42612 vdd.n11635 vdd.t2355 7.146
R42613 vdd.n11635 vdd.t2176 7.146
R42614 vdd.n11634 vdd.t1222 7.146
R42615 vdd.n11634 vdd.t1027 7.146
R42616 vdd.n11633 vdd.t105 7.146
R42617 vdd.n11633 vdd.t2909 7.146
R42618 vdd.n11632 vdd.t583 7.146
R42619 vdd.n11632 vdd.t395 7.146
R42620 vdd.n11631 vdd.t2419 7.146
R42621 vdd.n11631 vdd.t2249 7.146
R42622 vdd.n11630 vdd.t2192 7.146
R42623 vdd.n11630 vdd.t1995 7.146
R42624 vdd.n11629 vdd.t1770 7.146
R42625 vdd.n11629 vdd.t1577 7.146
R42626 vdd.n179 vdd.t41 7.146
R42627 vdd.n179 vdd.t2164 7.146
R42628 vdd.n168 vdd.t298 7.146
R42629 vdd.n168 vdd.t2402 7.146
R42630 vdd.n167 vdd.t391 7.146
R42631 vdd.n167 vdd.t711 7.146
R42632 vdd.n166 vdd.t623 7.146
R42633 vdd.n166 vdd.t928 7.146
R42634 vdd.n165 vdd.t1754 7.146
R42635 vdd.n165 vdd.t2084 7.146
R42636 vdd.n164 vdd.t2169 7.146
R42637 vdd.n164 vdd.t2481 7.146
R42638 vdd.n163 vdd.t2403 7.146
R42639 vdd.n163 vdd.t2746 7.146
R42640 vdd.n162 vdd.t567 7.146
R42641 vdd.n162 vdd.t868 7.146
R42642 vdd.n161 vdd.t82 7.146
R42643 vdd.n161 vdd.t412 7.146
R42644 vdd.n160 vdd.t1204 7.146
R42645 vdd.n160 vdd.t1523 7.146
R42646 vdd.n159 vdd.t1619 7.146
R42647 vdd.n159 vdd.t1942 7.146
R42648 vdd.n158 vdd.t1411 7.146
R42649 vdd.n158 vdd.t676 7.146
R42650 vdd.n157 vdd.t533 7.146
R42651 vdd.n157 vdd.t844 7.146
R42652 vdd.n156 vdd.t1842 7.146
R42653 vdd.n156 vdd.t969 7.146
R42654 vdd.n155 vdd.t736 7.146
R42655 vdd.n155 vdd.t2847 7.146
R42656 vdd.n154 vdd.t2591 7.146
R42657 vdd.n154 vdd.t1709 7.146
R42658 vdd.n153 vdd.t68 7.146
R42659 vdd.n153 vdd.t2196 7.146
R42660 vdd.n152 vdd.t1921 7.146
R42661 vdd.n152 vdd.t1052 7.146
R42662 vdd.n151 vdd.t1670 7.146
R42663 vdd.n151 vdd.t815 7.146
R42664 vdd.n150 vdd.t1256 7.146
R42665 vdd.n150 vdd.t411 7.146
R42666 vdd.n359 vdd.t1836 7.146
R42667 vdd.n359 vdd.t964 7.146
R42668 vdd.n348 vdd.t2097 7.146
R42669 vdd.n348 vdd.t1218 7.146
R42670 vdd.n347 vdd.t1683 7.146
R42671 vdd.n347 vdd.t2011 7.146
R42672 vdd.n346 vdd.t1929 7.146
R42673 vdd.n346 vdd.t2263 7.146
R42674 vdd.n345 vdd.t79 7.146
R42675 vdd.n345 vdd.t409 7.146
R42676 vdd.n344 vdd.t491 7.146
R42677 vdd.n344 vdd.t813 7.146
R42678 vdd.n343 vdd.t751 7.146
R42679 vdd.n343 vdd.t1046 7.146
R42680 vdd.n342 vdd.t1858 7.146
R42681 vdd.n342 vdd.t2191 7.146
R42682 vdd.n341 vdd.t1388 7.146
R42683 vdd.n341 vdd.t1706 7.146
R42684 vdd.n340 vdd.t2517 7.146
R42685 vdd.n340 vdd.t2844 7.146
R42686 vdd.n339 vdd.t2938 7.146
R42687 vdd.n339 vdd.t284 7.146
R42688 vdd.n338 vdd.t19 7.146
R42689 vdd.n338 vdd.t2268 7.146
R42690 vdd.n337 vdd.t1827 7.146
R42691 vdd.n337 vdd.t2158 7.146
R42692 vdd.n336 vdd.t675 7.146
R42693 vdd.n336 vdd.t2793 7.146
R42694 vdd.n335 vdd.t2523 7.146
R42695 vdd.n335 vdd.t1650 7.146
R42696 vdd.n334 vdd.t1391 7.146
R42697 vdd.n334 vdd.t531 7.146
R42698 vdd.n333 vdd.t1864 7.146
R42699 vdd.n333 vdd.t986 7.146
R42700 vdd.n332 vdd.t753 7.146
R42701 vdd.n332 vdd.t2870 7.146
R42702 vdd.n331 vdd.t496 7.146
R42703 vdd.n331 vdd.t2619 7.146
R42704 vdd.n330 vdd.t84 7.146
R42705 vdd.n330 vdd.t2210 7.146
R42706 vdd.n539 vdd.t668 7.146
R42707 vdd.n539 vdd.t66 7.146
R42708 vdd.n528 vdd.t898 7.146
R42709 vdd.n528 vdd.t311 7.146
R42710 vdd.n527 vdd.t2 7.146
R42711 vdd.n527 vdd.t364 7.146
R42712 vdd.n526 vdd.t268 7.146
R42713 vdd.n526 vdd.t609 7.146
R42714 vdd.n525 vdd.t1385 7.146
R42715 vdd.n525 vdd.t1732 7.146
R42716 vdd.n524 vdd.t1792 7.146
R42717 vdd.n524 vdd.t2145 7.146
R42718 vdd.n523 vdd.t2053 7.146
R42719 vdd.n523 vdd.t2384 7.146
R42720 vdd.n522 vdd.t197 7.146
R42721 vdd.n522 vdd.t538 7.146
R42722 vdd.n521 vdd.t2721 7.146
R42723 vdd.n521 vdd.t56 7.146
R42724 vdd.n520 vdd.t840 7.146
R42725 vdd.n520 vdd.t1179 7.146
R42726 vdd.n519 vdd.t1252 7.146
R42727 vdd.n519 vdd.t1596 7.146
R42728 vdd.n518 vdd.t1608 7.146
R42729 vdd.n518 vdd.t1513 7.146
R42730 vdd.n517 vdd.t173 7.146
R42731 vdd.n517 vdd.t512 7.146
R42732 vdd.n516 vdd.t2472 7.146
R42733 vdd.n516 vdd.t1867 7.146
R42734 vdd.n515 vdd.t1334 7.146
R42735 vdd.n515 vdd.t755 7.146
R42736 vdd.n514 vdd.t222 7.146
R42737 vdd.n514 vdd.t2606 7.146
R42738 vdd.n513 vdd.t699 7.146
R42739 vdd.n513 vdd.t90 7.146
R42740 vdd.n512 vdd.t2545 7.146
R42741 vdd.n512 vdd.t1934 7.146
R42742 vdd.n511 vdd.t2299 7.146
R42743 vdd.n511 vdd.t1694 7.146
R42744 vdd.n510 vdd.t1882 7.146
R42745 vdd.n510 vdd.t1269 7.146
R42746 vdd.n719 vdd.t2468 7.146
R42747 vdd.n719 vdd.t1863 7.146
R42748 vdd.n708 vdd.t2732 7.146
R42749 vdd.n708 vdd.t2112 7.146
R42750 vdd.n707 vdd.t1309 7.146
R42751 vdd.n707 vdd.t1658 7.146
R42752 vdd.n706 vdd.t1567 7.146
R42753 vdd.n706 vdd.t1913 7.146
R42754 vdd.n705 vdd.t2717 7.146
R42755 vdd.n705 vdd.t52 7.146
R42756 vdd.n704 vdd.t132 7.146
R42757 vdd.n704 vdd.t470 7.146
R42758 vdd.n703 vdd.t381 7.146
R42759 vdd.n703 vdd.t726 7.146
R42760 vdd.n702 vdd.t1491 7.146
R42761 vdd.n702 vdd.t1830 7.146
R42762 vdd.n701 vdd.t1009 7.146
R42763 vdd.n701 vdd.t1364 7.146
R42764 vdd.n700 vdd.t2156 7.146
R42765 vdd.n700 vdd.t2493 7.146
R42766 vdd.n699 vdd.t2584 7.146
R42767 vdd.n699 vdd.t2923 7.146
R42768 vdd.n698 vdd.t234 7.146
R42769 vdd.n698 vdd.t140 7.146
R42770 vdd.n697 vdd.t1460 7.146
R42771 vdd.n697 vdd.t1808 7.146
R42772 vdd.n696 vdd.t1276 7.146
R42773 vdd.n696 vdd.t702 7.146
R42774 vdd.n695 vdd.t170 7.146
R42775 vdd.n695 vdd.t2547 7.146
R42776 vdd.n694 vdd.t2022 7.146
R42777 vdd.n694 vdd.t1403 7.146
R42778 vdd.n693 vdd.t2486 7.146
R42779 vdd.n693 vdd.t1886 7.146
R42780 vdd.n692 vdd.t1357 7.146
R42781 vdd.n692 vdd.t770 7.146
R42782 vdd.n691 vdd.t1111 7.146
R42783 vdd.n691 vdd.t520 7.146
R42784 vdd.n690 vdd.t718 7.146
R42785 vdd.n690 vdd.t107 7.146
R42786 vdd.n899 vdd.t1547 7.146
R42787 vdd.n899 vdd.t698 7.146
R42788 vdd.n888 vdd.t1786 7.146
R42789 vdd.n888 vdd.t915 7.146
R42790 vdd.n887 vdd.t2663 7.146
R42791 vdd.n887 vdd.t2977 7.146
R42792 vdd.n886 vdd.t2913 7.146
R42793 vdd.n886 vdd.t248 7.146
R42794 vdd.n885 vdd.t1037 7.146
R42795 vdd.n885 vdd.t1363 7.146
R42796 vdd.n884 vdd.t1450 7.146
R42797 vdd.n884 vdd.t1775 7.146
R42798 vdd.n883 vdd.t1701 7.146
R42799 vdd.n883 vdd.t2029 7.146
R42800 vdd.n882 vdd.t2835 7.146
R42801 vdd.n882 vdd.t175 7.146
R42802 vdd.n881 vdd.t2350 7.146
R42803 vdd.n881 vdd.t2694 7.146
R42804 vdd.n880 vdd.t504 7.146
R42805 vdd.n880 vdd.t826 7.146
R42806 vdd.n879 vdd.t904 7.146
R42807 vdd.n879 vdd.t1231 7.146
R42808 vdd.n878 vdd.t2467 7.146
R42809 vdd.n878 vdd.t1720 7.146
R42810 vdd.n877 vdd.t2807 7.146
R42811 vdd.n877 vdd.t154 7.146
R42812 vdd.n876 vdd.t386 7.146
R42813 vdd.n876 vdd.t2490 7.146
R42814 vdd.n875 vdd.t2239 7.146
R42815 vdd.n875 vdd.t1361 7.146
R42816 vdd.n874 vdd.t1095 7.146
R42817 vdd.n874 vdd.t246 7.146
R42818 vdd.n873 vdd.t1570 7.146
R42819 vdd.n873 vdd.t722 7.146
R42820 vdd.n872 vdd.t449 7.146
R42821 vdd.n872 vdd.t2576 7.146
R42822 vdd.n871 vdd.t208 7.146
R42823 vdd.n871 vdd.t2315 7.146
R42824 vdd.n870 vdd.t2778 7.146
R42825 vdd.n870 vdd.t1908 7.146
R42826 vdd.n1079 vdd.t380 7.146
R42827 vdd.n1079 vdd.t2152 7.146
R42828 vdd.n1068 vdd.t617 7.146
R42829 vdd.n1068 vdd.t2388 7.146
R42830 vdd.n1067 vdd.t960 7.146
R42831 vdd.n1067 vdd.t2309 7.146
R42832 vdd.n1066 vdd.t1214 7.146
R42833 vdd.n1066 vdd.t2569 7.146
R42834 vdd.n1065 vdd.t2346 7.146
R42835 vdd.n1065 vdd.t717 7.146
R42836 vdd.n1064 vdd.t2777 7.146
R42837 vdd.n1064 vdd.t1108 7.146
R42838 vdd.n1063 vdd.t18 7.146
R42839 vdd.n1063 vdd.t1354 7.146
R42840 vdd.n1062 vdd.t1142 7.146
R42841 vdd.n1062 vdd.t2483 7.146
R42842 vdd.n1061 vdd.t692 7.146
R42843 vdd.n1061 vdd.t2018 7.146
R42844 vdd.n1060 vdd.t1802 7.146
R42845 vdd.n1060 vdd.t169 7.146
R42846 vdd.n1059 vdd.t2238 7.146
R42847 vdd.n1059 vdd.t586 7.146
R42848 vdd.n1058 vdd.t1076 7.146
R42849 vdd.n1058 vdd.t2578 7.146
R42850 vdd.n1057 vdd.t1121 7.146
R42851 vdd.n1057 vdd.t2459 7.146
R42852 vdd.n1056 vdd.t2183 7.146
R42853 vdd.n1056 vdd.t957 7.146
R42854 vdd.n1055 vdd.t1036 7.146
R42855 vdd.n1055 vdd.t2832 7.146
R42856 vdd.n1054 vdd.t2912 7.146
R42857 vdd.n1054 vdd.t1696 7.146
R42858 vdd.n1053 vdd.t404 7.146
R42859 vdd.n1053 vdd.t2179 7.146
R42860 vdd.n1052 vdd.t2257 7.146
R42861 vdd.n1052 vdd.t1029 7.146
R42862 vdd.n1051 vdd.t2004 7.146
R42863 vdd.n1051 vdd.t807 7.146
R42864 vdd.n1050 vdd.t1585 7.146
R42865 vdd.n1050 vdd.t399 7.146
R42866 vdd.n1259 vdd.t2178 7.146
R42867 vdd.n1259 vdd.t1979 7.146
R42868 vdd.n1248 vdd.t2407 7.146
R42869 vdd.n1248 vdd.t2237 7.146
R42870 vdd.n1247 vdd.t2291 7.146
R42871 vdd.n1247 vdd.t2889 7.146
R42872 vdd.n1246 vdd.t2536 7.146
R42873 vdd.n1246 vdd.t139 7.146
R42874 vdd.n1245 vdd.t688 7.146
R42875 vdd.n1245 vdd.t1255 7.146
R42876 vdd.n1244 vdd.t1094 7.146
R42877 vdd.n1244 vdd.t1668 7.146
R42878 vdd.n1243 vdd.t1326 7.146
R42879 vdd.n1243 vdd.t1919 7.146
R42880 vdd.n1242 vdd.t2463 7.146
R42881 vdd.n1242 vdd.t62 7.146
R42882 vdd.n1241 vdd.t1990 7.146
R42883 vdd.n1241 vdd.t2590 7.146
R42884 vdd.n1240 vdd.t148 7.146
R42885 vdd.n1240 vdd.t735 7.146
R42886 vdd.n1239 vdd.t557 7.146
R42887 vdd.n1239 vdd.t1125 7.146
R42888 vdd.n1238 vdd.t2680 7.146
R42889 vdd.n1238 vdd.t1940 7.146
R42890 vdd.n1237 vdd.t2436 7.146
R42891 vdd.n1237 vdd.t32 7.146
R42892 vdd.n1236 vdd.t976 7.146
R42893 vdd.n1236 vdd.t809 7.146
R42894 vdd.n1235 vdd.t2855 7.146
R42895 vdd.n1235 vdd.t2666 7.146
R42896 vdd.n1234 vdd.t1716 7.146
R42897 vdd.n1234 vdd.t1518 7.146
R42898 vdd.n1233 vdd.t2204 7.146
R42899 vdd.n1233 vdd.t2006 7.146
R42900 vdd.n1232 vdd.t1058 7.146
R42901 vdd.n1232 vdd.t864 7.146
R42902 vdd.n1231 vdd.t822 7.146
R42903 vdd.n1231 vdd.t631 7.146
R42904 vdd.n1230 vdd.t417 7.146
R42905 vdd.n1230 vdd.t226 7.146
R42906 vdd.n1439 vdd.t2005 7.146
R42907 vdd.n1439 vdd.t47 7.146
R42908 vdd.n1428 vdd.t2256 7.146
R42909 vdd.n1428 vdd.t300 7.146
R42910 vdd.n1427 vdd.t2859 7.146
R42911 vdd.n1427 vdd.t1963 7.146
R42912 vdd.n1426 vdd.t115 7.146
R42913 vdd.n1426 vdd.t2227 7.146
R42914 vdd.n1425 vdd.t1234 7.146
R42915 vdd.n1425 vdd.t365 7.146
R42916 vdd.n1424 vdd.t1643 7.146
R42917 vdd.n1424 vdd.t792 7.146
R42918 vdd.n1423 vdd.t1896 7.146
R42919 vdd.n1423 vdd.t1001 7.146
R42920 vdd.n1422 vdd.t36 7.146
R42921 vdd.n1422 vdd.t2147 7.146
R42922 vdd.n1421 vdd.t2561 7.146
R42923 vdd.n1421 vdd.t1663 7.146
R42924 vdd.n1420 vdd.t710 7.146
R42925 vdd.n1420 vdd.t2802 7.146
R42926 vdd.n1419 vdd.t1106 7.146
R42927 vdd.n1419 vdd.t245 7.146
R42928 vdd.n1418 vdd.t2061 7.146
R42929 vdd.n1418 vdd.t443 7.146
R42930 vdd.n1417 vdd.t8 7.146
R42931 vdd.n1417 vdd.t2119 7.146
R42932 vdd.n1416 vdd.t825 7.146
R42933 vdd.n1416 vdd.t1849 7.146
R42934 vdd.n1415 vdd.t2693 7.146
R42935 vdd.n1415 vdd.t743 7.146
R42936 vdd.n1414 vdd.t1543 7.146
R42937 vdd.n1414 vdd.t2595 7.146
R42938 vdd.n1413 vdd.t2031 7.146
R42939 vdd.n1413 vdd.t74 7.146
R42940 vdd.n1412 vdd.t883 7.146
R42941 vdd.n1412 vdd.t1924 7.146
R42942 vdd.n1411 vdd.t648 7.146
R42943 vdd.n1411 vdd.t1677 7.146
R42944 vdd.n1410 vdd.t250 7.146
R42945 vdd.n1410 vdd.t1263 7.146
R42946 vdd.n1619 vdd.t479 7.146
R42947 vdd.n1619 vdd.t1843 7.146
R42948 vdd.n1608 vdd.t738 7.146
R42949 vdd.n1608 vdd.t2099 7.146
R42950 vdd.n1607 vdd.t2200 7.146
R42951 vdd.n1607 vdd.t303 7.146
R42952 vdd.n1606 vdd.t2426 7.146
R42953 vdd.n1606 vdd.t542 7.146
R42954 vdd.n1605 vdd.t590 7.146
R42955 vdd.n1605 vdd.t1659 7.146
R42956 vdd.n1604 vdd.t971 7.146
R42957 vdd.n1604 vdd.t2092 7.146
R42958 vdd.n1603 vdd.t1226 7.146
R42959 vdd.n1603 vdd.t2318 7.146
R42960 vdd.n1602 vdd.t2360 7.146
R42961 vdd.n1602 vdd.t472 7.146
R42962 vdd.n1601 vdd.t1885 7.146
R42963 vdd.n1601 vdd.t2981 7.146
R42964 vdd.n1600 vdd.t28 7.146
R42965 vdd.n1600 vdd.t1118 7.146
R42966 vdd.n1599 vdd.t456 7.146
R42967 vdd.n1599 vdd.t1534 7.146
R42968 vdd.n1598 vdd.t2903 7.146
R42969 vdd.n1598 vdd.t2030 7.146
R42970 vdd.n1597 vdd.t2327 7.146
R42971 vdd.n1597 vdd.t454 7.146
R42972 vdd.n1596 vdd.t2290 7.146
R42973 vdd.n1596 vdd.t683 7.146
R42974 vdd.n1595 vdd.t1144 7.146
R42975 vdd.n1595 vdd.t2531 7.146
R42976 vdd.n1594 vdd.t23 7.146
R42977 vdd.n1594 vdd.t1396 7.146
R42978 vdd.n1593 vdd.t503 7.146
R42979 vdd.n1593 vdd.t1872 7.146
R42980 vdd.n1592 vdd.t2349 7.146
R42981 vdd.n1592 vdd.t757 7.146
R42982 vdd.n1591 vdd.t2115 7.146
R42983 vdd.n1591 vdd.t501 7.146
R42984 vdd.n1590 vdd.t1700 7.146
R42985 vdd.n1590 vdd.t97 7.146
R42986 vdd.n1799 vdd.t273 7.146
R42987 vdd.n1799 vdd.t419 7.146
R42988 vdd.n1788 vdd.t502 7.146
R42989 vdd.n1788 vdd.t650 7.146
R42990 vdd.n1787 vdd.t1614 7.146
R42991 vdd.n1787 vdd.t1181 7.146
R42992 vdd.n1786 vdd.t1857 7.146
R42993 vdd.n1786 vdd.t1424 7.146
R42994 vdd.n1785 vdd.t0 7.146
R42995 vdd.n1785 vdd.t2580 7.146
R42996 vdd.n1784 vdd.t433 7.146
R42997 vdd.n1784 vdd.t2980 7.146
R42998 vdd.n1783 vdd.t667 7.146
R42999 vdd.n1783 vdd.t251 7.146
R43000 vdd.n1782 vdd.t1789 7.146
R43001 vdd.n1782 vdd.t1367 7.146
R43002 vdd.n1781 vdd.t1311 7.146
R43003 vdd.n1781 vdd.t886 7.146
R43004 vdd.n1780 vdd.t2451 7.146
R43005 vdd.n1780 vdd.t2034 7.146
R43006 vdd.n1779 vdd.t2878 7.146
R43007 vdd.n1779 vdd.t2432 7.146
R43008 vdd.n1778 vdd.t374 7.146
R43009 vdd.n1778 vdd.t403 7.146
R43010 vdd.n1777 vdd.t1771 7.146
R43011 vdd.n1777 vdd.t1333 7.146
R43012 vdd.n1776 vdd.t2080 7.146
R43013 vdd.n1776 vdd.t2229 7.146
R43014 vdd.n1775 vdd.t923 7.146
R43015 vdd.n1775 vdd.t1082 7.146
R43016 vdd.n1774 vdd.t2792 7.146
R43017 vdd.n1774 vdd.t2945 7.146
R43018 vdd.n1773 vdd.t294 7.146
R43019 vdd.n1773 vdd.t437 7.146
R43020 vdd.n1772 vdd.t2131 7.146
R43021 vdd.n1772 vdd.t2285 7.146
R43022 vdd.n1771 vdd.t1891 7.146
R43023 vdd.n1771 vdd.t2049 7.146
R43024 vdd.n1770 vdd.t1466 7.146
R43025 vdd.n1770 vdd.t1618 7.146
R43026 vdd.n1979 vdd.t100 7.146
R43027 vdd.n1979 vdd.t2223 7.146
R43028 vdd.n1968 vdd.t335 7.146
R43029 vdd.n1968 vdd.t2450 7.146
R43030 vdd.n1967 vdd.t2189 7.146
R43031 vdd.n1967 vdd.t2496 7.146
R43032 vdd.n1966 vdd.t2418 7.146
R43033 vdd.n1966 vdd.t2759 7.146
R43034 vdd.n1965 vdd.t580 7.146
R43035 vdd.n1965 vdd.t882 7.146
R43036 vdd.n1964 vdd.t965 7.146
R43037 vdd.n1964 vdd.t1286 7.146
R43038 vdd.n1963 vdd.t1219 7.146
R43039 vdd.n1963 vdd.t1542 7.146
R43040 vdd.n1962 vdd.t2351 7.146
R43041 vdd.n1962 vdd.t2692 7.146
R43042 vdd.n1961 vdd.t1881 7.146
R43043 vdd.n1961 vdd.t2212 7.146
R43044 vdd.n1960 vdd.t22 7.146
R43045 vdd.n1960 vdd.t352 7.146
R43046 vdd.n1959 vdd.t450 7.146
R43047 vdd.n1959 vdd.t775 7.146
R43048 vdd.n1958 vdd.t2745 7.146
R43049 vdd.n1958 vdd.t1978 7.146
R43050 vdd.n1957 vdd.t2322 7.146
R43051 vdd.n1957 vdd.t2657 7.146
R43052 vdd.n1956 vdd.t1899 7.146
R43053 vdd.n1956 vdd.t1020 7.146
R43054 vdd.n1955 vdd.t779 7.146
R43055 vdd.n1955 vdd.t2902 7.146
R43056 vdd.n1954 vdd.t2628 7.146
R43057 vdd.n1954 vdd.t1758 7.146
R43058 vdd.n1953 vdd.t118 7.146
R43059 vdd.n1953 vdd.t2241 7.146
R43060 vdd.n1952 vdd.t1955 7.146
R43061 vdd.n1952 vdd.t1100 7.146
R43062 vdd.n1951 vdd.t1722 7.146
R43063 vdd.n1951 vdd.t849 7.146
R43064 vdd.n1950 vdd.t1293 7.146
R43065 vdd.n1950 vdd.t451 7.146
R43066 vdd.n2159 vdd.t1894 7.146
R43067 vdd.n2159 vdd.t1014 7.146
R43068 vdd.n2148 vdd.t2132 7.146
R43069 vdd.n2148 vdd.t1264 7.146
R43070 vdd.n2147 vdd.t511 7.146
R43071 vdd.n2147 vdd.t828 7.146
R43072 vdd.n2146 vdd.t765 7.146
R43073 vdd.n2146 vdd.t1066 7.146
R43074 vdd.n2145 vdd.t1875 7.146
R43075 vdd.n2145 vdd.t2209 7.146
R43076 vdd.n2144 vdd.t2294 7.146
R43077 vdd.n2144 vdd.t2616 7.146
R43078 vdd.n2143 vdd.t2538 7.146
R43079 vdd.n2143 vdd.t2865 7.146
R43080 vdd.n2142 vdd.t691 7.146
R43081 vdd.n2142 vdd.t984 7.146
R43082 vdd.n2141 vdd.t215 7.146
R43083 vdd.n2141 vdd.t530 7.146
R43084 vdd.n2140 vdd.t1328 7.146
R43085 vdd.n2140 vdd.t1648 7.146
R43086 vdd.n2139 vdd.t1753 7.146
R43087 vdd.n2139 vdd.t2083 7.146
R43088 vdd.n2138 vdd.t1325 7.146
R43089 vdd.n2138 vdd.t599 7.146
R43090 vdd.n2137 vdd.t658 7.146
R43091 vdd.n2137 vdd.t958 7.146
R43092 vdd.n2136 vdd.t729 7.146
R43093 vdd.n2136 vdd.t2839 7.146
R43094 vdd.n2135 vdd.t2585 7.146
R43095 vdd.n2135 vdd.t1703 7.146
R43096 vdd.n2134 vdd.t1429 7.146
R43097 vdd.n2134 vdd.t587 7.146
R43098 vdd.n2133 vdd.t1915 7.146
R43099 vdd.n2133 vdd.t1040 7.146
R43100 vdd.n2132 vdd.t794 7.146
R43101 vdd.n2132 vdd.t2916 7.146
R43102 vdd.n2131 vdd.t547 7.146
R43103 vdd.n2131 vdd.t2672 7.146
R43104 vdd.n2130 vdd.t135 7.146
R43105 vdd.n2130 vdd.t2259 7.146
R43106 vdd.n2339 vdd.t725 7.146
R43107 vdd.n2339 vdd.t2770 7.146
R43108 vdd.n2328 vdd.t937 7.146
R43109 vdd.n2328 vdd.t4 7.146
R43110 vdd.n2327 vdd.t1806 7.146
R43111 vdd.n2327 vdd.t196 7.146
R43112 vdd.n2326 vdd.t2069 7.146
R43113 vdd.n2326 vdd.t442 7.146
R43114 vdd.n2325 vdd.t212 7.146
R43115 vdd.n2325 vdd.t1562 7.146
R43116 vdd.n2324 vdd.t621 7.146
R43117 vdd.n2324 vdd.t1970 7.146
R43118 vdd.n2323 vdd.t857 7.146
R43119 vdd.n2323 vdd.t2231 7.146
R43120 vdd.n2322 vdd.t1992 7.146
R43121 vdd.n2322 vdd.t372 7.146
R43122 vdd.n2321 vdd.t1510 7.146
R43123 vdd.n2321 vdd.t2888 7.146
R43124 vdd.n2320 vdd.t2655 7.146
R43125 vdd.n2320 vdd.t1004 7.146
R43126 vdd.n2319 vdd.t78 7.146
R43127 vdd.n2319 vdd.t1423 7.146
R43128 vdd.n2318 vdd.t2934 7.146
R43129 vdd.n2318 vdd.t2091 7.146
R43130 vdd.n2317 vdd.t1957 7.146
R43131 vdd.n2317 vdd.t340 7.146
R43132 vdd.n2316 vdd.t2516 7.146
R43133 vdd.n2316 vdd.t1576 7.146
R43134 vdd.n2315 vdd.t1386 7.146
R43135 vdd.n2315 vdd.t458 7.146
R43136 vdd.n2314 vdd.t271 7.146
R43137 vdd.n2314 vdd.t2302 7.146
R43138 vdd.n2313 vdd.t748 7.146
R43139 vdd.n2313 vdd.t2782 7.146
R43140 vdd.n2312 vdd.t2600 7.146
R43141 vdd.n2312 vdd.t1638 7.146
R43142 vdd.n2311 vdd.t2336 7.146
R43143 vdd.n2311 vdd.t1400 7.146
R43144 vdd.n2310 vdd.t1928 7.146
R43145 vdd.n2310 vdd.t972 7.146
R43146 vdd.n2519 vdd.t545 7.146
R43147 vdd.n2519 vdd.t1573 7.146
R43148 vdd.n2508 vdd.t795 7.146
R43149 vdd.n2508 vdd.t1807 7.146
R43150 vdd.n2507 vdd.t2369 7.146
R43151 vdd.n2507 vdd.t1488 7.146
R43152 vdd.n2506 vdd.t2626 7.146
R43153 vdd.n2506 vdd.t1741 7.146
R43154 vdd.n2505 vdd.t777 7.146
R43155 vdd.n2505 vdd.t2883 7.146
R43156 vdd.n2504 vdd.t1169 7.146
R43157 vdd.n2504 vdd.t305 7.146
R43158 vdd.n2503 vdd.t1414 7.146
R43159 vdd.n2503 vdd.t546 7.146
R43160 vdd.n2502 vdd.t2560 7.146
R43161 vdd.n2502 vdd.t1662 7.146
R43162 vdd.n2501 vdd.t2087 7.146
R43163 vdd.n2501 vdd.t1187 7.146
R43164 vdd.n2500 vdd.t232 7.146
R43165 vdd.n2500 vdd.t2319 7.146
R43166 vdd.n2499 vdd.t636 7.146
R43167 vdd.n2499 vdd.t2755 7.146
R43168 vdd.n2498 vdd.t2303 7.146
R43169 vdd.n2498 vdd.t701 7.146
R43170 vdd.n2497 vdd.t2526 7.146
R43171 vdd.n2497 vdd.t1637 7.146
R43172 vdd.n2496 vdd.t2344 7.146
R43173 vdd.n2496 vdd.t410 7.146
R43174 vdd.n2495 vdd.t1213 7.146
R43175 vdd.n2495 vdd.t2264 7.146
R43176 vdd.n2494 vdd.t96 7.146
R43177 vdd.n2494 vdd.t1116 7.146
R43178 vdd.n2493 vdd.t574 7.146
R43179 vdd.n2493 vdd.t1593 7.146
R43180 vdd.n2492 vdd.t2408 7.146
R43181 vdd.n2492 vdd.t466 7.146
R43182 vdd.n2491 vdd.t2182 7.146
R43183 vdd.n2491 vdd.t233 7.146
R43184 vdd.n2490 vdd.t1761 7.146
R43185 vdd.n2490 vdd.t2795 7.146
R43186 vdd.n2699 vdd.t1592 7.146
R43187 vdd.n2699 vdd.t406 7.146
R43188 vdd.n2688 vdd.t1826 7.146
R43189 vdd.n2688 vdd.t633 7.146
R43190 vdd.n2687 vdd.t1463 7.146
R43191 vdd.n2687 vdd.t2805 7.146
R43192 vdd.n2686 vdd.t1715 7.146
R43193 vdd.n2686 vdd.t65 7.146
R43194 vdd.n2685 vdd.t2854 7.146
R43195 vdd.n2685 vdd.t1182 7.146
R43196 vdd.n2684 vdd.t292 7.146
R43197 vdd.n2684 vdd.t1598 7.146
R43198 vdd.n2683 vdd.t524 7.146
R43199 vdd.n2683 vdd.t1839 7.146
R43200 vdd.n2682 vdd.t1641 7.146
R43201 vdd.n2682 vdd.t2986 7.146
R43202 vdd.n2681 vdd.t1163 7.146
R43203 vdd.n2681 vdd.t2501 7.146
R43204 vdd.n2680 vdd.t2304 7.146
R43205 vdd.n2680 vdd.t653 7.146
R43206 vdd.n2679 vdd.t2738 7.146
R43207 vdd.n2679 vdd.t1064 7.146
R43208 vdd.n2678 vdd.t802 7.146
R43209 vdd.n2678 vdd.t2283 7.146
R43210 vdd.n2677 vdd.t1617 7.146
R43211 vdd.n2677 vdd.t2961 7.146
R43212 vdd.n2676 vdd.t432 7.146
R43213 vdd.n2676 vdd.t2211 7.146
R43214 vdd.n2675 vdd.t2276 7.146
R43215 vdd.n2675 vdd.t1070 7.146
R43216 vdd.n2674 vdd.t1131 7.146
R43217 vdd.n2674 vdd.t2931 7.146
R43218 vdd.n2673 vdd.t1607 7.146
R43219 vdd.n2673 vdd.t427 7.146
R43220 vdd.n2672 vdd.t483 7.146
R43221 vdd.n2672 vdd.t2271 7.146
R43222 vdd.n2671 vdd.t256 7.146
R43223 vdd.n2671 vdd.t2036 7.146
R43224 vdd.n2670 vdd.t2815 7.146
R43225 vdd.n2670 vdd.t1603 7.146
R43226 vdd.n2879 vdd.t426 7.146
R43227 vdd.n2879 vdd.t237 7.146
R43228 vdd.n2868 vdd.t656 7.146
R43229 vdd.n2868 vdd.t467 7.146
R43230 vdd.n2867 vdd.t2786 7.146
R43231 vdd.n2867 vdd.t394 7.146
R43232 vdd.n2866 vdd.t37 7.146
R43233 vdd.n2866 vdd.t626 7.146
R43234 vdd.n2865 vdd.t1157 7.146
R43235 vdd.n2865 vdd.t1757 7.146
R43236 vdd.n2864 vdd.t1586 7.146
R43237 vdd.n2864 vdd.t2173 7.146
R43238 vdd.n2863 vdd.t1820 7.146
R43239 vdd.n2863 vdd.t2405 7.146
R43240 vdd.n2862 vdd.t2963 7.146
R43241 vdd.n2862 vdd.t571 7.146
R43242 vdd.n2861 vdd.t2478 7.146
R43243 vdd.n2861 vdd.t83 7.146
R43244 vdd.n2860 vdd.t632 7.146
R43245 vdd.n2860 vdd.t1207 7.146
R43246 vdd.n2859 vdd.t1035 7.146
R43247 vdd.n2859 vdd.t1622 7.146
R43248 vdd.n2858 vdd.t2381 7.146
R43249 vdd.n2858 vdd.t1652 7.146
R43250 vdd.n2857 vdd.t2939 7.146
R43251 vdd.n2857 vdd.t535 7.146
R43252 vdd.n2856 vdd.t2234 7.146
R43253 vdd.n2856 vdd.t2041 7.146
R43254 vdd.n2855 vdd.t1089 7.146
R43255 vdd.n2855 vdd.t894 7.146
R43256 vdd.n2854 vdd.t2953 7.146
R43257 vdd.n2854 vdd.t2768 7.146
R43258 vdd.n2853 vdd.t447 7.146
R43259 vdd.n2853 vdd.t259 7.146
R43260 vdd.n2852 vdd.t2287 7.146
R43261 vdd.n2852 vdd.t2102 7.146
R43262 vdd.n2851 vdd.t2060 7.146
R43263 vdd.n2851 vdd.t1848 7.146
R43264 vdd.n2850 vdd.t1628 7.146
R43265 vdd.n2850 vdd.t1433 7.146
R43266 vdd.n3059 vdd.t2908 7.146
R43267 vdd.n3059 vdd.t2038 7.146
R43268 vdd.n3048 vdd.t160 7.146
R43269 vdd.n3048 vdd.t2274 7.146
R43270 vdd.n3047 vdd.t1370 7.146
R43271 vdd.n3047 vdd.t1686 7.146
R43272 vdd.n3046 vdd.t1604 7.146
R43273 vdd.n3046 vdd.t1930 7.146
R43274 vdd.n3045 vdd.t2758 7.146
R43275 vdd.n3045 vdd.t81 7.146
R43276 vdd.n3044 vdd.t183 7.146
R43277 vdd.n3044 vdd.t494 7.146
R43278 vdd.n3043 vdd.t429 7.146
R43279 vdd.n3043 vdd.t752 7.146
R43280 vdd.n3042 vdd.t1541 7.146
R43281 vdd.n3042 vdd.t1861 7.146
R43282 vdd.n3041 vdd.t1072 7.146
R43283 vdd.n3041 vdd.t1389 7.146
R43284 vdd.n3040 vdd.t2214 7.146
R43285 vdd.n3040 vdd.t2522 7.146
R43286 vdd.n3039 vdd.t2623 7.146
R43287 vdd.n3039 vdd.t2943 7.146
R43288 vdd.n3038 vdd.t1000 7.146
R43289 vdd.n3038 vdd.t279 7.146
R43290 vdd.n3037 vdd.t1511 7.146
R43291 vdd.n3037 vdd.t1828 7.146
R43292 vdd.n3036 vdd.t1712 7.146
R43293 vdd.n3036 vdd.t843 7.146
R43294 vdd.n3035 vdd.t597 7.146
R43295 vdd.n3035 vdd.t2724 7.146
R43296 vdd.n3034 vdd.t2429 7.146
R43297 vdd.n3034 vdd.t1572 7.146
R43298 vdd.n3033 vdd.t2922 7.146
R43299 vdd.n3033 vdd.t2062 7.146
R43300 vdd.n3032 vdd.t1778 7.146
R43301 vdd.n3032 vdd.t903 7.146
R43302 vdd.n3031 vdd.t1533 7.146
R43303 vdd.n3031 vdd.t682 7.146
R43304 vdd.n3030 vdd.t1117 7.146
R43305 vdd.n3030 vdd.t275 7.146
R43306 vdd.n3239 vdd.t1708 7.146
R43307 vdd.n3239 vdd.t103 7.146
R43308 vdd.n3228 vdd.t1946 7.146
R43309 vdd.n3228 vdd.t339 7.146
R43310 vdd.n3227 vdd.t2700 7.146
R43311 vdd.n3227 vdd.t799 7.146
R43312 vdd.n3226 vdd.t2930 7.146
R43313 vdd.n3226 vdd.t1019 7.146
R43314 vdd.n3225 vdd.t1065 7.146
R43315 vdd.n3225 vdd.t2162 7.146
R43316 vdd.n3224 vdd.t1475 7.146
R43317 vdd.n3224 vdd.t2593 7.146
R43318 vdd.n3223 vdd.t1727 7.146
R43319 vdd.n3223 vdd.t2821 7.146
R43320 vdd.n3222 vdd.t2869 7.146
R43321 vdd.n3222 vdd.t949 7.146
R43322 vdd.n3221 vdd.t2375 7.146
R43323 vdd.n3221 vdd.t488 7.146
R43324 vdd.n3220 vdd.t529 7.146
R43325 vdd.n3220 vdd.t1612 7.146
R43326 vdd.n3219 vdd.t927 7.146
R43327 vdd.n3219 vdd.t2045 7.146
R43328 vdd.n3218 vdd.t2615 7.146
R43329 vdd.n3218 vdd.t1740 7.146
R43330 vdd.n3217 vdd.t2834 7.146
R43331 vdd.n3217 vdd.t926 7.146
R43332 vdd.n3216 vdd.t534 7.146
R43333 vdd.n3216 vdd.t1907 7.146
R43334 vdd.n3215 vdd.t2382 7.146
R43335 vdd.n3215 vdd.t788 7.146
R43336 vdd.n3214 vdd.t1250 7.146
R43337 vdd.n3214 vdd.t2633 7.146
R43338 vdd.n3213 vdd.t1731 7.146
R43339 vdd.n3213 vdd.t125 7.146
R43340 vdd.n3212 vdd.t608 7.146
R43341 vdd.n3212 vdd.t1962 7.146
R43342 vdd.n3211 vdd.t363 7.146
R43343 vdd.n3211 vdd.t1730 7.146
R43344 vdd.n3210 vdd.t2935 7.146
R43345 vdd.n3210 vdd.t1304 7.146
R43346 vdd.n3419 vdd.t528 7.146
R43347 vdd.n3419 vdd.t2921 7.146
R43348 vdd.n3408 vdd.t783 7.146
R43349 vdd.n3408 vdd.t176 7.146
R43350 vdd.n3407 vdd.t990 7.146
R43351 vdd.n3407 vdd.t1342 7.146
R43352 vdd.n3406 vdd.t1245 7.146
R43353 vdd.n3406 vdd.t1589 7.146
R43354 vdd.n3405 vdd.t2371 7.146
R43355 vdd.n3405 vdd.t2739 7.146
R43356 vdd.n3404 vdd.t2794 7.146
R43357 vdd.n3404 vdd.t164 7.146
R43358 vdd.n3403 vdd.t46 7.146
R43359 vdd.n3403 vdd.t405 7.146
R43360 vdd.n3402 vdd.t1170 7.146
R43361 vdd.n3402 vdd.t1515 7.146
R43362 vdd.n3401 vdd.t721 7.146
R43363 vdd.n3401 vdd.t1044 7.146
R43364 vdd.n3400 vdd.t1825 7.146
R43365 vdd.n3400 vdd.t2188 7.146
R43366 vdd.n3399 vdd.t2262 7.146
R43367 vdd.n3399 vdd.t2608 7.146
R43368 vdd.n3398 vdd.t1206 7.146
R43369 vdd.n3398 vdd.t1115 7.146
R43370 vdd.n3397 vdd.t1139 7.146
R43371 vdd.n3397 vdd.t1492 7.146
R43372 vdd.n3396 vdd.t2325 7.146
R43373 vdd.n3396 vdd.t1735 7.146
R43374 vdd.n3395 vdd.t1198 7.146
R43375 vdd.n3395 vdd.t613 7.146
R43376 vdd.n3394 vdd.t75 7.146
R43377 vdd.n3394 vdd.t2454 7.146
R43378 vdd.n3393 vdd.t554 7.146
R43379 vdd.n3393 vdd.t2936 7.146
R43380 vdd.n3392 vdd.t2395 7.146
R43381 vdd.n3392 vdd.t1791 7.146
R43382 vdd.n3391 vdd.t2160 7.146
R43383 vdd.n3391 vdd.t1556 7.146
R43384 vdd.n3390 vdd.t1747 7.146
R43385 vdd.n3390 vdd.t1132 7.146
R43386 vdd.n3599 vdd.t2605 7.146
R43387 vdd.n3599 vdd.t1729 7.146
R43388 vdd.n3588 vdd.t2838 7.146
R43389 vdd.n3588 vdd.t1966 7.146
R43390 vdd.n3587 vdd.t2331 7.146
R43391 vdd.n3587 vdd.t2665 7.146
R43392 vdd.n3586 vdd.t2594 7.146
R43393 vdd.n3586 vdd.t2915 7.146
R43394 vdd.n3585 vdd.t742 7.146
R43395 vdd.n3585 vdd.t1039 7.146
R43396 vdd.n3584 vdd.t1130 7.146
R43397 vdd.n3584 vdd.t1453 7.146
R43398 vdd.n3583 vdd.t1382 7.146
R43399 vdd.n3583 vdd.t1702 7.146
R43400 vdd.n3582 vdd.t2509 7.146
R43401 vdd.n3582 vdd.t2837 7.146
R43402 vdd.n3581 vdd.t2052 7.146
R43403 vdd.n3581 vdd.t2354 7.146
R43404 vdd.n3580 vdd.t194 7.146
R43405 vdd.n3580 vdd.t508 7.146
R43406 vdd.n3579 vdd.t610 7.146
R43407 vdd.n3579 vdd.t906 7.146
R43408 vdd.n3578 vdd.t473 7.146
R43409 vdd.n3578 vdd.t2731 7.146
R43410 vdd.n3577 vdd.t2485 7.146
R43411 vdd.n3577 vdd.t2811 7.146
R43412 vdd.n3576 vdd.t1407 7.146
R43413 vdd.n3576 vdd.t562 7.146
R43414 vdd.n3575 vdd.t297 7.146
R43415 vdd.n3575 vdd.t2400 7.146
R43416 vdd.n3574 vdd.t2138 7.146
R43417 vdd.n3574 vdd.t1266 7.146
R43418 vdd.n3573 vdd.t2618 7.146
R43419 vdd.n3573 vdd.t1751 7.146
R43420 vdd.n3572 vdd.t1474 7.146
R43421 vdd.n3572 vdd.t622 7.146
R43422 vdd.n3571 vdd.t1237 7.146
R43423 vdd.n3571 vdd.t387 7.146
R43424 vdd.n3570 vdd.t827 7.146
R43425 vdd.n3570 vdd.t2956 7.146
R43426 vdd.n3779 vdd.t145 7.146
R43427 vdd.n3779 vdd.t221 7.146
R43428 vdd.n3768 vdd.t388 7.146
R43429 vdd.n3768 vdd.t462 7.146
R43430 vdd.n3767 vdd.t980 7.146
R43431 vdd.n3767 vdd.t1997 7.146
R43432 vdd.n3766 vdd.t1240 7.146
R43433 vdd.n3766 vdd.t2251 7.146
R43434 vdd.n3765 vdd.t2367 7.146
R43435 vdd.n3765 vdd.t397 7.146
R43436 vdd.n3764 vdd.t2789 7.146
R43437 vdd.n3764 vdd.t806 7.146
R43438 vdd.n3763 vdd.t40 7.146
R43439 vdd.n3763 vdd.t1026 7.146
R43440 vdd.n3762 vdd.t1162 7.146
R43441 vdd.n3762 vdd.t2175 7.146
R43442 vdd.n3761 vdd.t716 7.146
R43443 vdd.n3761 vdd.t1693 7.146
R43444 vdd.n3760 vdd.t1822 7.146
R43445 vdd.n3760 vdd.t2830 7.146
R43446 vdd.n3759 vdd.t2258 7.146
R43447 vdd.n3759 vdd.t270 7.146
R43448 vdd.n3758 vdd.t1050 7.146
R43449 vdd.n3758 vdd.t578 7.146
R43450 vdd.n3757 vdd.t1136 7.146
R43451 vdd.n3757 vdd.t2146 7.146
R43452 vdd.n3756 vdd.t1939 7.146
R43453 vdd.n3756 vdd.t2027 7.146
R43454 vdd.n3755 vdd.t814 7.146
R43455 vdd.n3755 vdd.t880 7.146
R43456 vdd.n3754 vdd.t2679 7.146
R43457 vdd.n3754 vdd.t2754 7.146
R43458 vdd.n3753 vdd.t166 7.146
R43459 vdd.n3753 vdd.t244 7.146
R43460 vdd.n3752 vdd.t2012 7.146
R43461 vdd.n3752 vdd.t2095 7.146
R43462 vdd.n3751 vdd.t1767 7.146
R43463 vdd.n3751 vdd.t1832 7.146
R43464 vdd.n3750 vdd.t1347 7.146
R43465 vdd.n3750 vdd.t1419 7.146
R43466 vdd.n3959 vdd.t1933 7.146
R43467 vdd.n3959 vdd.t1750 7.146
R43468 vdd.n3948 vdd.t2186 7.146
R43469 vdd.n3948 vdd.t1989 7.146
R43470 vdd.n3947 vdd.t2306 7.146
R43471 vdd.n3947 vdd.t2907 7.146
R43472 vdd.n3946 vdd.t2559 7.146
R43473 vdd.n3946 vdd.t159 7.146
R43474 vdd.n3945 vdd.t709 7.146
R43475 vdd.n3945 vdd.t1267 7.146
R43476 vdd.n3944 vdd.t1105 7.146
R43477 vdd.n3944 vdd.t1692 7.146
R43478 vdd.n3943 vdd.t1346 7.146
R43479 vdd.n3943 vdd.t1931 7.146
R43480 vdd.n3942 vdd.t2477 7.146
R43481 vdd.n3942 vdd.t87 7.146
R43482 vdd.n3941 vdd.t2016 7.146
R43483 vdd.n3941 vdd.t2604 7.146
R43484 vdd.n3940 vdd.t167 7.146
R43485 vdd.n3940 vdd.t754 7.146
R43486 vdd.n3939 vdd.t581 7.146
R43487 vdd.n3939 vdd.t1137 7.146
R43488 vdd.n3938 vdd.t2651 7.146
R43489 vdd.n3938 vdd.t1923 7.146
R43490 vdd.n3937 vdd.t2457 7.146
R43491 vdd.n3937 vdd.t55 7.146
R43492 vdd.n3936 vdd.t773 7.146
R43493 vdd.n3936 vdd.t582 7.146
R43494 vdd.n3935 vdd.t2617 7.146
R43495 vdd.n3935 vdd.t2417 7.146
R43496 vdd.n3934 vdd.t1473 7.146
R43497 vdd.n3934 vdd.t1278 7.146
R43498 vdd.n3933 vdd.t1951 7.146
R43499 vdd.n3933 vdd.t1769 7.146
R43500 vdd.n3932 vdd.t829 7.146
R43501 vdd.n3932 vdd.t637 7.146
R43502 vdd.n3931 vdd.t598 7.146
R43503 vdd.n3931 vdd.t408 7.146
R43504 vdd.n3930 vdd.t180 7.146
R43505 vdd.n3930 vdd.t2970 7.146
R43506 vdd.n4139 vdd.t1766 7.146
R43507 vdd.n4139 vdd.t2801 7.146
R43508 vdd.n4128 vdd.t2015 7.146
R43509 vdd.n4128 vdd.t58 7.146
R43510 vdd.n4127 vdd.t2882 7.146
R43511 vdd.n4127 vdd.t1988 7.146
R43512 vdd.n4126 vdd.t134 7.146
R43513 vdd.n4126 vdd.t2243 7.146
R43514 vdd.n4125 vdd.t1251 7.146
R43515 vdd.n4125 vdd.t390 7.146
R43516 vdd.n4124 vdd.t1661 7.146
R43517 vdd.n4124 vdd.t801 7.146
R43518 vdd.n4123 vdd.t1917 7.146
R43519 vdd.n4123 vdd.t1021 7.146
R43520 vdd.n4122 vdd.t61 7.146
R43521 vdd.n4122 vdd.t2168 7.146
R43522 vdd.n4121 vdd.t2587 7.146
R43523 vdd.n4121 vdd.t1685 7.146
R43524 vdd.n4120 vdd.t732 7.146
R43525 vdd.n4120 vdd.t2823 7.146
R43526 vdd.n4119 vdd.t1120 7.146
R43527 vdd.n4119 vdd.t264 7.146
R43528 vdd.n4118 vdd.t2033 7.146
R43529 vdd.n4118 vdd.t422 7.146
R43530 vdd.n4117 vdd.t30 7.146
R43531 vdd.n4117 vdd.t2142 7.146
R43532 vdd.n4116 vdd.t602 7.146
R43533 vdd.n4116 vdd.t1616 7.146
R43534 vdd.n4115 vdd.t2441 7.146
R43535 vdd.n4115 vdd.t495 7.146
R43536 vdd.n4114 vdd.t1303 7.146
R43537 vdd.n4114 vdd.t2343 7.146
R43538 vdd.n4113 vdd.t1784 7.146
R43539 vdd.n4113 vdd.t2824 7.146
R43540 vdd.n4112 vdd.t657 7.146
R43541 vdd.n4112 vdd.t1687 7.146
R43542 vdd.n4111 vdd.t428 7.146
R43543 vdd.n4111 vdd.t1439 7.146
R43544 vdd.n4110 vdd.t2991 7.146
R43545 vdd.n4110 vdd.t1022 7.146
R43546 vdd.n4319 vdd.t263 7.146
R43547 vdd.n4319 vdd.t1611 7.146
R43548 vdd.n4308 vdd.t493 7.146
R43549 vdd.n4308 vdd.t1855 7.146
R43550 vdd.n4307 vdd.t2219 7.146
R43551 vdd.n4307 vdd.t320 7.146
R43552 vdd.n4306 vdd.t2447 7.146
R43553 vdd.n4306 vdd.t570 7.146
R43554 vdd.n4305 vdd.t605 7.146
R43555 vdd.n4305 vdd.t1681 7.146
R43556 vdd.n4304 vdd.t993 7.146
R43557 vdd.n4304 vdd.t2105 7.146
R43558 vdd.n4303 vdd.t1247 7.146
R43559 vdd.n4303 vdd.t2339 7.146
R43560 vdd.n4302 vdd.t2374 7.146
R43561 vdd.n4302 vdd.t487 7.146
R43562 vdd.n4301 vdd.t1911 7.146
R43563 vdd.n4301 vdd.t7 7.146
R43564 vdd.n4300 vdd.t50 7.146
R43565 vdd.n4300 vdd.t1133 7.146
R43566 vdd.n4299 vdd.t469 7.146
R43567 vdd.n4299 vdd.t1561 7.146
R43568 vdd.n4298 vdd.t2876 7.146
R43569 vdd.n4298 vdd.t2003 7.146
R43570 vdd.n4297 vdd.t2348 7.146
R43571 vdd.n4297 vdd.t465 7.146
R43572 vdd.n4296 vdd.t2068 7.146
R43573 vdd.n4296 vdd.t452 7.146
R43574 vdd.n4295 vdd.t914 7.146
R43575 vdd.n4295 vdd.t2298 7.146
R43576 vdd.n4294 vdd.t2783 7.146
R43577 vdd.n4294 vdd.t1152 7.146
R43578 vdd.n4293 vdd.t285 7.146
R43579 vdd.n4293 vdd.t1635 7.146
R43580 vdd.n4292 vdd.t2122 7.146
R43581 vdd.n4292 vdd.t515 7.146
R43582 vdd.n4291 vdd.t1880 7.146
R43583 vdd.n4291 vdd.t280 7.146
R43584 vdd.n4290 vdd.t1456 7.146
R43585 vdd.n4290 vdd.t2843 7.146
R43586 vdd.n4499 vdd.t1285 7.146
R43587 vdd.n4499 vdd.t1443 7.146
R43588 vdd.n4488 vdd.t1540 7.146
R43589 vdd.n4488 vdd.t1691 7.146
R43590 vdd.n4487 vdd.t1284 7.146
R43591 vdd.n4487 vdd.t867 7.146
R43592 vdd.n4486 vdd.t1539 7.146
R43593 vdd.n4486 vdd.t1113 7.146
R43594 vdd.n4485 vdd.t2691 7.146
R43595 vdd.n4485 vdd.t2261 7.146
R43596 vdd.n4484 vdd.t113 7.146
R43597 vdd.n4484 vdd.t2675 7.146
R43598 vdd.n4483 vdd.t354 7.146
R43599 vdd.n4483 vdd.t2918 7.146
R43600 vdd.n4482 vdd.t1469 7.146
R43601 vdd.n4482 vdd.t1043 7.146
R43602 vdd.n4481 vdd.t989 7.146
R43603 vdd.n4481 vdd.t589 7.146
R43604 vdd.n4480 vdd.t2134 7.146
R43605 vdd.n4480 vdd.t1705 7.146
R43606 vdd.n4479 vdd.t2556 7.146
R43607 vdd.n4479 vdd.t2118 7.146
R43608 vdd.n4478 vdd.t1345 7.146
R43609 vdd.n4478 vdd.t1379 7.146
R43610 vdd.n4477 vdd.t1445 7.146
R43611 vdd.n4477 vdd.t1012 7.146
R43612 vdd.n4476 vdd.t133 7.146
R43613 vdd.n4476 vdd.t288 7.146
R43614 vdd.n4475 vdd.t1977 7.146
R43615 vdd.n4475 vdd.t2125 7.146
R43616 vdd.n4474 vdd.t842 7.146
R43617 vdd.n4474 vdd.t979 7.146
R43618 vdd.n4473 vdd.t1313 7.146
R43619 vdd.n4473 vdd.t1459 7.146
R43620 vdd.n4472 vdd.t205 7.146
R43621 vdd.n4472 vdd.t345 7.146
R43622 vdd.n4471 vdd.t2942 7.146
R43623 vdd.n4471 vdd.t106 7.146
R43624 vdd.n4470 vdd.t2520 7.146
R43625 vdd.n4470 vdd.t2686 7.146
R43626 vdd.n4679 vdd.t1124 7.146
R43627 vdd.n4679 vdd.t283 7.146
R43628 vdd.n4668 vdd.t1378 7.146
R43629 vdd.n4668 vdd.t517 7.146
R43630 vdd.n4667 vdd.t1860 7.146
R43631 vdd.n4667 vdd.t2195 7.146
R43632 vdd.n4666 vdd.t2110 7.146
R43633 vdd.n4666 vdd.t2423 7.146
R43634 vdd.n4665 vdd.t266 7.146
R43635 vdd.n4665 vdd.t585 7.146
R43636 vdd.n4664 vdd.t671 7.146
R43637 vdd.n4664 vdd.t966 7.146
R43638 vdd.n4663 vdd.t899 7.146
R43639 vdd.n4663 vdd.t1221 7.146
R43640 vdd.n4662 vdd.t2051 7.146
R43641 vdd.n4662 vdd.t2353 7.146
R43642 vdd.n4661 vdd.t1566 7.146
R43643 vdd.n4661 vdd.t1884 7.146
R43644 vdd.n4660 vdd.t2716 7.146
R43645 vdd.n4660 vdd.t26 7.146
R43646 vdd.n4659 vdd.t131 7.146
R43647 vdd.n4659 vdd.t453 7.146
R43648 vdd.n4658 vdd.t750 7.146
R43649 vdd.n4658 vdd.t2972 7.146
R43650 vdd.n4657 vdd.t2024 7.146
R43651 vdd.n4657 vdd.t2323 7.146
R43652 vdd.n4656 vdd.t2948 7.146
R43653 vdd.n4656 vdd.t2086 7.146
R43654 vdd.n4655 vdd.t1800 7.146
R43655 vdd.n4655 vdd.t931 7.146
R43656 vdd.n4654 vdd.t687 7.146
R43657 vdd.n4654 vdd.t2800 7.146
R43658 vdd.n4653 vdd.t1138 7.146
R43659 vdd.n4653 vdd.t299 7.146
R43660 vdd.n4652 vdd.t17 7.146
R43661 vdd.n4652 vdd.t2144 7.146
R43662 vdd.n4651 vdd.t2776 7.146
R43663 vdd.n4651 vdd.t1906 7.146
R43664 vdd.n4650 vdd.t2345 7.146
R43665 vdd.n4650 vdd.t1479 7.146
R43666 vdd.n4859 vdd.t2941 7.146
R43667 vdd.n4859 vdd.t2082 7.146
R43668 vdd.n4848 vdd.t204 7.146
R43669 vdd.n4848 vdd.t2312 7.146
R43670 vdd.n4847 vdd.t200 7.146
R43671 vdd.n4847 vdd.t513 7.146
R43672 vdd.n4846 vdd.t444 7.146
R43673 vdd.n4846 vdd.t768 7.146
R43674 vdd.n4845 vdd.t1564 7.146
R43675 vdd.n4845 vdd.t1879 7.146
R43676 vdd.n4844 vdd.t1973 7.146
R43677 vdd.n4844 vdd.t2296 7.146
R43678 vdd.n4843 vdd.t2232 7.146
R43679 vdd.n4843 vdd.t2543 7.146
R43680 vdd.n4842 vdd.t373 7.146
R43681 vdd.n4842 vdd.t697 7.146
R43682 vdd.n4841 vdd.t2892 7.146
R43683 vdd.n4841 vdd.t218 7.146
R43684 vdd.n4840 vdd.t1006 7.146
R43685 vdd.n4840 vdd.t1332 7.146
R43686 vdd.n4839 vdd.t1425 7.146
R43687 vdd.n4839 vdd.t1756 7.146
R43688 vdd.n4838 vdd.t2317 7.146
R43689 vdd.n4838 vdd.t1574 7.146
R43690 vdd.n4837 vdd.t342 7.146
R43691 vdd.n4837 vdd.t660 7.146
R43692 vdd.n4836 vdd.t1760 7.146
R43693 vdd.n4836 vdd.t888 7.146
R43694 vdd.n4835 vdd.t630 7.146
R43695 vdd.n4835 vdd.t2763 7.146
R43696 vdd.n4834 vdd.t2476 7.146
R43697 vdd.n4834 vdd.t1610 7.146
R43698 vdd.n4833 vdd.t2960 7.146
R43699 vdd.n4833 vdd.t2098 7.146
R43700 vdd.n4832 vdd.t1819 7.146
R43701 vdd.n4832 vdd.t946 7.146
R43702 vdd.n4831 vdd.t1584 7.146
R43703 vdd.n4831 vdd.t734 7.146
R43704 vdd.n4830 vdd.t1156 7.146
R43705 vdd.n4830 vdd.t310 7.146
R43706 vdd.n5039 vdd.t1755 7.146
R43707 vdd.n5039 vdd.t821 7.146
R43708 vdd.n5028 vdd.t1998 7.146
R43709 vdd.n5028 vdd.t1056 7.146
R43710 vdd.n5027 vdd.t1490 7.146
R43711 vdd.n5027 vdd.t2864 7.146
R43712 vdd.n5026 vdd.t1743 7.146
R43713 vdd.n5026 vdd.t120 7.146
R43714 vdd.n5025 vdd.t2887 7.146
R43715 vdd.n5025 vdd.t1239 7.146
R43716 vdd.n5024 vdd.t308 7.146
R43717 vdd.n5024 vdd.t1646 7.146
R43718 vdd.n5023 vdd.t551 7.146
R43719 vdd.n5023 vdd.t1902 7.146
R43720 vdd.n5022 vdd.t1667 7.146
R43721 vdd.n5022 vdd.t39 7.146
R43722 vdd.n5021 vdd.t1191 7.146
R43723 vdd.n5021 vdd.t2570 7.146
R43724 vdd.n5020 vdd.t2321 7.146
R43725 vdd.n5020 vdd.t715 7.146
R43726 vdd.n5019 vdd.t2757 7.146
R43727 vdd.n5019 vdd.t1110 7.146
R43728 vdd.n5018 vdd.t919 7.146
R43729 vdd.n5018 vdd.t99 7.146
R43730 vdd.n5017 vdd.t1640 7.146
R43731 vdd.n5017 vdd.t13 7.146
R43732 vdd.n5016 vdd.t593 7.146
R43733 vdd.n5016 vdd.t2632 7.146
R43734 vdd.n5015 vdd.t2428 7.146
R43735 vdd.n5015 vdd.t1482 7.146
R43736 vdd.n5014 vdd.t1281 7.146
R43737 vdd.n5014 vdd.t371 7.146
R43738 vdd.n5013 vdd.t1773 7.146
R43739 vdd.n5013 vdd.t834 7.146
R43740 vdd.n5012 vdd.t645 7.146
R43741 vdd.n5012 vdd.t2712 7.146
R43742 vdd.n5011 vdd.t416 7.146
R43743 vdd.n5011 vdd.t2446 7.146
R43744 vdd.n5010 vdd.t2975 7.146
R43745 vdd.n5010 vdd.t2044 7.146
R43746 vdd.n5219 vdd.t584 7.146
R43747 vdd.n5219 vdd.t2625 7.146
R43748 vdd.n5208 vdd.t820 7.146
R43749 vdd.n5208 vdd.t2874 7.146
R43750 vdd.n5207 vdd.t2810 7.146
R43751 vdd.n5207 vdd.t1168 7.146
R43752 vdd.n5206 vdd.t67 7.146
R43753 vdd.n5206 vdd.t1413 7.146
R43754 vdd.n5205 vdd.t1185 7.146
R43755 vdd.n5205 vdd.t2558 7.146
R43756 vdd.n5204 vdd.t1601 7.146
R43757 vdd.n5204 vdd.t2969 7.146
R43758 vdd.n5203 vdd.t1841 7.146
R43759 vdd.n5203 vdd.t236 7.146
R43760 vdd.n5202 vdd.t2988 7.146
R43761 vdd.n5202 vdd.t1350 7.146
R43762 vdd.n5201 vdd.t2504 7.146
R43763 vdd.n5201 vdd.t872 7.146
R43764 vdd.n5200 vdd.t655 7.146
R43765 vdd.n5200 vdd.t2014 7.146
R43766 vdd.n5199 vdd.t1067 7.146
R43767 vdd.n5199 vdd.t2416 7.146
R43768 vdd.n5198 vdd.t2521 7.146
R43769 vdd.n5198 vdd.t1671 7.146
R43770 vdd.n5197 vdd.t2962 7.146
R43771 vdd.n5197 vdd.t1318 7.146
R43772 vdd.n5196 vdd.t2373 7.146
R43773 vdd.n5196 vdd.t1432 7.146
R43774 vdd.n5195 vdd.t1246 7.146
R43775 vdd.n5195 vdd.t316 7.146
R43776 vdd.n5194 vdd.t126 7.146
R43777 vdd.n5194 vdd.t2167 7.146
R43778 vdd.n5193 vdd.t604 7.146
R43779 vdd.n5193 vdd.t2647 7.146
R43780 vdd.n5192 vdd.t2445 7.146
R43781 vdd.n5192 vdd.t1501 7.146
R43782 vdd.n5191 vdd.t2216 7.146
R43783 vdd.n5191 vdd.t1259 7.146
R43784 vdd.n5190 vdd.t1785 7.146
R43785 vdd.n5190 vdd.t845 7.146
R43786 vdd.n5399 vdd.t2645 7.146
R43787 vdd.n5399 vdd.t1428 7.146
R43788 vdd.n5388 vdd.t2898 7.146
R43789 vdd.n5388 vdd.t1674 7.146
R43790 vdd.n5387 vdd.t1141 7.146
R43791 vdd.n5387 vdd.t2484 7.146
R43792 vdd.n5386 vdd.t1395 7.146
R43793 vdd.n5386 vdd.t2749 7.146
R43794 vdd.n5385 vdd.t2530 7.146
R43795 vdd.n5385 vdd.t871 7.146
R43796 vdd.n5384 vdd.t2952 7.146
R43797 vdd.n5384 vdd.t1275 7.146
R43798 vdd.n5383 vdd.t210 7.146
R43799 vdd.n5383 vdd.t1526 7.146
R43800 vdd.n5382 vdd.t1324 7.146
R43801 vdd.n5382 vdd.t2676 7.146
R43802 vdd.n5381 vdd.t853 7.146
R43803 vdd.n5381 vdd.t2201 7.146
R43804 vdd.n5380 vdd.t1984 7.146
R43805 vdd.n5380 vdd.t338 7.146
R43806 vdd.n5379 vdd.t2397 7.146
R43807 vdd.n5379 vdd.t764 7.146
R43808 vdd.n5378 vdd.t1780 7.146
R43809 vdd.n5378 vdd.t296 7.146
R43810 vdd.n5377 vdd.t1292 7.146
R43811 vdd.n5377 vdd.t2646 7.146
R43812 vdd.n5376 vdd.t1452 7.146
R43813 vdd.n5376 vdd.t274 7.146
R43814 vdd.n5375 vdd.t334 7.146
R43815 vdd.n5375 vdd.t2114 7.146
R43816 vdd.n5374 vdd.t2194 7.146
R43817 vdd.n5374 vdd.t963 7.146
R43818 vdd.n5373 vdd.t2668 7.146
R43819 vdd.n5373 vdd.t1449 7.146
R43820 vdd.n5372 vdd.t1520 7.146
R43821 vdd.n5372 vdd.t330 7.146
R43822 vdd.n5371 vdd.t1273 7.146
R43823 vdd.n5371 vdd.t94 7.146
R43824 vdd.n5370 vdd.t865 7.146
R43825 vdd.n5370 vdd.t2660 7.146
R43826 vdd.n5579 vdd.t1448 7.146
R43827 vdd.n5579 vdd.t269 7.146
R43828 vdd.n5568 vdd.t1698 7.146
R43829 vdd.n5568 vdd.t498 7.146
R43830 vdd.n5567 vdd.t2465 7.146
R43831 vdd.n5567 vdd.t816 7.146
R43832 vdd.n5566 vdd.t2727 7.146
R43833 vdd.n5566 vdd.t1051 7.146
R43834 vdd.n5565 vdd.t848 7.146
R43835 vdd.n5565 vdd.t2197 7.146
R43836 vdd.n5564 vdd.t1262 7.146
R43837 vdd.n5564 vdd.t2611 7.146
R43838 vdd.n5563 vdd.t1502 7.146
R43839 vdd.n5563 vdd.t2846 7.146
R43840 vdd.n5562 vdd.t2649 7.146
R43841 vdd.n5562 vdd.t968 7.146
R43842 vdd.n5561 vdd.t2170 7.146
R43843 vdd.n5561 vdd.t519 7.146
R43844 vdd.n5560 vdd.t318 7.146
R43845 vdd.n5560 vdd.t1636 7.146
R43846 vdd.n5559 vdd.t741 7.146
R43847 vdd.n5559 vdd.t2070 7.146
R43848 vdd.n5558 vdd.t402 7.146
R43849 vdd.n5558 vdd.t1874 7.146
R43850 vdd.n5557 vdd.t2622 7.146
R43851 vdd.n5557 vdd.t948 7.146
R43852 vdd.n5556 vdd.t293 7.146
R43853 vdd.n5556 vdd.t2073 7.146
R43854 vdd.n5555 vdd.t2130 7.146
R43855 vdd.n5555 vdd.t921 7.146
R43856 vdd.n5554 vdd.t985 7.146
R43857 vdd.n5554 vdd.t2788 7.146
R43858 vdd.n5553 vdd.t1465 7.146
R43859 vdd.n5553 vdd.t291 7.146
R43860 vdd.n5552 vdd.t350 7.146
R43861 vdd.n5552 vdd.t2128 7.146
R43862 vdd.n5551 vdd.t111 7.146
R43863 vdd.n5551 vdd.t1889 7.146
R43864 vdd.n5550 vdd.t2690 7.146
R43865 vdd.n5550 vdd.t1462 7.146
R43866 vdd.n5759 vdd.t2929 7.146
R43867 vdd.n5759 vdd.t93 7.146
R43868 vdd.n5748 vdd.t188 7.146
R43869 vdd.n5748 vdd.t329 7.146
R43870 vdd.n5747 vdd.t1795 7.146
R43871 vdd.n5747 vdd.t1373 7.146
R43872 vdd.n5746 vdd.t2059 7.146
R43873 vdd.n5746 vdd.t1606 7.146
R43874 vdd.n5745 vdd.t201 7.146
R43875 vdd.n5745 vdd.t2762 7.146
R43876 vdd.n5744 vdd.t615 7.146
R43877 vdd.n5744 vdd.t186 7.146
R43878 vdd.n5743 vdd.t841 7.146
R43879 vdd.n5743 vdd.t431 7.146
R43880 vdd.n5742 vdd.t1976 7.146
R43881 vdd.n5742 vdd.t1546 7.146
R43882 vdd.n5741 vdd.t1497 7.146
R43883 vdd.n5741 vdd.t1073 7.146
R43884 vdd.n5740 vdd.t2641 7.146
R43885 vdd.n5740 vdd.t2215 7.146
R43886 vdd.n5739 vdd.t64 7.146
R43887 vdd.n5739 vdd.t2624 7.146
R43888 vdd.n5738 vdd.t1225 7.146
R43889 vdd.n5738 vdd.t1249 7.146
R43890 vdd.n5737 vdd.t1948 7.146
R43891 vdd.n5737 vdd.t1514 7.146
R43892 vdd.n5736 vdd.t1746 7.146
R43893 vdd.n5736 vdd.t1893 7.146
R43894 vdd.n5735 vdd.t619 7.146
R43895 vdd.n5735 vdd.t774 7.146
R43896 vdd.n5734 vdd.t2466 7.146
R43897 vdd.n5734 vdd.t2621 7.146
R43898 vdd.n5733 vdd.t2951 7.146
R43899 vdd.n5733 vdd.t112 7.146
R43900 vdd.n5732 vdd.t1801 7.146
R43901 vdd.n5732 vdd.t1952 7.146
R43902 vdd.n5731 vdd.t1571 7.146
R43903 vdd.n5731 vdd.t1718 7.146
R43904 vdd.n5730 vdd.t1140 7.146
R43905 vdd.n5730 vdd.t1283 7.146
R43906 vdd.n5939 vdd.t1464 7.146
R43907 vdd.n5939 vdd.t2853 7.146
R43908 vdd.n5928 vdd.t1719 7.146
R43909 vdd.n5928 vdd.t110 7.146
R43910 vdd.n5927 vdd.t2722 7.146
R43911 vdd.n5927 vdd.t812 7.146
R43912 vdd.n5926 vdd.t2950 7.146
R43913 vdd.n5926 vdd.t1042 7.146
R43914 vdd.n5925 vdd.t1088 7.146
R43915 vdd.n5925 vdd.t2187 7.146
R43916 vdd.n5924 vdd.t1495 7.146
R43917 vdd.n5924 vdd.t2607 7.146
R43918 vdd.n5923 vdd.t1745 7.146
R43919 vdd.n5923 vdd.t2842 7.146
R43920 vdd.n5922 vdd.t2891 7.146
R43921 vdd.n5922 vdd.t962 7.146
R43922 vdd.n5921 vdd.t2393 7.146
R43923 vdd.n5921 vdd.t514 7.146
R43924 vdd.n5920 vdd.t553 7.146
R43925 vdd.n5920 vdd.t1634 7.146
R43926 vdd.n5919 vdd.t945 7.146
R43927 vdd.n5919 vdd.t2064 7.146
R43928 vdd.n5918 vdd.t2597 7.146
R43929 vdd.n5918 vdd.t1714 7.146
R43930 vdd.n5917 vdd.t2858 7.146
R43931 vdd.n5917 vdd.t944 7.146
R43932 vdd.n5916 vdd.t306 7.146
R43933 vdd.n5916 vdd.t1660 7.146
R43934 vdd.n5915 vdd.t2155 7.146
R43935 vdd.n5915 vdd.t544 7.146
R43936 vdd.n5914 vdd.t1008 7.146
R43937 vdd.n5914 vdd.t2387 7.146
R43938 vdd.n5913 vdd.t1489 7.146
R43939 vdd.n5913 vdd.t2877 7.146
R43940 vdd.n5912 vdd.t379 7.146
R43941 vdd.n5912 vdd.t1737 7.146
R43942 vdd.n5911 vdd.t130 7.146
R43943 vdd.n5911 vdd.t1483 7.146
R43944 vdd.n5910 vdd.t2715 7.146
R43945 vdd.n5910 vdd.t1079 7.146
R43946 vdd.n6119 vdd.t302 7.146
R43947 vdd.n6119 vdd.t1655 7.146
R43948 vdd.n6108 vdd.t541 7.146
R43949 vdd.n6108 vdd.t1912 7.146
R43950 vdd.n6107 vdd.t1011 7.146
R43951 vdd.n6107 vdd.t2116 7.146
R43952 vdd.n6106 vdd.t1258 7.146
R43953 vdd.n6106 vdd.t2352 7.146
R43954 vdd.n6105 vdd.t2392 7.146
R43955 vdd.n6105 vdd.t507 7.146
R43956 vdd.n6104 vdd.t2814 7.146
R43957 vdd.n6104 vdd.t905 7.146
R43958 vdd.n6103 vdd.t72 7.146
R43959 vdd.n6103 vdd.t1148 7.146
R43960 vdd.n6102 vdd.t1190 7.146
R43961 vdd.n6102 vdd.t2293 7.146
R43962 vdd.n6101 vdd.t740 7.146
R43963 vdd.n6101 vdd.t1810 7.146
R43964 vdd.n6100 vdd.t1847 7.146
R43965 vdd.n6100 vdd.t2957 7.146
R43966 vdd.n6099 vdd.t2275 7.146
R43967 vdd.n6099 vdd.t389 7.146
R43968 vdd.n6098 vdd.t1180 7.146
R43969 vdd.n6098 vdd.t327 7.146
R43970 vdd.n6097 vdd.t1160 7.146
R43971 vdd.n6097 vdd.t2273 7.146
R43972 vdd.n6096 vdd.t2106 7.146
R43973 vdd.n6096 vdd.t486 7.146
R43974 vdd.n6095 vdd.t954 7.146
R43975 vdd.n6095 vdd.t2335 7.146
R43976 vdd.n6094 vdd.t2827 7.146
R43977 vdd.n6094 vdd.t1205 7.146
R43978 vdd.n6093 vdd.t321 7.146
R43979 vdd.n6093 vdd.t1680 7.146
R43980 vdd.n6092 vdd.t2174 7.146
R43981 vdd.n6092 vdd.t569 7.146
R43982 vdd.n6091 vdd.t1926 7.146
R43983 vdd.n6091 vdd.t317 7.146
R43984 vdd.n6090 vdd.t1503 7.146
R43985 vdd.n6090 vdd.t2901 7.146
R43986 vdd.n6299 vdd.t1341 7.146
R43987 vdd.n6299 vdd.t1487 7.146
R43988 vdd.n6288 vdd.t1588 7.146
R43989 vdd.n6288 vdd.t1739 7.146
R43990 vdd.n6287 vdd.t129 7.146
R43991 vdd.n6287 vdd.t2696 7.146
R43992 vdd.n6286 vdd.t376 7.146
R43993 vdd.n6286 vdd.t2928 7.146
R43994 vdd.n6285 vdd.t1486 7.146
R43995 vdd.n6285 vdd.t1063 7.146
R43996 vdd.n6284 vdd.t1914 7.146
R43997 vdd.n6284 vdd.t1468 7.146
R43998 vdd.n6283 vdd.t2154 7.146
R43999 vdd.n6283 vdd.t1721 7.146
R44000 vdd.n6282 vdd.t304 7.146
R44001 vdd.n6282 vdd.t2860 7.146
R44002 vdd.n6281 vdd.t2809 7.146
R44003 vdd.n6281 vdd.t2370 7.146
R44004 vdd.n6280 vdd.t939 7.146
R44005 vdd.n6280 vdd.t525 7.146
R44006 vdd.n6279 vdd.t1366 7.146
R44007 vdd.n6279 vdd.t925 7.146
R44008 vdd.n6278 vdd.t2674 7.146
R44009 vdd.n6278 vdd.t2710 7.146
R44010 vdd.n6277 vdd.t287 7.146
R44011 vdd.n6277 vdd.t2831 7.146
R44012 vdd.n6276 vdd.t179 7.146
R44013 vdd.n6276 vdd.t324 7.146
R44014 vdd.n6275 vdd.t2035 7.146
R44015 vdd.n6275 vdd.t2181 7.146
R44016 vdd.n6274 vdd.t887 7.146
R44017 vdd.n6274 vdd.t1033 7.146
R44018 vdd.n6273 vdd.t1368 7.146
R44019 vdd.n6273 vdd.t1509 7.146
R44020 vdd.n6272 vdd.t253 7.146
R44021 vdd.n6272 vdd.t401 7.146
R44022 vdd.n6271 vdd.t2985 7.146
R44023 vdd.n6271 vdd.t157 7.146
R44024 vdd.n6270 vdd.t2583 7.146
R44025 vdd.n6270 vdd.t2736 7.146
R44026 vdd.n6479 vdd.t1167 7.146
R44027 vdd.n6479 vdd.t2965 7.146
R44028 vdd.n6468 vdd.t1412 7.146
R44029 vdd.n6468 vdd.t229 7.146
R44030 vdd.n6467 vdd.t695 7.146
R44031 vdd.n6467 vdd.t2021 7.146
R44032 vdd.n6466 vdd.t912 7.146
R44033 vdd.n6466 vdd.t2266 7.146
R44034 vdd.n6465 vdd.t2065 7.146
R44035 vdd.n6465 vdd.t415 7.146
R44036 vdd.n6464 vdd.t2470 7.146
R44037 vdd.n6464 vdd.t819 7.146
R44038 vdd.n6463 vdd.t2733 7.146
R44039 vdd.n6463 vdd.t1057 7.146
R44040 vdd.n6462 vdd.t852 7.146
R44041 vdd.n6462 vdd.t2203 7.146
R44042 vdd.n6461 vdd.t398 7.146
R44043 vdd.n6461 vdd.t1713 7.146
R44044 vdd.n6460 vdd.t1505 7.146
R44045 vdd.n6460 vdd.t2852 7.146
R44046 vdd.n6459 vdd.t1927 7.146
R44047 vdd.n6459 vdd.t289 7.146
R44048 vdd.n6458 vdd.t2058 7.146
R44049 vdd.n6458 vdd.t552 7.146
R44050 vdd.n6457 vdd.t833 7.146
R44051 vdd.n6457 vdd.t2166 7.146
R44052 vdd.n6456 vdd.t2990 7.146
R44053 vdd.n6456 vdd.t1782 7.146
R44054 vdd.n6455 vdd.t1845 7.146
R44055 vdd.n6455 vdd.t654 7.146
R44056 vdd.n6454 vdd.t739 7.146
R44057 vdd.n6454 vdd.t2503 7.146
R44058 vdd.n6453 vdd.t1189 7.146
R44059 vdd.n6453 vdd.t2987 7.146
R44060 vdd.n6452 vdd.t71 7.146
R44061 vdd.n6452 vdd.t1840 7.146
R44062 vdd.n6451 vdd.t2813 7.146
R44063 vdd.n6451 vdd.t1600 7.146
R44064 vdd.n6450 vdd.t2391 7.146
R44065 vdd.n6450 vdd.t1184 7.146
R44066 vdd.n6659 vdd.t2984 7.146
R44067 vdd.n6659 vdd.t1777 7.146
R44068 vdd.n6648 vdd.t252 7.146
R44069 vdd.n6648 vdd.t2032 7.146
R44070 vdd.n6647 vdd.t1991 7.146
R44071 vdd.n6647 vdd.t341 7.146
R44072 vdd.n6646 vdd.t2244 7.146
R44073 vdd.n6646 vdd.t595 7.146
R44074 vdd.n6645 vdd.t392 7.146
R44075 vdd.n6645 vdd.t1710 7.146
R44076 vdd.n6644 vdd.t804 7.146
R44077 vdd.n6644 vdd.t2124 7.146
R44078 vdd.n6643 vdd.t1025 7.146
R44079 vdd.n6643 vdd.t2364 7.146
R44080 vdd.n6642 vdd.t2172 7.146
R44081 vdd.n6642 vdd.t518 7.146
R44082 vdd.n6641 vdd.t1690 7.146
R44083 vdd.n6641 vdd.t34 7.146
R44084 vdd.n6640 vdd.t2826 7.146
R44085 vdd.n6640 vdd.t1155 7.146
R44086 vdd.n6639 vdd.t265 7.146
R44087 vdd.n6639 vdd.t1583 7.146
R44088 vdd.n6638 vdd.t649 7.146
R44089 vdd.n6638 vdd.t2133 7.146
R44090 vdd.n6637 vdd.t2143 7.146
R44091 vdd.n6637 vdd.t485 7.146
R44092 vdd.n6636 vdd.t1798 7.146
R44093 vdd.n6636 vdd.t612 7.146
R44094 vdd.n6635 vdd.t681 7.146
R44095 vdd.n6635 vdd.t2453 7.146
R44096 vdd.n6634 vdd.t2529 7.146
R44097 vdd.n6634 vdd.t1314 7.146
R44098 vdd.n6633 vdd.t10 7.146
R44099 vdd.n6633 vdd.t1794 7.146
R44100 vdd.n6632 vdd.t1866 7.146
R44101 vdd.n6632 vdd.t674 7.146
R44102 vdd.n6631 vdd.t1626 7.146
R44103 vdd.n6631 vdd.t439 7.146
R44104 vdd.n6630 vdd.t1212 7.146
R44105 vdd.n6630 vdd.t3 7.146
R44106 vdd.n6839 vdd.t1790 7.146
R44107 vdd.n6839 vdd.t856 7.146
R44108 vdd.n6828 vdd.t2057 7.146
R44109 vdd.n6828 vdd.t1103 7.146
R44110 vdd.n6827 vdd.t322 7.146
R44111 vdd.n6827 vdd.t1666 7.146
R44112 vdd.n6826 vdd.t573 7.146
R44113 vdd.n6826 vdd.t1916 7.146
R44114 vdd.n6825 vdd.t1684 7.146
R44115 vdd.n6825 vdd.t60 7.146
R44116 vdd.n6824 vdd.t2107 7.146
R44117 vdd.n6824 vdd.t474 7.146
R44118 vdd.n6823 vdd.t2340 7.146
R44119 vdd.n6823 vdd.t731 7.146
R44120 vdd.n6822 vdd.t492 7.146
R44121 vdd.n6822 vdd.t1835 7.146
R44122 vdd.n6821 vdd.t9 7.146
R44123 vdd.n6821 vdd.t1374 7.146
R44124 vdd.n6820 vdd.t1134 7.146
R44125 vdd.n6820 vdd.t2499 7.146
R44126 vdd.n6819 vdd.t1563 7.146
R44127 vdd.n6819 vdd.t2925 7.146
R44128 vdd.n6818 vdd.t2254 7.146
R44129 vdd.n6818 vdd.t1394 7.146
R44130 vdd.n6817 vdd.t468 7.146
R44131 vdd.n6817 vdd.t1816 7.146
R44132 vdd.n6816 vdd.t625 7.146
R44133 vdd.n6816 vdd.t2685 7.146
R44134 vdd.n6815 vdd.t2473 7.146
R44135 vdd.n6815 vdd.t1532 7.146
R44136 vdd.n6814 vdd.t1337 7.146
R44137 vdd.n6814 vdd.t421 7.146
R44138 vdd.n6813 vdd.t1812 7.146
R44139 vdd.n6813 vdd.t874 7.146
R44140 vdd.n6812 vdd.t706 7.146
R44141 vdd.n6812 vdd.t2752 7.146
R44142 vdd.n6811 vdd.t455 7.146
R44143 vdd.n6811 vdd.t2491 7.146
R44144 vdd.n6810 vdd.t27 7.146
R44145 vdd.n6810 vdd.t2090 7.146
R44146 vdd.n7019 vdd.t1277 7.146
R44147 vdd.n7019 vdd.t2678 7.146
R44148 vdd.n7008 vdd.t1529 7.146
R44149 vdd.n7008 vdd.t2920 7.146
R44150 vdd.n7007 vdd.t1888 7.146
R44151 vdd.n7007 vdd.t2983 7.146
R44152 vdd.n7006 vdd.t2127 7.146
R44153 vdd.n7006 vdd.t254 7.146
R44154 vdd.n7005 vdd.t290 7.146
R44155 vdd.n7005 vdd.t1369 7.146
R44156 vdd.n7004 vdd.t705 7.146
R44157 vdd.n7004 vdd.t1781 7.146
R44158 vdd.n7003 vdd.t922 7.146
R44159 vdd.n7003 vdd.t2037 7.146
R44160 vdd.n7002 vdd.t2076 7.146
R44161 vdd.n7002 vdd.t182 7.146
R44162 vdd.n7001 vdd.t1587 7.146
R44163 vdd.n7001 vdd.t2704 7.146
R44164 vdd.n7000 vdd.t2737 7.146
R44165 vdd.n7000 vdd.t830 7.146
R44166 vdd.n6999 vdd.t162 7.146
R44167 vdd.n6999 vdd.t1238 7.146
R44168 vdd.n6998 vdd.t863 7.146
R44169 vdd.n6998 vdd.t2994 7.146
R44170 vdd.n6997 vdd.t2050 7.146
R44171 vdd.n6997 vdd.t158 7.146
R44172 vdd.n6996 vdd.t124 7.146
R44173 vdd.n6996 vdd.t1478 7.146
R44174 vdd.n6995 vdd.t1961 7.146
R44175 vdd.n6995 vdd.t362 7.146
R44176 vdd.n6994 vdd.t836 7.146
R44177 vdd.n6994 vdd.t2222 7.146
R44178 vdd.n6993 vdd.t1302 7.146
R44179 vdd.n6993 vdd.t2709 7.146
R44180 vdd.n6992 vdd.t190 7.146
R44181 vdd.n6992 vdd.t1554 7.146
R44182 vdd.n6991 vdd.t2933 7.146
R44183 vdd.n6991 vdd.t1300 7.146
R44184 vdd.n6990 vdd.t2508 7.146
R44185 vdd.n6990 vdd.t892 7.146
R44186 vdd.n7199 vdd.t2342 7.146
R44187 vdd.n7199 vdd.t1472 7.146
R44188 vdd.n7188 vdd.t2602 7.146
R44189 vdd.n7188 vdd.t1726 7.146
R44190 vdd.n7187 vdd.t967 7.146
R44191 vdd.n7187 vdd.t1289 7.146
R44192 vdd.n7186 vdd.t1223 7.146
R44193 vdd.n7186 vdd.t1545 7.146
R44194 vdd.n7185 vdd.t2357 7.146
R44195 vdd.n7185 vdd.t2699 7.146
R44196 vdd.n7184 vdd.t2780 7.146
R44197 vdd.n7184 vdd.t116 7.146
R44198 vdd.n7183 vdd.t25 7.146
R44199 vdd.n7183 vdd.t355 7.146
R44200 vdd.n7182 vdd.t1147 7.146
R44201 vdd.n7182 vdd.t1470 7.146
R44202 vdd.n7181 vdd.t700 7.146
R44203 vdd.n7181 vdd.t991 7.146
R44204 vdd.n7180 vdd.t1809 7.146
R44205 vdd.n7180 vdd.t2136 7.146
R44206 vdd.n7179 vdd.t2242 7.146
R44207 vdd.n7179 vdd.t2565 7.146
R44208 vdd.n7178 vdd.t2334 7.146
R44209 vdd.n7178 vdd.t1591 7.146
R44210 vdd.n7177 vdd.t1127 7.146
R44211 vdd.n7177 vdd.t1447 7.146
R44212 vdd.n7176 vdd.t1154 7.146
R44213 vdd.n7176 vdd.t309 7.146
R44214 vdd.n7175 vdd.t33 7.146
R44215 vdd.n7175 vdd.t2159 7.146
R44216 vdd.n7174 vdd.t1892 7.146
R44217 vdd.n7174 vdd.t1013 7.146
R44218 vdd.n7173 vdd.t2363 7.146
R44219 vdd.n7173 vdd.t1496 7.146
R44220 vdd.n7172 vdd.t1230 7.146
R44221 vdd.n7172 vdd.t385 7.146
R44222 vdd.n7171 vdd.t978 7.146
R44223 vdd.n7171 vdd.t143 7.146
R44224 vdd.n7170 vdd.t594 7.146
R44225 vdd.n7170 vdd.t2723 7.146
R44226 vdd.n7379 vdd.t1151 7.146
R44227 vdd.n7379 vdd.t1299 7.146
R44228 vdd.n7368 vdd.t1401 7.146
R44229 vdd.n7368 vdd.t1553 7.146
R44230 vdd.n7367 vdd.t2297 7.146
R44231 vdd.n7367 vdd.t1862 7.146
R44232 vdd.n7366 vdd.t2541 7.146
R44233 vdd.n7366 vdd.t2111 7.146
R44234 vdd.n7365 vdd.t696 7.146
R44235 vdd.n7365 vdd.t267 7.146
R44236 vdd.n7364 vdd.t1099 7.146
R44237 vdd.n7364 vdd.t672 7.146
R44238 vdd.n7363 vdd.t1331 7.146
R44239 vdd.n7363 vdd.t900 7.146
R44240 vdd.n7362 vdd.t2471 7.146
R44241 vdd.n7362 vdd.t2054 7.146
R44242 vdd.n7361 vdd.t1999 7.146
R44243 vdd.n7361 vdd.t1568 7.146
R44244 vdd.n7360 vdd.t156 7.146
R44245 vdd.n7360 vdd.t2718 7.146
R44246 vdd.n7359 vdd.t572 7.146
R44247 vdd.n7359 vdd.t136 7.146
R44248 vdd.n7358 vdd.t933 7.146
R44249 vdd.n7358 vdd.t956 7.146
R44250 vdd.n7357 vdd.t2442 7.146
R44251 vdd.n7357 vdd.t2026 7.146
R44252 vdd.n7356 vdd.t2974 7.146
R44253 vdd.n7356 vdd.t144 7.146
R44254 vdd.n7355 vdd.t1829 7.146
R44255 vdd.n7355 vdd.t1983 7.146
R44256 vdd.n7354 vdd.t724 7.146
R44257 vdd.n7354 vdd.t850 7.146
R44258 vdd.n7353 vdd.t1177 7.146
R44259 vdd.n7353 vdd.t1323 7.146
R44260 vdd.n7352 vdd.t51 7.146
R44261 vdd.n7352 vdd.t209 7.146
R44262 vdd.n7351 vdd.t2798 7.146
R44263 vdd.n7351 vdd.t2954 7.146
R44264 vdd.n7350 vdd.t2379 7.146
R44265 vdd.n7350 vdd.t2533 7.146
R44266 vdd.n7559 vdd.t977 7.146
R44267 vdd.n7559 vdd.t141 7.146
R44268 vdd.n7548 vdd.t1233 7.146
R44269 vdd.n7548 vdd.t384 7.146
R44270 vdd.n7547 vdd.t2866 7.146
R44271 vdd.n7547 vdd.t202 7.146
R44272 vdd.n7546 vdd.t122 7.146
R44273 vdd.n7546 vdd.t446 7.146
R44274 vdd.n7545 vdd.t1242 7.146
R44275 vdd.n7545 vdd.t1565 7.146
R44276 vdd.n7544 vdd.t1649 7.146
R44277 vdd.n7544 vdd.t1975 7.146
R44278 vdd.n7543 vdd.t1904 7.146
R44279 vdd.n7543 vdd.t2233 7.146
R44280 vdd.n7542 vdd.t42 7.146
R44281 vdd.n7542 vdd.t377 7.146
R44282 vdd.n7541 vdd.t2571 7.146
R44283 vdd.n7541 vdd.t2893 7.146
R44284 vdd.n7540 vdd.t719 7.146
R44285 vdd.n7540 vdd.t1007 7.146
R44286 vdd.n7539 vdd.t1112 7.146
R44287 vdd.n7539 vdd.t1426 7.146
R44288 vdd.n7538 vdd.t332 7.146
R44289 vdd.n7538 vdd.t2581 7.146
R44290 vdd.n7537 vdd.t15 7.146
R44291 vdd.n7537 vdd.t346 7.146
R44292 vdd.n7536 vdd.t2804 7.146
R44293 vdd.n7536 vdd.t1935 7.146
R44294 vdd.n7535 vdd.t1665 7.146
R44295 vdd.n7535 vdd.t811 7.146
R44296 vdd.n7534 vdd.t549 7.146
R44297 vdd.n7534 vdd.t2673 7.146
R44298 vdd.n7533 vdd.t999 7.146
R44299 vdd.n7533 vdd.t163 7.146
R44300 vdd.n7532 vdd.t2885 7.146
R44301 vdd.n7532 vdd.t2009 7.146
R44302 vdd.n7531 vdd.t2635 7.146
R44303 vdd.n7531 vdd.t1765 7.146
R44304 vdd.n7530 vdd.t2225 7.146
R44305 vdd.n7530 vdd.t1339 7.146
R44306 vdd.n7739 vdd.t2799 7.146
R44307 vdd.n7739 vdd.t1174 7.146
R44308 vdd.n7728 vdd.t54 7.146
R44309 vdd.n7728 vdd.t1418 7.146
R44310 vdd.n7727 vdd.t1172 7.146
R44311 vdd.n7727 vdd.t2279 7.146
R44312 vdd.n7726 vdd.t1415 7.146
R44313 vdd.n7726 vdd.t2513 7.146
R44314 vdd.n7725 vdd.t2567 7.146
R44315 vdd.n7725 vdd.t664 7.146
R44316 vdd.n7724 vdd.t2971 7.146
R44317 vdd.n7724 vdd.t1077 7.146
R44318 vdd.n7723 vdd.t240 7.146
R44319 vdd.n7723 vdd.t1307 7.146
R44320 vdd.n7722 vdd.t1352 7.146
R44321 vdd.n7722 vdd.t2448 7.146
R44322 vdd.n7721 vdd.t873 7.146
R44323 vdd.n7721 vdd.t1971 7.146
R44324 vdd.n7720 vdd.t2017 7.146
R44325 vdd.n7720 vdd.t128 7.146
R44326 vdd.n7719 vdd.t2421 7.146
R44327 vdd.n7719 vdd.t539 7.146
R44328 vdd.n7718 vdd.t1922 7.146
R44329 vdd.n7718 vdd.t1047 7.146
R44330 vdd.n7717 vdd.t1319 7.146
R44331 vdd.n7717 vdd.t2415 7.146
R44332 vdd.n7716 vdd.t1613 7.146
R44333 vdd.n7716 vdd.t2998 7.146
R44334 vdd.n7715 vdd.t489 7.146
R44335 vdd.n7715 vdd.t1854 7.146
R44336 vdd.n7714 vdd.t2337 7.146
R44337 vdd.n7714 vdd.t747 7.146
R44338 vdd.n7713 vdd.t2822 7.146
R44339 vdd.n7713 vdd.t1196 7.146
R44340 vdd.n7712 vdd.t1682 7.146
R44341 vdd.n7712 vdd.t77 7.146
R44342 vdd.n7711 vdd.t1434 7.146
R44343 vdd.n7711 vdd.t2820 7.146
R44344 vdd.n7710 vdd.t1017 7.146
R44345 vdd.n7710 vdd.t2396 7.146
R44346 vdd.n7919 vdd.t343 7.146
R44347 vdd.n7919 vdd.t686 7.146
R44348 vdd.n7908 vdd.t596 7.146
R44349 vdd.n7908 vdd.t907 7.146
R44350 vdd.n7907 vdd.t2828 7.146
R44351 vdd.n7907 vdd.t858 7.146
R44352 vdd.n7906 vdd.t88 7.146
R44353 vdd.n7906 vdd.t1102 7.146
R44354 vdd.n7905 vdd.t1210 7.146
R44355 vdd.n7905 vdd.t2247 7.146
R44356 vdd.n7904 vdd.t1624 7.146
R44357 vdd.n7904 vdd.t2656 7.146
R44358 vdd.n7903 vdd.t1868 7.146
R44359 vdd.n7903 vdd.t2905 7.146
R44360 vdd.n7902 vdd.t11 7.146
R44361 vdd.n7902 vdd.t1024 7.146
R44362 vdd.n7901 vdd.t2527 7.146
R44363 vdd.n7901 vdd.t575 7.146
R44364 vdd.n7900 vdd.t679 7.146
R44365 vdd.n7900 vdd.t1688 7.146
R44366 vdd.n7899 vdd.t1087 7.146
R44367 vdd.n7899 vdd.t2109 7.146
R44368 vdd.n7898 vdd.t2495 7.146
R44369 vdd.n7898 vdd.t2683 7.146
R44370 vdd.n7897 vdd.t2978 7.146
R44371 vdd.n7897 vdd.t997 7.146
R44372 vdd.n7896 vdd.t2149 7.146
R44373 vdd.n7896 vdd.t2479 7.146
R44374 vdd.n7895 vdd.t1003 7.146
R44375 vdd.n7895 vdd.t1348 7.146
R44376 vdd.n7894 vdd.t2886 7.146
R44377 vdd.n7894 vdd.t235 7.146
R44378 vdd.n7893 vdd.t368 7.146
R44379 vdd.n7893 vdd.t712 7.146
R44380 vdd.n7892 vdd.t2228 7.146
R44381 vdd.n7892 vdd.t2562 7.146
R44382 vdd.n7891 vdd.t1967 7.146
R44383 vdd.n7891 vdd.t2307 7.146
R44384 vdd.n7890 vdd.t1557 7.146
R44385 vdd.n7890 vdd.t1897 7.146
R44386 vdd.n8099 vdd.t2399 7.146
R44387 vdd.n8099 vdd.t1197 7.146
R44388 vdd.n8088 vdd.t2654 7.146
R44389 vdd.n8088 vdd.t1436 7.146
R44390 vdd.n8087 vdd.t1165 7.146
R44391 vdd.n8087 vdd.t2502 7.146
R44392 vdd.n8086 vdd.t1409 7.146
R44393 vdd.n8086 vdd.t2764 7.146
R44394 vdd.n8085 vdd.t2555 7.146
R44395 vdd.n8085 vdd.t889 7.146
R44396 vdd.n8084 vdd.t2966 7.146
R44397 vdd.n8084 vdd.t1294 7.146
R44398 vdd.n8083 vdd.t230 7.146
R44399 vdd.n8083 vdd.t1549 7.146
R44400 vdd.n8082 vdd.t1344 7.146
R44401 vdd.n8082 vdd.t2703 7.146
R44402 vdd.n8081 vdd.t870 7.146
R44403 vdd.n8081 vdd.t2220 7.146
R44404 vdd.n8080 vdd.t2010 7.146
R44405 vdd.n8080 vdd.t359 7.146
R44406 vdd.n8079 vdd.t2412 7.146
R44407 vdd.n8079 vdd.t781 7.146
R44408 vdd.n8078 vdd.t1764 7.146
R44409 vdd.n8078 vdd.t276 7.146
R44410 vdd.n8077 vdd.t1316 7.146
R44411 vdd.n8077 vdd.t2664 7.146
R44412 vdd.n8076 vdd.t1220 7.146
R44413 vdd.n8076 vdd.t21 7.146
R44414 vdd.n8075 vdd.t104 7.146
R44415 vdd.n8075 vdd.t1878 7.146
R44416 vdd.n8074 vdd.t1943 7.146
R44417 vdd.n8074 vdd.t766 7.146
R44418 vdd.n8073 vdd.t2422 7.146
R44419 vdd.n8073 vdd.t1217 7.146
R44420 vdd.n8072 vdd.t1279 7.146
R44421 vdd.n8072 vdd.t101 7.146
R44422 vdd.n8071 vdd.t1048 7.146
R44423 vdd.n8071 vdd.t2840 7.146
R44424 vdd.n8070 vdd.t640 7.146
R44425 vdd.n8070 vdd.t2413 7.146
R44426 vdd.n8279 vdd.t1215 7.146
R44427 vdd.n8279 vdd.t16 7.146
R44428 vdd.n8268 vdd.t1454 7.146
R44429 vdd.n8268 vdd.t278 7.146
R44430 vdd.n8267 vdd.t2480 7.146
R44431 vdd.n8267 vdd.t831 7.146
R44432 vdd.n8266 vdd.t2743 7.146
R44433 vdd.n8266 vdd.t1074 7.146
R44434 vdd.n8265 vdd.t866 7.146
R44435 vdd.n8265 vdd.t2218 7.146
R44436 vdd.n8264 vdd.t1274 7.146
R44437 vdd.n8264 vdd.t2627 7.146
R44438 vdd.n8263 vdd.t1521 7.146
R44439 vdd.n8263 vdd.t2873 7.146
R44440 vdd.n8262 vdd.t2669 7.146
R44441 vdd.n8262 vdd.t992 7.146
R44442 vdd.n8261 vdd.t2198 7.146
R44443 vdd.n8261 vdd.t537 7.146
R44444 vdd.n8260 vdd.t336 7.146
R44445 vdd.n8260 vdd.t1654 7.146
R44446 vdd.n8259 vdd.t761 7.146
R44447 vdd.n8259 vdd.t2088 7.146
R44448 vdd.n8258 vdd.t378 7.146
R44449 vdd.n8258 vdd.t1844 7.146
R44450 vdd.n8257 vdd.t2642 7.146
R44451 vdd.n8257 vdd.t961 7.146
R44452 vdd.n8256 vdd.t43 7.146
R44453 vdd.n8256 vdd.t1821 7.146
R44454 vdd.n8255 vdd.t1905 7.146
R44455 vdd.n8255 vdd.t713 7.146
R44456 vdd.n8254 vdd.t784 7.146
R44457 vdd.n8254 vdd.t2563 7.146
R44458 vdd.n8253 vdd.t1241 7.146
R44459 vdd.n8253 vdd.t38 7.146
R44460 vdd.n8252 vdd.t121 7.146
R44461 vdd.n8252 vdd.t1898 7.146
R44462 vdd.n8251 vdd.t2867 7.146
R44463 vdd.n8251 vdd.t1644 7.146
R44464 vdd.n8250 vdd.t2437 7.146
R44465 vdd.n8250 vdd.t1235 7.146
R44466 vdd.n8459 vdd.t2711 7.146
R44467 vdd.n8459 vdd.t2841 7.146
R44468 vdd.n8448 vdd.t2937 7.146
R44469 vdd.n8448 vdd.t102 7.146
R44470 vdd.n8447 vdd.t1815 7.146
R44471 vdd.n8447 vdd.t1390 7.146
R44472 vdd.n8446 vdd.t2075 7.146
R44473 vdd.n8446 vdd.t1631 7.146
R44474 vdd.n8445 vdd.t219 7.146
R44475 vdd.n8445 vdd.t2775 7.146
R44476 vdd.n8444 vdd.t627 7.146
R44477 vdd.n8444 vdd.t206 7.146
R44478 vdd.n8443 vdd.t859 7.146
R44479 vdd.n8443 vdd.t448 7.146
R44480 vdd.n8442 vdd.t2000 7.146
R44481 vdd.n8442 vdd.t1569 7.146
R44482 vdd.n8441 vdd.t1512 7.146
R44483 vdd.n8441 vdd.t1093 7.146
R44484 vdd.n8440 vdd.t2658 7.146
R44485 vdd.n8440 vdd.t2236 7.146
R44486 vdd.n8439 vdd.t85 7.146
R44487 vdd.n8439 vdd.t2644 7.146
R44488 vdd.n8438 vdd.t1203 7.146
R44489 vdd.n8438 vdd.t1227 7.146
R44490 vdd.n8437 vdd.t1968 7.146
R44491 vdd.n8437 vdd.t1538 7.146
R44492 vdd.n8436 vdd.t1504 7.146
R44493 vdd.n8436 vdd.t1651 7.146
R44494 vdd.n8435 vdd.t396 7.146
R44495 vdd.n8435 vdd.t532 7.146
R44496 vdd.n8434 vdd.t2250 7.146
R44497 vdd.n8434 vdd.t2380 7.146
R44498 vdd.n8433 vdd.t2729 7.146
R44499 vdd.n8433 vdd.t2871 7.146
R44500 vdd.n8432 vdd.t1578 7.146
R44501 vdd.n8432 vdd.t1728 7.146
R44502 vdd.n8431 vdd.t1327 7.146
R44503 vdd.n8431 vdd.t1476 7.146
R44504 vdd.n8430 vdd.t910 7.146
R44505 vdd.n8430 vdd.t1068 7.146
R44506 vdd.n8639 vdd.t2519 7.146
R44507 vdd.n8639 vdd.t897 7.146
R44508 vdd.n8628 vdd.t2773 7.146
R44509 vdd.n8628 vdd.t1135 7.146
R44510 vdd.n8627 vdd.t2377 7.146
R44511 vdd.n8627 vdd.t490 7.146
R44512 vdd.n8626 vdd.t2630 7.146
R44513 vdd.n8626 vdd.t749 7.146
R44514 vdd.n8625 vdd.t785 7.146
R44515 vdd.n8625 vdd.t1856 7.146
R44516 vdd.n8624 vdd.t1175 7.146
R44517 vdd.n8624 vdd.t2281 7.146
R44518 vdd.n8623 vdd.t1416 7.146
R44519 vdd.n8623 vdd.t2518 7.146
R44520 vdd.n8622 vdd.t2572 7.146
R44521 vdd.n8622 vdd.t669 7.146
R44522 vdd.n8621 vdd.t2093 7.146
R44523 vdd.n8621 vdd.t203 7.146
R44524 vdd.n8620 vdd.t242 7.146
R44525 vdd.n8620 vdd.t1310 7.146
R44526 vdd.n8619 vdd.t644 7.146
R44527 vdd.n8619 vdd.t1736 7.146
R44528 vdd.n8618 vdd.t601 7.146
R44529 vdd.n8618 vdd.t2725 7.146
R44530 vdd.n8617 vdd.t2535 7.146
R44531 vdd.n8617 vdd.t642 7.146
R44532 vdd.n8616 vdd.t1335 7.146
R44533 vdd.n8616 vdd.t2735 7.146
R44534 vdd.n8615 vdd.t223 7.146
R44535 vdd.n8615 vdd.t1581 7.146
R44536 vdd.n8614 vdd.t2078 7.146
R44537 vdd.n8614 vdd.t460 7.146
R44538 vdd.n8613 vdd.t2546 7.146
R44539 vdd.n8613 vdd.t916 7.146
R44540 vdd.n8612 vdd.t1402 7.146
R44541 vdd.n8612 vdd.t2784 7.146
R44542 vdd.n8611 vdd.t1153 7.146
R44543 vdd.n8611 vdd.t2542 7.146
R44544 vdd.n8610 vdd.t769 7.146
R44545 vdd.n8610 vdd.t2121 7.146
R44546 vdd.n8819 vdd.t1329 7.146
R44547 vdd.n8819 vdd.t2730 7.146
R44548 vdd.n8808 vdd.t1579 7.146
R44549 vdd.n8808 vdd.t2959 7.146
R44550 vdd.n8807 vdd.t723 7.146
R44551 vdd.n8807 vdd.t1793 7.146
R44552 vdd.n8806 vdd.t934 7.146
R44553 vdd.n8806 vdd.t2055 7.146
R44554 vdd.n8805 vdd.t2089 7.146
R44555 vdd.n8805 vdd.t199 7.146
R44556 vdd.n8804 vdd.t2492 7.146
R44557 vdd.n8804 vdd.t611 7.146
R44558 vdd.n8803 vdd.t2751 7.146
R44559 vdd.n8803 vdd.t838 7.146
R44560 vdd.n8802 vdd.t877 7.146
R44561 vdd.n8802 vdd.t1972 7.146
R44562 vdd.n8801 vdd.t420 7.146
R44563 vdd.n8801 vdd.t1493 7.146
R44564 vdd.n8800 vdd.t1531 7.146
R44565 vdd.n8800 vdd.t2638 7.146
R44566 vdd.n8799 vdd.t1947 7.146
R44567 vdd.n8799 vdd.t59 7.146
R44568 vdd.n8798 vdd.t2185 7.146
R44569 vdd.n8798 vdd.t1297 7.146
R44570 vdd.n8797 vdd.t851 7.146
R44571 vdd.n8797 vdd.t1944 7.146
R44572 vdd.n8796 vdd.t171 7.146
R44573 vdd.n8796 vdd.t1525 7.146
R44574 vdd.n8795 vdd.t2023 7.146
R44575 vdd.n8795 vdd.t414 7.146
R44576 vdd.n8794 vdd.t879 7.146
R44577 vdd.n8794 vdd.t2265 7.146
R44578 vdd.n8793 vdd.t1358 7.146
R44579 vdd.n8793 vdd.t2748 7.146
R44580 vdd.n8792 vdd.t241 7.146
R44581 vdd.n8792 vdd.t1595 7.146
R44582 vdd.n8791 vdd.t2973 7.146
R44583 vdd.n8791 vdd.t1356 7.146
R44584 vdd.n8790 vdd.t2573 7.146
R44585 vdd.n8790 vdd.t930 7.146
R44586 vdd.n8999 vdd.t2386 7.146
R44587 vdd.n8999 vdd.t2544 7.146
R44588 vdd.n8988 vdd.t2640 7.146
R44589 vdd.n8988 vdd.t2785 7.146
R44590 vdd.n8987 vdd.t2791 7.146
R44591 vdd.n8987 vdd.t2356 7.146
R44592 vdd.n8986 vdd.t44 7.146
R44593 vdd.n8986 vdd.t2613 7.146
R44594 vdd.n8985 vdd.t1166 7.146
R44595 vdd.n8985 vdd.t763 7.146
R44596 vdd.n8984 vdd.t1590 7.146
R44597 vdd.n8984 vdd.t1146 7.146
R44598 vdd.n8983 vdd.t1823 7.146
R44599 vdd.n8983 vdd.t1398 7.146
R44600 vdd.n8982 vdd.t2967 7.146
R44601 vdd.n8982 vdd.t2537 7.146
R44602 vdd.n8981 vdd.t2487 7.146
R44603 vdd.n8981 vdd.t2072 7.146
R44604 vdd.n8980 vdd.t635 7.146
R44605 vdd.n8980 vdd.t216 7.146
R44606 vdd.n8979 vdd.t1041 7.146
R44607 vdd.n8979 vdd.t624 7.146
R44608 vdd.n8978 vdd.t670 7.146
R44609 vdd.n8978 vdd.t707 7.146
R44610 vdd.n8977 vdd.t2946 7.146
R44611 vdd.n8977 vdd.t2505 7.146
R44612 vdd.n8976 vdd.t1211 7.146
R44613 vdd.n8976 vdd.t1360 7.146
R44614 vdd.n8975 vdd.t89 7.146
R44615 vdd.n8975 vdd.t243 7.146
R44616 vdd.n8974 vdd.t1932 7.146
R44617 vdd.n8974 vdd.t2094 7.146
R44618 vdd.n8973 vdd.t2406 7.146
R44619 vdd.n8973 vdd.t2577 7.146
R44620 vdd.n8972 vdd.t1268 7.146
R44621 vdd.n8972 vdd.t1421 7.146
R44622 vdd.n8971 vdd.t1028 7.146
R44623 vdd.n8971 vdd.t1178 7.146
R44624 vdd.n8970 vdd.t628 7.146
R44625 vdd.n8970 vdd.t790 7.146
R44626 vdd.n9179 vdd.t2235 7.146
R44627 vdd.n9179 vdd.t1005 7.146
R44628 vdd.n9168 vdd.t2462 7.146
R44629 vdd.n9168 vdd.t1257 7.146
R44630 vdd.n9167 vdd.t375 7.146
R44631 vdd.n9167 vdd.t1695 7.146
R44632 vdd.n9166 vdd.t616 7.146
R44633 vdd.n9166 vdd.t1936 7.146
R44634 vdd.n9165 vdd.t1738 7.146
R44635 vdd.n9165 vdd.t91 7.146
R44636 vdd.n9164 vdd.t2153 7.146
R44637 vdd.n9164 vdd.t499 7.146
R44638 vdd.n9163 vdd.t2390 7.146
R44639 vdd.n9163 vdd.t756 7.146
R44640 vdd.n9162 vdd.t543 7.146
R44641 vdd.n9162 vdd.t1869 7.146
R44642 vdd.n9161 vdd.t69 7.146
R44643 vdd.n9161 vdd.t1393 7.146
R44644 vdd.n9160 vdd.t1186 7.146
R44645 vdd.n9160 vdd.t2528 7.146
R44646 vdd.n9159 vdd.t1602 7.146
R44647 vdd.n9159 vdd.t2949 7.146
R44648 vdd.n9158 vdd.t45 7.146
R44649 vdd.n9158 vdd.t1527 7.146
R44650 vdd.n9157 vdd.t521 7.146
R44651 vdd.n9157 vdd.t1834 7.146
R44652 vdd.n9156 vdd.t1038 7.146
R44653 vdd.n9156 vdd.t2833 7.146
R44654 vdd.n9155 vdd.t2914 7.146
R44655 vdd.n9155 vdd.t1697 7.146
R44656 vdd.n9154 vdd.t1768 7.146
R44657 vdd.n9154 vdd.t579 7.146
R44658 vdd.n9153 vdd.t2255 7.146
R44659 vdd.n9153 vdd.t1031 7.146
R44660 vdd.n9152 vdd.t1107 7.146
R44661 vdd.n9152 vdd.t2910 7.146
R44662 vdd.n9151 vdd.t860 7.146
R44663 vdd.n9151 vdd.t2659 7.146
R44664 vdd.n9150 vdd.t463 7.146
R44665 vdd.n9150 vdd.t2252 7.146
R44666 vdd.n9359 vdd.t1032 7.146
R44667 vdd.n9359 vdd.t2825 7.146
R44668 vdd.n9348 vdd.t1270 7.146
R44669 vdd.n9348 vdd.t86 7.146
R44670 vdd.n9347 vdd.t1669 7.146
R44671 vdd.n9347 vdd.t14 7.146
R44672 vdd.n9346 vdd.t1920 7.146
R44673 vdd.n9346 vdd.t277 7.146
R44674 vdd.n9345 vdd.t63 7.146
R44675 vdd.n9345 vdd.t1392 7.146
R44676 vdd.n9344 vdd.t475 7.146
R44677 vdd.n9344 vdd.t1799 7.146
R44678 vdd.n9343 vdd.t733 7.146
R44679 vdd.n9343 vdd.t2063 7.146
R44680 vdd.n9342 vdd.t1837 7.146
R44681 vdd.n9342 vdd.t207 7.146
R44682 vdd.n9341 vdd.t1375 7.146
R44683 vdd.n9341 vdd.t2726 7.146
R44684 vdd.n9340 vdd.t2500 7.146
R44685 vdd.n9340 vdd.t846 7.146
R44686 vdd.n9339 vdd.t2927 7.146
R44687 vdd.n9339 vdd.t1261 7.146
R44688 vdd.n9338 vdd.t1633 7.146
R44689 vdd.n9338 vdd.t151 7.146
R44690 vdd.n9337 vdd.t1818 7.146
R44691 vdd.n9337 vdd.t178 7.146
R44692 vdd.n9336 vdd.t2857 7.146
R44693 vdd.n9336 vdd.t1639 7.146
R44694 vdd.n9335 vdd.t1717 7.146
R44695 vdd.n9335 vdd.t523 7.146
R44696 vdd.n9334 vdd.t600 7.146
R44697 vdd.n9334 vdd.t2366 7.146
R44698 vdd.n9333 vdd.t1059 7.146
R44699 vdd.n9333 vdd.t2848 7.146
R44700 vdd.n9332 vdd.t2924 7.146
R44701 vdd.n9332 vdd.t1711 7.146
R44702 vdd.n9331 vdd.t2688 7.146
R44703 vdd.n9331 vdd.t1457 7.146
R44704 vdd.n9330 vdd.t2267 7.146
R44705 vdd.n9330 vdd.t1055 7.146
R44706 vdd.n9539 vdd.t2849 7.146
R44707 vdd.n9539 vdd.t1910 7.146
R44708 vdd.n9528 vdd.t109 7.146
R44709 vdd.n9528 vdd.t2150 7.146
R44710 vdd.n9527 vdd.t2989 7.146
R44711 vdd.n9527 vdd.t1349 7.146
R44712 vdd.n9526 vdd.t255 7.146
R44713 vdd.n9526 vdd.t1594 7.146
R44714 vdd.n9525 vdd.t1372 7.146
R44715 vdd.n9525 vdd.t2744 7.146
R44716 vdd.n9524 vdd.t1783 7.146
R44717 vdd.n9524 vdd.t168 7.146
R44718 vdd.n9523 vdd.t2040 7.146
R44719 vdd.n9523 vdd.t413 7.146
R44720 vdd.n9522 vdd.t185 7.146
R44721 vdd.n9522 vdd.t1524 7.146
R44722 vdd.n9521 vdd.t2707 7.146
R44723 vdd.n9521 vdd.t1053 7.146
R44724 vdd.n9520 vdd.t832 7.146
R44725 vdd.n9520 vdd.t2199 7.146
R44726 vdd.n9519 vdd.t1243 7.146
R44727 vdd.n9519 vdd.t2612 7.146
R44728 vdd.n9518 vdd.t257 7.146
R44729 vdd.n9518 vdd.t2383 7.146
R44730 vdd.n9517 vdd.t161 7.146
R44731 vdd.n9517 vdd.t1500 7.146
R44732 vdd.n9516 vdd.t1657 7.146
R44733 vdd.n9516 vdd.t744 7.146
R44734 vdd.n9515 vdd.t540 7.146
R44735 vdd.n9515 vdd.t2596 7.146
R44736 vdd.n9514 vdd.t2385 7.146
R44737 vdd.n9514 vdd.t1441 7.146
R44738 vdd.n9513 vdd.t2875 7.146
R44739 vdd.n9513 vdd.t1925 7.146
R44740 vdd.n9512 vdd.t1734 7.146
R44741 vdd.n9512 vdd.t805 7.146
R44742 vdd.n9511 vdd.t1480 7.146
R44743 vdd.n9511 vdd.t564 7.146
R44744 vdd.n9510 vdd.t1078 7.146
R44745 vdd.n9510 vdd.t149 7.146
R44746 vdd.n9719 vdd.t1653 7.146
R44747 vdd.n9719 vdd.t737 7.146
R44748 vdd.n9708 vdd.t1909 7.146
R44749 vdd.n9708 vdd.t951 7.146
R44750 vdd.n9707 vdd.t1290 7.146
R44751 vdd.n9707 vdd.t2677 7.146
R44752 vdd.n9706 vdd.t1550 7.146
R44753 vdd.n9706 vdd.t2919 7.146
R44754 vdd.n9705 vdd.t2702 7.146
R44755 vdd.n9705 vdd.t1049 7.146
R44756 vdd.n9704 vdd.t119 7.146
R44757 vdd.n9704 vdd.t1455 7.146
R44758 vdd.n9703 vdd.t358 7.146
R44759 vdd.n9703 vdd.t1707 7.146
R44760 vdd.n9702 vdd.t1477 7.146
R44761 vdd.n9702 vdd.t2845 7.146
R44762 vdd.n9701 vdd.t995 7.146
R44763 vdd.n9701 vdd.t2361 7.146
R44764 vdd.n9700 vdd.t2141 7.146
R44765 vdd.n9700 vdd.t516 7.146
R44766 vdd.n9699 vdd.t2568 7.146
R44767 vdd.n9699 vdd.t911 7.146
R44768 vdd.n9698 vdd.t1824 7.146
R44769 vdd.n9698 vdd.t974 7.146
R44770 vdd.n9697 vdd.t1451 7.146
R44771 vdd.n9697 vdd.t2818 7.146
R44772 vdd.n9696 vdd.t482 7.146
R44773 vdd.n9696 vdd.t2534 7.146
R44774 vdd.n9695 vdd.t2330 7.146
R44775 vdd.n9695 vdd.t1397 7.146
R44776 vdd.n9694 vdd.t1201 7.146
R44777 vdd.n9694 vdd.t282 7.146
R44778 vdd.n9693 vdd.t1676 7.146
R44779 vdd.n9693 vdd.t759 7.146
R44780 vdd.n9692 vdd.t561 7.146
R44781 vdd.n9692 vdd.t2609 7.146
R44782 vdd.n9691 vdd.t314 7.146
R44783 vdd.n9691 vdd.t2347 7.146
R44784 vdd.n9690 vdd.t2897 7.146
R44785 vdd.n9690 vdd.t1937 7.146
R44786 vdd.n9899 vdd.t418 7.146
R44787 vdd.n9899 vdd.t2525 7.146
R44788 vdd.n9888 vdd.t647 7.146
R44789 vdd.n9888 vdd.t2779 7.146
R44790 vdd.n9887 vdd.t673 7.146
R44791 vdd.n9887 vdd.t970 7.146
R44792 vdd.n9886 vdd.t901 7.146
R44793 vdd.n9886 vdd.t1224 7.146
R44794 vdd.n9885 vdd.t2056 7.146
R44795 vdd.n9885 vdd.t2359 7.146
R44796 vdd.n9884 vdd.t2452 7.146
R44797 vdd.n9884 vdd.t2781 7.146
R44798 vdd.n9883 vdd.t2719 7.146
R44799 vdd.n9883 vdd.t29 7.146
R44800 vdd.n9882 vdd.t839 7.146
R44801 vdd.n9882 vdd.t1150 7.146
R44802 vdd.n9881 vdd.t382 7.146
R44803 vdd.n9881 vdd.t703 7.146
R44804 vdd.n9880 vdd.t1494 7.146
R44805 vdd.n9880 vdd.t1813 7.146
R44806 vdd.n9879 vdd.t1918 7.146
R44807 vdd.n9879 vdd.t2248 7.146
R44808 vdd.n9878 vdd.t351 7.146
R44809 vdd.n9878 vdd.t2598 7.146
R44810 vdd.n9877 vdd.t823 7.146
R44811 vdd.n9877 vdd.t1128 7.146
R44812 vdd.n9876 vdd.t2226 7.146
R44813 vdd.n9876 vdd.t1340 7.146
R44814 vdd.n9875 vdd.t1081 7.146
R44815 vdd.n9875 vdd.t228 7.146
R44816 vdd.n9874 vdd.t2944 7.146
R44817 vdd.n9874 vdd.t2081 7.146
R44818 vdd.n9873 vdd.t436 7.146
R44819 vdd.n9873 vdd.t2552 7.146
R44820 vdd.n9872 vdd.t2282 7.146
R44821 vdd.n9872 vdd.t1406 7.146
R44822 vdd.n9871 vdd.t2048 7.146
R44823 vdd.n9871 vdd.t1159 7.146
R44824 vdd.n9870 vdd.t1615 7.146
R44825 vdd.n9870 vdd.t772 7.146
R44826 vdd.n10079 vdd.t920 7.146
R44827 vdd.n10079 vdd.t70 7.146
R44828 vdd.n10068 vdd.t1161 7.146
R44829 vdd.n10068 vdd.t315 7.146
R44830 vdd.n10067 vdd.t2313 7.146
R44831 vdd.n10067 vdd.t2643 7.146
R44832 vdd.n10066 vdd.t2575 7.146
R44833 vdd.n10066 vdd.t2895 7.146
R44834 vdd.n10065 vdd.t720 7.146
R44835 vdd.n10065 vdd.t1010 7.146
R44836 vdd.n10064 vdd.t1114 7.146
R44837 vdd.n10064 vdd.t1427 7.146
R44838 vdd.n10063 vdd.t1359 7.146
R44839 vdd.n10063 vdd.t1672 7.146
R44840 vdd.n10062 vdd.t2489 7.146
R44841 vdd.n10062 vdd.t2812 7.146
R44842 vdd.n10061 vdd.t2025 7.146
R44843 vdd.n10061 vdd.t2324 7.146
R44844 vdd.n10060 vdd.t172 7.146
R44845 vdd.n10060 vdd.t477 7.146
R44846 vdd.n10059 vdd.t591 7.146
R44847 vdd.n10059 vdd.t890 7.146
R44848 vdd.n10058 vdd.t917 7.146
R44849 vdd.n10058 vdd.t187 7.146
R44850 vdd.n10057 vdd.t2464 7.146
R44851 vdd.n10057 vdd.t2787 7.146
R44852 vdd.n10056 vdd.t2753 7.146
R44853 vdd.n10056 vdd.t1873 7.146
R44854 vdd.n10055 vdd.t1599 7.146
R44855 vdd.n10055 vdd.t760 7.146
R44856 vdd.n10054 vdd.t476 7.146
R44857 vdd.n10054 vdd.t2610 7.146
R44858 vdd.n10053 vdd.t935 7.146
R44859 vdd.n10053 vdd.t98 7.146
R44860 vdd.n10052 vdd.t2806 7.146
R44861 vdd.n10052 vdd.t1938 7.146
R44862 vdd.n10051 vdd.t2579 7.146
R44863 vdd.n10051 vdd.t1699 7.146
R44864 vdd.n10050 vdd.t2151 7.146
R44865 vdd.n10050 vdd.t1272 7.146
R44866 vdd.n10259 vdd.t2750 7.146
R44867 vdd.n10259 vdd.t2900 7.146
R44868 vdd.n10248 vdd.t2979 7.146
R44869 vdd.n10248 vdd.t152 7.146
R44870 vdd.n10247 vdd.t643 7.146
R44871 vdd.n10247 vdd.t220 7.146
R44872 vdd.n10246 vdd.t878 7.146
R44873 vdd.n10246 vdd.t461 7.146
R44874 vdd.n10245 vdd.t2020 7.146
R44875 vdd.n10245 vdd.t1582 7.146
R44876 vdd.n10244 vdd.t2424 7.146
R44877 vdd.n10244 vdd.t2001 7.146
R44878 vdd.n10243 vdd.t2684 7.146
R44879 vdd.n10243 vdd.t2253 7.146
R44880 vdd.n10242 vdd.t818 7.146
R44881 vdd.n10242 vdd.t400 7.146
R44882 vdd.n10241 vdd.t344 7.146
R44883 vdd.n10241 vdd.t2911 7.146
R44884 vdd.n10240 vdd.t1458 7.146
R44885 vdd.n10240 vdd.t1034 7.146
R44886 vdd.n10239 vdd.t1883 7.146
R44887 vdd.n10239 vdd.t1446 7.146
R44888 vdd.n10238 vdd.t2515 7.146
R44889 vdd.n10238 vdd.t2548 7.146
R44890 vdd.n10237 vdd.t800 7.146
R44891 vdd.n10237 vdd.t369 7.146
R44892 vdd.n10236 vdd.t1558 7.146
R44893 vdd.n10236 vdd.t1704 7.146
R44894 vdd.n10235 vdd.t438 7.146
R44895 vdd.n10235 vdd.t588 7.146
R44896 vdd.n10234 vdd.t2284 7.146
R44897 vdd.n10234 vdd.t2425 7.146
R44898 vdd.n10233 vdd.t2769 7.146
R44899 vdd.n10233 vdd.t2917 7.146
R44900 vdd.n10232 vdd.t1620 7.146
R44901 vdd.n10232 vdd.t1772 7.146
R44902 vdd.n10231 vdd.t1381 7.146
R44903 vdd.n10231 vdd.t1522 7.146
R44904 vdd.n10230 vdd.t952 7.146
R44905 vdd.n10230 vdd.t1109 7.146
R44906 vdd.n10439 vdd.t2582 7.146
R44907 vdd.n10439 vdd.t936 7.146
R44908 vdd.n10428 vdd.t2808 7.146
R44909 vdd.n10428 vdd.t1183 7.146
R44910 vdd.n10427 vdd.t1193 7.146
R44911 vdd.n10427 vdd.t2292 7.146
R44912 vdd.n10426 vdd.t1430 7.146
R44913 vdd.n10426 vdd.t2540 7.146
R44914 vdd.n10425 vdd.t2588 7.146
R44915 vdd.n10425 vdd.t690 7.146
R44916 vdd.n10424 vdd.t2993 7.146
R44917 vdd.n10424 vdd.t1098 7.146
R44918 vdd.n10423 vdd.t260 7.146
R44919 vdd.n10423 vdd.t1330 7.146
R44920 vdd.n10422 vdd.t1376 7.146
R44921 vdd.n10422 vdd.t2469 7.146
R44922 vdd.n10421 vdd.t895 7.146
R44923 vdd.n10421 vdd.t1996 7.146
R44924 vdd.n10420 vdd.t2043 7.146
R44925 vdd.n10420 vdd.t153 7.146
R44926 vdd.n10419 vdd.t2443 7.146
R44927 vdd.n10419 vdd.t566 7.146
R44928 vdd.n10418 vdd.t1901 7.146
R44929 vdd.n10418 vdd.t1018 7.146
R44930 vdd.n10417 vdd.t1343 7.146
R44931 vdd.n10417 vdd.t2440 7.146
R44932 vdd.n10416 vdd.t1387 7.146
R44933 vdd.n10416 vdd.t2772 7.146
R44934 vdd.n10415 vdd.t272 7.146
R44935 vdd.n10415 vdd.t1625 7.146
R44936 vdd.n10414 vdd.t2113 7.146
R44937 vdd.n10414 vdd.t497 7.146
R44938 vdd.n10413 vdd.t2601 7.146
R44939 vdd.n10413 vdd.t955 7.146
R44940 vdd.n10412 vdd.t1444 7.146
R44941 vdd.n10412 vdd.t2829 7.146
R44942 vdd.n10411 vdd.t1208 7.146
R44943 vdd.n10411 vdd.t2599 7.146
R44944 vdd.n10410 vdd.t808 7.146
R44945 vdd.n10410 vdd.t2177 7.146
R44946 vdd.n10619 vdd.t1383 7.146
R44947 vdd.n10619 vdd.t2410 7.146
R44948 vdd.n10608 vdd.t1621 7.146
R44949 vdd.n10608 vdd.t2670 7.146
R44950 vdd.n10607 vdd.t2506 7.146
R44951 vdd.n10607 vdd.t1627 7.146
R44952 vdd.n10606 vdd.t2767 7.146
R44953 vdd.n10606 vdd.t1870 7.146
R44954 vdd.n10605 vdd.t893 7.146
R44955 vdd.n10605 vdd.t12 7.146
R44956 vdd.n10604 vdd.t1298 7.146
R44957 vdd.n10604 vdd.t445 7.146
R44958 vdd.n10603 vdd.t1552 7.146
R44959 vdd.n10603 vdd.t680 7.146
R44960 vdd.n10602 vdd.t2708 7.146
R44961 vdd.n10602 vdd.t1797 7.146
R44962 vdd.n10601 vdd.t2221 7.146
R44963 vdd.n10601 vdd.t1320 7.146
R44964 vdd.n10600 vdd.t361 7.146
R44965 vdd.n10600 vdd.t2458 7.146
R44966 vdd.n10599 vdd.t786 7.146
R44967 vdd.n10599 vdd.t2894 7.146
R44968 vdd.n10598 vdd.t506 7.146
R44969 vdd.n10598 vdd.t1871 7.146
R44970 vdd.n10597 vdd.t2671 7.146
R44971 vdd.n10597 vdd.t1776 7.146
R44972 vdd.n10596 vdd.t214 7.146
R44973 vdd.n10596 vdd.t1236 7.146
R44974 vdd.n10595 vdd.t2071 7.146
R44975 vdd.n10595 vdd.t117 7.146
R44976 vdd.n10594 vdd.t918 7.146
R44977 vdd.n10594 vdd.t1954 7.146
R44978 vdd.n10593 vdd.t1399 7.146
R44979 vdd.n10593 vdd.t2434 7.146
R44980 vdd.n10592 vdd.t286 7.146
R44981 vdd.n10592 vdd.t1291 7.146
R44982 vdd.n10591 vdd.t24 7.146
R44983 vdd.n10591 vdd.t1061 7.146
R44984 vdd.n10590 vdd.t2614 7.146
R44985 vdd.n10590 vdd.t651 7.146
R44986 vdd.n10799 vdd.t2431 7.146
R44987 vdd.n10799 vdd.t2260 7.146
R44988 vdd.n10788 vdd.t2698 7.146
R44989 vdd.n10788 vdd.t2488 7.146
R44990 vdd.n10787 vdd.t1597 7.146
R44991 vdd.n10787 vdd.t2202 7.146
R44992 vdd.n10786 vdd.t1838 7.146
R44993 vdd.n10786 vdd.t2427 7.146
R44994 vdd.n10785 vdd.t2982 7.146
R44995 vdd.n10785 vdd.t592 7.146
R44996 vdd.n10784 vdd.t424 7.146
R44997 vdd.n10784 vdd.t975 7.146
R44998 vdd.n10783 vdd.t652 7.146
R44999 vdd.n10783 vdd.t1229 7.146
R45000 vdd.n10782 vdd.t1779 7.146
R45001 vdd.n10782 vdd.t2362 7.146
R45002 vdd.n10781 vdd.t1295 7.146
R45003 vdd.n10781 vdd.t1890 7.146
R45004 vdd.n10780 vdd.t2435 7.146
R45005 vdd.n10780 vdd.t31 7.146
R45006 vdd.n10779 vdd.t2863 7.146
R45007 vdd.n10779 vdd.t459 7.146
R45008 vdd.n10778 vdd.t1974 7.146
R45009 vdd.n10778 vdd.t1248 7.146
R45010 vdd.n10777 vdd.t1759 7.146
R45011 vdd.n10777 vdd.t2333 7.146
R45012 vdd.n10776 vdd.t1254 7.146
R45013 vdd.n10776 vdd.t1069 7.146
R45014 vdd.n10775 vdd.t142 7.146
R45015 vdd.n10775 vdd.t2932 7.146
R45016 vdd.n10774 vdd.t1981 7.146
R45017 vdd.n10774 vdd.t1788 7.146
R45018 vdd.n10773 vdd.t2456 7.146
R45019 vdd.n10773 vdd.t2272 7.146
R45020 vdd.n10772 vdd.t1317 7.146
R45021 vdd.n10772 vdd.t1126 7.146
R45022 vdd.n10771 vdd.t1084 7.146
R45023 vdd.n10771 vdd.t891 7.146
R45024 vdd.n10770 vdd.t678 7.146
R45025 vdd.n10770 vdd.t478 7.146
R45026 vdd.n10979 vdd.t2270 7.146
R45027 vdd.n10979 vdd.t1062 7.146
R45028 vdd.n10968 vdd.t2507 7.146
R45029 vdd.n10968 vdd.t1296 7.146
R45030 vdd.n10967 vdd.t2171 7.146
R45031 vdd.n10967 vdd.t522 7.146
R45032 vdd.n10966 vdd.t2404 7.146
R45033 vdd.n10966 vdd.t771 7.146
R45034 vdd.n10965 vdd.t568 7.146
R45035 vdd.n10965 vdd.t1887 7.146
R45036 vdd.n10964 vdd.t953 7.146
R45037 vdd.n10964 vdd.t2300 7.146
R45038 vdd.n10963 vdd.t1209 7.146
R45039 vdd.n10963 vdd.t2549 7.146
R45040 vdd.n10962 vdd.t2338 7.146
R45041 vdd.n10962 vdd.t704 7.146
R45042 vdd.n10961 vdd.t1865 7.146
R45043 vdd.n10961 vdd.t225 7.146
R45044 vdd.n10960 vdd.t6 7.146
R45045 vdd.n10960 vdd.t1336 7.146
R45046 vdd.n10959 vdd.t441 7.146
R45047 vdd.n10959 vdd.t1762 7.146
R45048 vdd.n10958 vdd.t1353 7.146
R45049 vdd.n10958 vdd.t2850 7.146
R45050 vdd.n10957 vdd.t2316 7.146
R45051 vdd.n10957 vdd.t666 7.146
R45052 vdd.n10956 vdd.t1092 7.146
R45053 vdd.n10956 vdd.t2890 7.146
R45054 vdd.n10955 vdd.t2955 7.146
R45055 vdd.n10955 vdd.t1744 7.146
R45056 vdd.n10954 vdd.t1804 7.146
R45057 vdd.n10954 vdd.t618 7.146
R45058 vdd.n10953 vdd.t2289 7.146
R45059 vdd.n10953 vdd.t1086 7.146
R45060 vdd.n10952 vdd.t1143 7.146
R45061 vdd.n10952 vdd.t2947 7.146
R45062 vdd.n10951 vdd.t902 7.146
R45063 vdd.n10951 vdd.t2720 7.146
R45064 vdd.n10950 vdd.t500 7.146
R45065 vdd.n10950 vdd.t2286 7.146
R45066 vdd.n11159 vdd.t767 7.146
R45067 vdd.n11159 vdd.t2881 7.146
R45068 vdd.n11148 vdd.t973 7.146
R45069 vdd.n11148 vdd.t137 7.146
R45070 vdd.n11147 vdd.t1499 7.146
R45071 vdd.n11147 vdd.t1817 7.146
R45072 vdd.n11146 vdd.t1749 7.146
R45073 vdd.n11146 vdd.t2079 7.146
R45074 vdd.n11145 vdd.t2896 7.146
R45075 vdd.n11145 vdd.t224 7.146
R45076 vdd.n11144 vdd.t312 7.146
R45077 vdd.n11144 vdd.t629 7.146
R45078 vdd.n11143 vdd.t555 7.146
R45079 vdd.n11143 vdd.t861 7.146
R45080 vdd.n11142 vdd.t1673 7.146
R45081 vdd.n11142 vdd.t2002 7.146
R45082 vdd.n11141 vdd.t1199 7.146
R45083 vdd.n11141 vdd.t1517 7.146
R45084 vdd.n11140 vdd.t2326 7.146
R45085 vdd.n11140 vdd.t2662 7.146
R45086 vdd.n11139 vdd.t2766 7.146
R45087 vdd.n11139 vdd.t92 7.146
R45088 vdd.n11138 vdd.t2208 7.146
R45089 vdd.n11138 vdd.t1442 7.146
R45090 vdd.n11137 vdd.t1645 7.146
R45091 vdd.n11137 vdd.t1969 7.146
R45092 vdd.n11136 vdd.t2574 7.146
R45093 vdd.n11136 vdd.t1689 7.146
R45094 vdd.n11135 vdd.t1417 7.146
R45095 vdd.n11135 vdd.t576 7.146
R45096 vdd.n11134 vdd.t301 7.146
R45097 vdd.n11134 vdd.t2409 7.146
R45098 vdd.n11133 vdd.t787 7.146
R45099 vdd.n11133 vdd.t2906 7.146
R45100 vdd.n11132 vdd.t2631 7.146
R45101 vdd.n11132 vdd.t1763 7.146
R45102 vdd.n11131 vdd.t2378 7.146
R45103 vdd.n11131 vdd.t1508 7.146
R45104 vdd.n11130 vdd.t1959 7.146
R45105 vdd.n11130 vdd.t1101 7.146
R45106 vdd.n11339 vdd.t2564 7.146
R45107 vdd.n11339 vdd.t1945 7.146
R45108 vdd.n11328 vdd.t2796 7.146
R45109 vdd.n11328 vdd.t2205 7.146
R45110 vdd.n11327 vdd.t2817 7.146
R45111 vdd.n11327 vdd.t181 7.146
R45112 vdd.n11326 vdd.t73 7.146
R45113 vdd.n11326 vdd.t430 7.146
R45114 vdd.n11325 vdd.t1195 7.146
R45115 vdd.n11325 vdd.t1544 7.146
R45116 vdd.n11324 vdd.t1609 7.146
R45117 vdd.n11324 vdd.t1953 7.146
R45118 vdd.n11323 vdd.t1852 7.146
R45119 vdd.n11323 vdd.t2213 7.146
R45120 vdd.n11322 vdd.t2995 7.146
R45121 vdd.n11322 vdd.t353 7.146
R45122 vdd.n11321 vdd.t2511 7.146
R45123 vdd.n11321 vdd.t2872 7.146
R45124 vdd.n11320 vdd.t663 7.146
R45125 vdd.n11320 vdd.t988 7.146
R45126 vdd.n11319 vdd.t1075 7.146
R45127 vdd.n11319 vdd.t1410 7.146
R45128 vdd.n11318 vdd.t810 7.146
R45129 vdd.n11318 vdd.t728 7.146
R45130 vdd.n11317 vdd.t2968 7.146
R45131 vdd.n11317 vdd.t328 7.146
R45132 vdd.n11316 vdd.t1377 7.146
R45133 vdd.n11316 vdd.t791 7.146
R45134 vdd.n11315 vdd.t258 7.146
R45135 vdd.n11315 vdd.t2636 7.146
R45136 vdd.n11314 vdd.t2101 7.146
R45137 vdd.n11314 vdd.t1485 7.146
R45138 vdd.n11313 vdd.t2589 7.146
R45139 vdd.n11313 vdd.t1965 7.146
R45140 vdd.n11312 vdd.t1431 7.146
R45141 vdd.n11312 vdd.t837 7.146
R45142 vdd.n11311 vdd.t1194 7.146
R45143 vdd.n11311 vdd.t607 7.146
R45144 vdd.n11310 vdd.t796 7.146
R45145 vdd.n11310 vdd.t192 7.146
R45146 vdd.n11415 vdd.t782 7.146
R45147 vdd.n11411 vdd.t996 7.146
R45148 vdd.n11408 vdd.t1471 7.146
R45149 vdd.n11405 vdd.t1725 7.146
R45150 vdd.n11402 vdd.t2868 7.146
R45151 vdd.n11399 vdd.t295 7.146
R45152 vdd.n11396 vdd.t527 7.146
R45153 vdd.n11393 vdd.t1647 7.146
R45154 vdd.n11390 vdd.t1176 7.146
R45155 vdd.n11387 vdd.t2314 7.146
R45156 vdd.n11386 vdd.t2747 7.146
R45157 vdd.n11383 vdd.t2301 7.146
R45158 vdd.n11380 vdd.t1629 7.146
R45159 vdd.n11377 vdd.t2592 7.146
R45160 vdd.n11374 vdd.t1435 7.146
R45161 vdd.n11371 vdd.t319 7.146
R45162 vdd.n11368 vdd.t798 7.146
R45163 vdd.n11365 vdd.t2650 7.146
R45164 vdd.n11362 vdd.t2394 7.146
R45165 vdd.n11359 vdd.t1982 7.146
R45166 vdd.n13506 vdd.n13505 0.261
R45167 vdd.n11387 vdd.n11386 0.261
R45168 vdd.n13535 vdd.n13534 0.2
R45169 vdd.n11416 vdd.n11415 0.197
R45170 vdd.n13458 vdd.n13447 0.151
R45171 vdd.n13447 vdd.n13446 0.151
R45172 vdd.n13446 vdd.n13445 0.151
R45173 vdd.n13445 vdd.n13444 0.151
R45174 vdd.n13444 vdd.n13443 0.151
R45175 vdd.n13443 vdd.n13442 0.151
R45176 vdd.n13442 vdd.n13441 0.151
R45177 vdd.n13441 vdd.n13440 0.151
R45178 vdd.n13440 vdd.n13439 0.151
R45179 vdd.n13439 vdd.n13438 0.151
R45180 vdd.n13438 vdd.n13437 0.151
R45181 vdd.n13437 vdd.n13436 0.151
R45182 vdd.n13436 vdd.n13435 0.151
R45183 vdd.n13435 vdd.n13434 0.151
R45184 vdd.n13434 vdd.n13433 0.151
R45185 vdd.n13433 vdd.n13432 0.151
R45186 vdd.n13432 vdd.n13431 0.151
R45187 vdd.n13431 vdd.n13430 0.151
R45188 vdd.n13430 vdd.n13429 0.151
R45189 vdd.n13278 vdd.n13267 0.151
R45190 vdd.n13267 vdd.n13266 0.151
R45191 vdd.n13266 vdd.n13265 0.151
R45192 vdd.n13265 vdd.n13264 0.151
R45193 vdd.n13264 vdd.n13263 0.151
R45194 vdd.n13263 vdd.n13262 0.151
R45195 vdd.n13262 vdd.n13261 0.151
R45196 vdd.n13261 vdd.n13260 0.151
R45197 vdd.n13260 vdd.n13259 0.151
R45198 vdd.n13259 vdd.n13258 0.151
R45199 vdd.n13258 vdd.n13257 0.151
R45200 vdd.n13257 vdd.n13256 0.151
R45201 vdd.n13256 vdd.n13255 0.151
R45202 vdd.n13255 vdd.n13254 0.151
R45203 vdd.n13254 vdd.n13253 0.151
R45204 vdd.n13253 vdd.n13252 0.151
R45205 vdd.n13252 vdd.n13251 0.151
R45206 vdd.n13251 vdd.n13250 0.151
R45207 vdd.n13250 vdd.n13249 0.151
R45208 vdd.n13098 vdd.n13087 0.151
R45209 vdd.n13087 vdd.n13086 0.151
R45210 vdd.n13086 vdd.n13085 0.151
R45211 vdd.n13085 vdd.n13084 0.151
R45212 vdd.n13084 vdd.n13083 0.151
R45213 vdd.n13083 vdd.n13082 0.151
R45214 vdd.n13082 vdd.n13081 0.151
R45215 vdd.n13081 vdd.n13080 0.151
R45216 vdd.n13080 vdd.n13079 0.151
R45217 vdd.n13079 vdd.n13078 0.151
R45218 vdd.n13078 vdd.n13077 0.151
R45219 vdd.n13077 vdd.n13076 0.151
R45220 vdd.n13076 vdd.n13075 0.151
R45221 vdd.n13075 vdd.n13074 0.151
R45222 vdd.n13074 vdd.n13073 0.151
R45223 vdd.n13073 vdd.n13072 0.151
R45224 vdd.n13072 vdd.n13071 0.151
R45225 vdd.n13071 vdd.n13070 0.151
R45226 vdd.n13070 vdd.n13069 0.151
R45227 vdd.n12918 vdd.n12907 0.151
R45228 vdd.n12907 vdd.n12906 0.151
R45229 vdd.n12906 vdd.n12905 0.151
R45230 vdd.n12905 vdd.n12904 0.151
R45231 vdd.n12904 vdd.n12903 0.151
R45232 vdd.n12903 vdd.n12902 0.151
R45233 vdd.n12902 vdd.n12901 0.151
R45234 vdd.n12901 vdd.n12900 0.151
R45235 vdd.n12900 vdd.n12899 0.151
R45236 vdd.n12899 vdd.n12898 0.151
R45237 vdd.n12898 vdd.n12897 0.151
R45238 vdd.n12897 vdd.n12896 0.151
R45239 vdd.n12896 vdd.n12895 0.151
R45240 vdd.n12895 vdd.n12894 0.151
R45241 vdd.n12894 vdd.n12893 0.151
R45242 vdd.n12893 vdd.n12892 0.151
R45243 vdd.n12892 vdd.n12891 0.151
R45244 vdd.n12891 vdd.n12890 0.151
R45245 vdd.n12890 vdd.n12889 0.151
R45246 vdd.n12738 vdd.n12727 0.151
R45247 vdd.n12727 vdd.n12726 0.151
R45248 vdd.n12726 vdd.n12725 0.151
R45249 vdd.n12725 vdd.n12724 0.151
R45250 vdd.n12724 vdd.n12723 0.151
R45251 vdd.n12723 vdd.n12722 0.151
R45252 vdd.n12722 vdd.n12721 0.151
R45253 vdd.n12721 vdd.n12720 0.151
R45254 vdd.n12720 vdd.n12719 0.151
R45255 vdd.n12719 vdd.n12718 0.151
R45256 vdd.n12718 vdd.n12717 0.151
R45257 vdd.n12717 vdd.n12716 0.151
R45258 vdd.n12716 vdd.n12715 0.151
R45259 vdd.n12715 vdd.n12714 0.151
R45260 vdd.n12714 vdd.n12713 0.151
R45261 vdd.n12713 vdd.n12712 0.151
R45262 vdd.n12712 vdd.n12711 0.151
R45263 vdd.n12711 vdd.n12710 0.151
R45264 vdd.n12710 vdd.n12709 0.151
R45265 vdd.n12558 vdd.n12547 0.151
R45266 vdd.n12547 vdd.n12546 0.151
R45267 vdd.n12546 vdd.n12545 0.151
R45268 vdd.n12545 vdd.n12544 0.151
R45269 vdd.n12544 vdd.n12543 0.151
R45270 vdd.n12543 vdd.n12542 0.151
R45271 vdd.n12542 vdd.n12541 0.151
R45272 vdd.n12541 vdd.n12540 0.151
R45273 vdd.n12540 vdd.n12539 0.151
R45274 vdd.n12539 vdd.n12538 0.151
R45275 vdd.n12538 vdd.n12537 0.151
R45276 vdd.n12537 vdd.n12536 0.151
R45277 vdd.n12536 vdd.n12535 0.151
R45278 vdd.n12535 vdd.n12534 0.151
R45279 vdd.n12534 vdd.n12533 0.151
R45280 vdd.n12533 vdd.n12532 0.151
R45281 vdd.n12532 vdd.n12531 0.151
R45282 vdd.n12531 vdd.n12530 0.151
R45283 vdd.n12530 vdd.n12529 0.151
R45284 vdd.n12378 vdd.n12367 0.151
R45285 vdd.n12367 vdd.n12366 0.151
R45286 vdd.n12366 vdd.n12365 0.151
R45287 vdd.n12365 vdd.n12364 0.151
R45288 vdd.n12364 vdd.n12363 0.151
R45289 vdd.n12363 vdd.n12362 0.151
R45290 vdd.n12362 vdd.n12361 0.151
R45291 vdd.n12361 vdd.n12360 0.151
R45292 vdd.n12360 vdd.n12359 0.151
R45293 vdd.n12359 vdd.n12358 0.151
R45294 vdd.n12358 vdd.n12357 0.151
R45295 vdd.n12357 vdd.n12356 0.151
R45296 vdd.n12356 vdd.n12355 0.151
R45297 vdd.n12355 vdd.n12354 0.151
R45298 vdd.n12354 vdd.n12353 0.151
R45299 vdd.n12353 vdd.n12352 0.151
R45300 vdd.n12352 vdd.n12351 0.151
R45301 vdd.n12351 vdd.n12350 0.151
R45302 vdd.n12350 vdd.n12349 0.151
R45303 vdd.n12198 vdd.n12187 0.151
R45304 vdd.n12187 vdd.n12186 0.151
R45305 vdd.n12186 vdd.n12185 0.151
R45306 vdd.n12185 vdd.n12184 0.151
R45307 vdd.n12184 vdd.n12183 0.151
R45308 vdd.n12183 vdd.n12182 0.151
R45309 vdd.n12182 vdd.n12181 0.151
R45310 vdd.n12181 vdd.n12180 0.151
R45311 vdd.n12180 vdd.n12179 0.151
R45312 vdd.n12179 vdd.n12178 0.151
R45313 vdd.n12178 vdd.n12177 0.151
R45314 vdd.n12177 vdd.n12176 0.151
R45315 vdd.n12176 vdd.n12175 0.151
R45316 vdd.n12175 vdd.n12174 0.151
R45317 vdd.n12174 vdd.n12173 0.151
R45318 vdd.n12173 vdd.n12172 0.151
R45319 vdd.n12172 vdd.n12171 0.151
R45320 vdd.n12171 vdd.n12170 0.151
R45321 vdd.n12170 vdd.n12169 0.151
R45322 vdd.n12018 vdd.n12007 0.151
R45323 vdd.n12007 vdd.n12006 0.151
R45324 vdd.n12006 vdd.n12005 0.151
R45325 vdd.n12005 vdd.n12004 0.151
R45326 vdd.n12004 vdd.n12003 0.151
R45327 vdd.n12003 vdd.n12002 0.151
R45328 vdd.n12002 vdd.n12001 0.151
R45329 vdd.n12001 vdd.n12000 0.151
R45330 vdd.n12000 vdd.n11999 0.151
R45331 vdd.n11999 vdd.n11998 0.151
R45332 vdd.n11998 vdd.n11997 0.151
R45333 vdd.n11997 vdd.n11996 0.151
R45334 vdd.n11996 vdd.n11995 0.151
R45335 vdd.n11995 vdd.n11994 0.151
R45336 vdd.n11994 vdd.n11993 0.151
R45337 vdd.n11993 vdd.n11992 0.151
R45338 vdd.n11992 vdd.n11991 0.151
R45339 vdd.n11991 vdd.n11990 0.151
R45340 vdd.n11990 vdd.n11989 0.151
R45341 vdd.n11838 vdd.n11827 0.151
R45342 vdd.n11827 vdd.n11826 0.151
R45343 vdd.n11826 vdd.n11825 0.151
R45344 vdd.n11825 vdd.n11824 0.151
R45345 vdd.n11824 vdd.n11823 0.151
R45346 vdd.n11823 vdd.n11822 0.151
R45347 vdd.n11822 vdd.n11821 0.151
R45348 vdd.n11821 vdd.n11820 0.151
R45349 vdd.n11820 vdd.n11819 0.151
R45350 vdd.n11819 vdd.n11818 0.151
R45351 vdd.n11818 vdd.n11817 0.151
R45352 vdd.n11817 vdd.n11816 0.151
R45353 vdd.n11816 vdd.n11815 0.151
R45354 vdd.n11815 vdd.n11814 0.151
R45355 vdd.n11814 vdd.n11813 0.151
R45356 vdd.n11813 vdd.n11812 0.151
R45357 vdd.n11812 vdd.n11811 0.151
R45358 vdd.n11811 vdd.n11810 0.151
R45359 vdd.n11810 vdd.n11809 0.151
R45360 vdd.n11658 vdd.n11647 0.151
R45361 vdd.n11647 vdd.n11646 0.151
R45362 vdd.n11646 vdd.n11645 0.151
R45363 vdd.n11645 vdd.n11644 0.151
R45364 vdd.n11644 vdd.n11643 0.151
R45365 vdd.n11643 vdd.n11642 0.151
R45366 vdd.n11642 vdd.n11641 0.151
R45367 vdd.n11641 vdd.n11640 0.151
R45368 vdd.n11640 vdd.n11639 0.151
R45369 vdd.n11639 vdd.n11638 0.151
R45370 vdd.n11638 vdd.n11637 0.151
R45371 vdd.n11637 vdd.n11636 0.151
R45372 vdd.n11636 vdd.n11635 0.151
R45373 vdd.n11635 vdd.n11634 0.151
R45374 vdd.n11634 vdd.n11633 0.151
R45375 vdd.n11633 vdd.n11632 0.151
R45376 vdd.n11632 vdd.n11631 0.151
R45377 vdd.n11631 vdd.n11630 0.151
R45378 vdd.n11630 vdd.n11629 0.151
R45379 vdd.n179 vdd.n168 0.151
R45380 vdd.n168 vdd.n167 0.151
R45381 vdd.n167 vdd.n166 0.151
R45382 vdd.n166 vdd.n165 0.151
R45383 vdd.n165 vdd.n164 0.151
R45384 vdd.n164 vdd.n163 0.151
R45385 vdd.n163 vdd.n162 0.151
R45386 vdd.n162 vdd.n161 0.151
R45387 vdd.n161 vdd.n160 0.151
R45388 vdd.n160 vdd.n159 0.151
R45389 vdd.n159 vdd.n158 0.151
R45390 vdd.n158 vdd.n157 0.151
R45391 vdd.n157 vdd.n156 0.151
R45392 vdd.n156 vdd.n155 0.151
R45393 vdd.n155 vdd.n154 0.151
R45394 vdd.n154 vdd.n153 0.151
R45395 vdd.n153 vdd.n152 0.151
R45396 vdd.n152 vdd.n151 0.151
R45397 vdd.n151 vdd.n150 0.151
R45398 vdd.n359 vdd.n348 0.151
R45399 vdd.n348 vdd.n347 0.151
R45400 vdd.n347 vdd.n346 0.151
R45401 vdd.n346 vdd.n345 0.151
R45402 vdd.n345 vdd.n344 0.151
R45403 vdd.n344 vdd.n343 0.151
R45404 vdd.n343 vdd.n342 0.151
R45405 vdd.n342 vdd.n341 0.151
R45406 vdd.n341 vdd.n340 0.151
R45407 vdd.n340 vdd.n339 0.151
R45408 vdd.n339 vdd.n338 0.151
R45409 vdd.n338 vdd.n337 0.151
R45410 vdd.n337 vdd.n336 0.151
R45411 vdd.n336 vdd.n335 0.151
R45412 vdd.n335 vdd.n334 0.151
R45413 vdd.n334 vdd.n333 0.151
R45414 vdd.n333 vdd.n332 0.151
R45415 vdd.n332 vdd.n331 0.151
R45416 vdd.n331 vdd.n330 0.151
R45417 vdd.n539 vdd.n528 0.151
R45418 vdd.n528 vdd.n527 0.151
R45419 vdd.n527 vdd.n526 0.151
R45420 vdd.n526 vdd.n525 0.151
R45421 vdd.n525 vdd.n524 0.151
R45422 vdd.n524 vdd.n523 0.151
R45423 vdd.n523 vdd.n522 0.151
R45424 vdd.n522 vdd.n521 0.151
R45425 vdd.n521 vdd.n520 0.151
R45426 vdd.n520 vdd.n519 0.151
R45427 vdd.n519 vdd.n518 0.151
R45428 vdd.n518 vdd.n517 0.151
R45429 vdd.n517 vdd.n516 0.151
R45430 vdd.n516 vdd.n515 0.151
R45431 vdd.n515 vdd.n514 0.151
R45432 vdd.n514 vdd.n513 0.151
R45433 vdd.n513 vdd.n512 0.151
R45434 vdd.n512 vdd.n511 0.151
R45435 vdd.n511 vdd.n510 0.151
R45436 vdd.n719 vdd.n708 0.151
R45437 vdd.n708 vdd.n707 0.151
R45438 vdd.n707 vdd.n706 0.151
R45439 vdd.n706 vdd.n705 0.151
R45440 vdd.n705 vdd.n704 0.151
R45441 vdd.n704 vdd.n703 0.151
R45442 vdd.n703 vdd.n702 0.151
R45443 vdd.n702 vdd.n701 0.151
R45444 vdd.n701 vdd.n700 0.151
R45445 vdd.n700 vdd.n699 0.151
R45446 vdd.n699 vdd.n698 0.151
R45447 vdd.n698 vdd.n697 0.151
R45448 vdd.n697 vdd.n696 0.151
R45449 vdd.n696 vdd.n695 0.151
R45450 vdd.n695 vdd.n694 0.151
R45451 vdd.n694 vdd.n693 0.151
R45452 vdd.n693 vdd.n692 0.151
R45453 vdd.n692 vdd.n691 0.151
R45454 vdd.n691 vdd.n690 0.151
R45455 vdd.n899 vdd.n888 0.151
R45456 vdd.n888 vdd.n887 0.151
R45457 vdd.n887 vdd.n886 0.151
R45458 vdd.n886 vdd.n885 0.151
R45459 vdd.n885 vdd.n884 0.151
R45460 vdd.n884 vdd.n883 0.151
R45461 vdd.n883 vdd.n882 0.151
R45462 vdd.n882 vdd.n881 0.151
R45463 vdd.n881 vdd.n880 0.151
R45464 vdd.n880 vdd.n879 0.151
R45465 vdd.n879 vdd.n878 0.151
R45466 vdd.n878 vdd.n877 0.151
R45467 vdd.n877 vdd.n876 0.151
R45468 vdd.n876 vdd.n875 0.151
R45469 vdd.n875 vdd.n874 0.151
R45470 vdd.n874 vdd.n873 0.151
R45471 vdd.n873 vdd.n872 0.151
R45472 vdd.n872 vdd.n871 0.151
R45473 vdd.n871 vdd.n870 0.151
R45474 vdd.n1079 vdd.n1068 0.151
R45475 vdd.n1068 vdd.n1067 0.151
R45476 vdd.n1067 vdd.n1066 0.151
R45477 vdd.n1066 vdd.n1065 0.151
R45478 vdd.n1065 vdd.n1064 0.151
R45479 vdd.n1064 vdd.n1063 0.151
R45480 vdd.n1063 vdd.n1062 0.151
R45481 vdd.n1062 vdd.n1061 0.151
R45482 vdd.n1061 vdd.n1060 0.151
R45483 vdd.n1060 vdd.n1059 0.151
R45484 vdd.n1059 vdd.n1058 0.151
R45485 vdd.n1058 vdd.n1057 0.151
R45486 vdd.n1057 vdd.n1056 0.151
R45487 vdd.n1056 vdd.n1055 0.151
R45488 vdd.n1055 vdd.n1054 0.151
R45489 vdd.n1054 vdd.n1053 0.151
R45490 vdd.n1053 vdd.n1052 0.151
R45491 vdd.n1052 vdd.n1051 0.151
R45492 vdd.n1051 vdd.n1050 0.151
R45493 vdd.n1259 vdd.n1248 0.151
R45494 vdd.n1248 vdd.n1247 0.151
R45495 vdd.n1247 vdd.n1246 0.151
R45496 vdd.n1246 vdd.n1245 0.151
R45497 vdd.n1245 vdd.n1244 0.151
R45498 vdd.n1244 vdd.n1243 0.151
R45499 vdd.n1243 vdd.n1242 0.151
R45500 vdd.n1242 vdd.n1241 0.151
R45501 vdd.n1241 vdd.n1240 0.151
R45502 vdd.n1240 vdd.n1239 0.151
R45503 vdd.n1239 vdd.n1238 0.151
R45504 vdd.n1238 vdd.n1237 0.151
R45505 vdd.n1237 vdd.n1236 0.151
R45506 vdd.n1236 vdd.n1235 0.151
R45507 vdd.n1235 vdd.n1234 0.151
R45508 vdd.n1234 vdd.n1233 0.151
R45509 vdd.n1233 vdd.n1232 0.151
R45510 vdd.n1232 vdd.n1231 0.151
R45511 vdd.n1231 vdd.n1230 0.151
R45512 vdd.n1439 vdd.n1428 0.151
R45513 vdd.n1428 vdd.n1427 0.151
R45514 vdd.n1427 vdd.n1426 0.151
R45515 vdd.n1426 vdd.n1425 0.151
R45516 vdd.n1425 vdd.n1424 0.151
R45517 vdd.n1424 vdd.n1423 0.151
R45518 vdd.n1423 vdd.n1422 0.151
R45519 vdd.n1422 vdd.n1421 0.151
R45520 vdd.n1421 vdd.n1420 0.151
R45521 vdd.n1420 vdd.n1419 0.151
R45522 vdd.n1419 vdd.n1418 0.151
R45523 vdd.n1418 vdd.n1417 0.151
R45524 vdd.n1417 vdd.n1416 0.151
R45525 vdd.n1416 vdd.n1415 0.151
R45526 vdd.n1415 vdd.n1414 0.151
R45527 vdd.n1414 vdd.n1413 0.151
R45528 vdd.n1413 vdd.n1412 0.151
R45529 vdd.n1412 vdd.n1411 0.151
R45530 vdd.n1411 vdd.n1410 0.151
R45531 vdd.n1619 vdd.n1608 0.151
R45532 vdd.n1608 vdd.n1607 0.151
R45533 vdd.n1607 vdd.n1606 0.151
R45534 vdd.n1606 vdd.n1605 0.151
R45535 vdd.n1605 vdd.n1604 0.151
R45536 vdd.n1604 vdd.n1603 0.151
R45537 vdd.n1603 vdd.n1602 0.151
R45538 vdd.n1602 vdd.n1601 0.151
R45539 vdd.n1601 vdd.n1600 0.151
R45540 vdd.n1600 vdd.n1599 0.151
R45541 vdd.n1599 vdd.n1598 0.151
R45542 vdd.n1598 vdd.n1597 0.151
R45543 vdd.n1597 vdd.n1596 0.151
R45544 vdd.n1596 vdd.n1595 0.151
R45545 vdd.n1595 vdd.n1594 0.151
R45546 vdd.n1594 vdd.n1593 0.151
R45547 vdd.n1593 vdd.n1592 0.151
R45548 vdd.n1592 vdd.n1591 0.151
R45549 vdd.n1591 vdd.n1590 0.151
R45550 vdd.n1799 vdd.n1788 0.151
R45551 vdd.n1788 vdd.n1787 0.151
R45552 vdd.n1787 vdd.n1786 0.151
R45553 vdd.n1786 vdd.n1785 0.151
R45554 vdd.n1785 vdd.n1784 0.151
R45555 vdd.n1784 vdd.n1783 0.151
R45556 vdd.n1783 vdd.n1782 0.151
R45557 vdd.n1782 vdd.n1781 0.151
R45558 vdd.n1781 vdd.n1780 0.151
R45559 vdd.n1780 vdd.n1779 0.151
R45560 vdd.n1779 vdd.n1778 0.151
R45561 vdd.n1778 vdd.n1777 0.151
R45562 vdd.n1777 vdd.n1776 0.151
R45563 vdd.n1776 vdd.n1775 0.151
R45564 vdd.n1775 vdd.n1774 0.151
R45565 vdd.n1774 vdd.n1773 0.151
R45566 vdd.n1773 vdd.n1772 0.151
R45567 vdd.n1772 vdd.n1771 0.151
R45568 vdd.n1771 vdd.n1770 0.151
R45569 vdd.n1979 vdd.n1968 0.151
R45570 vdd.n1968 vdd.n1967 0.151
R45571 vdd.n1967 vdd.n1966 0.151
R45572 vdd.n1966 vdd.n1965 0.151
R45573 vdd.n1965 vdd.n1964 0.151
R45574 vdd.n1964 vdd.n1963 0.151
R45575 vdd.n1963 vdd.n1962 0.151
R45576 vdd.n1962 vdd.n1961 0.151
R45577 vdd.n1961 vdd.n1960 0.151
R45578 vdd.n1960 vdd.n1959 0.151
R45579 vdd.n1959 vdd.n1958 0.151
R45580 vdd.n1958 vdd.n1957 0.151
R45581 vdd.n1957 vdd.n1956 0.151
R45582 vdd.n1956 vdd.n1955 0.151
R45583 vdd.n1955 vdd.n1954 0.151
R45584 vdd.n1954 vdd.n1953 0.151
R45585 vdd.n1953 vdd.n1952 0.151
R45586 vdd.n1952 vdd.n1951 0.151
R45587 vdd.n1951 vdd.n1950 0.151
R45588 vdd.n2159 vdd.n2148 0.151
R45589 vdd.n2148 vdd.n2147 0.151
R45590 vdd.n2147 vdd.n2146 0.151
R45591 vdd.n2146 vdd.n2145 0.151
R45592 vdd.n2145 vdd.n2144 0.151
R45593 vdd.n2144 vdd.n2143 0.151
R45594 vdd.n2143 vdd.n2142 0.151
R45595 vdd.n2142 vdd.n2141 0.151
R45596 vdd.n2141 vdd.n2140 0.151
R45597 vdd.n2140 vdd.n2139 0.151
R45598 vdd.n2139 vdd.n2138 0.151
R45599 vdd.n2138 vdd.n2137 0.151
R45600 vdd.n2137 vdd.n2136 0.151
R45601 vdd.n2136 vdd.n2135 0.151
R45602 vdd.n2135 vdd.n2134 0.151
R45603 vdd.n2134 vdd.n2133 0.151
R45604 vdd.n2133 vdd.n2132 0.151
R45605 vdd.n2132 vdd.n2131 0.151
R45606 vdd.n2131 vdd.n2130 0.151
R45607 vdd.n2339 vdd.n2328 0.151
R45608 vdd.n2328 vdd.n2327 0.151
R45609 vdd.n2327 vdd.n2326 0.151
R45610 vdd.n2326 vdd.n2325 0.151
R45611 vdd.n2325 vdd.n2324 0.151
R45612 vdd.n2324 vdd.n2323 0.151
R45613 vdd.n2323 vdd.n2322 0.151
R45614 vdd.n2322 vdd.n2321 0.151
R45615 vdd.n2321 vdd.n2320 0.151
R45616 vdd.n2320 vdd.n2319 0.151
R45617 vdd.n2319 vdd.n2318 0.151
R45618 vdd.n2318 vdd.n2317 0.151
R45619 vdd.n2317 vdd.n2316 0.151
R45620 vdd.n2316 vdd.n2315 0.151
R45621 vdd.n2315 vdd.n2314 0.151
R45622 vdd.n2314 vdd.n2313 0.151
R45623 vdd.n2313 vdd.n2312 0.151
R45624 vdd.n2312 vdd.n2311 0.151
R45625 vdd.n2311 vdd.n2310 0.151
R45626 vdd.n2519 vdd.n2508 0.151
R45627 vdd.n2508 vdd.n2507 0.151
R45628 vdd.n2507 vdd.n2506 0.151
R45629 vdd.n2506 vdd.n2505 0.151
R45630 vdd.n2505 vdd.n2504 0.151
R45631 vdd.n2504 vdd.n2503 0.151
R45632 vdd.n2503 vdd.n2502 0.151
R45633 vdd.n2502 vdd.n2501 0.151
R45634 vdd.n2501 vdd.n2500 0.151
R45635 vdd.n2500 vdd.n2499 0.151
R45636 vdd.n2499 vdd.n2498 0.151
R45637 vdd.n2498 vdd.n2497 0.151
R45638 vdd.n2497 vdd.n2496 0.151
R45639 vdd.n2496 vdd.n2495 0.151
R45640 vdd.n2495 vdd.n2494 0.151
R45641 vdd.n2494 vdd.n2493 0.151
R45642 vdd.n2493 vdd.n2492 0.151
R45643 vdd.n2492 vdd.n2491 0.151
R45644 vdd.n2491 vdd.n2490 0.151
R45645 vdd.n2699 vdd.n2688 0.151
R45646 vdd.n2688 vdd.n2687 0.151
R45647 vdd.n2687 vdd.n2686 0.151
R45648 vdd.n2686 vdd.n2685 0.151
R45649 vdd.n2685 vdd.n2684 0.151
R45650 vdd.n2684 vdd.n2683 0.151
R45651 vdd.n2683 vdd.n2682 0.151
R45652 vdd.n2682 vdd.n2681 0.151
R45653 vdd.n2681 vdd.n2680 0.151
R45654 vdd.n2680 vdd.n2679 0.151
R45655 vdd.n2679 vdd.n2678 0.151
R45656 vdd.n2678 vdd.n2677 0.151
R45657 vdd.n2677 vdd.n2676 0.151
R45658 vdd.n2676 vdd.n2675 0.151
R45659 vdd.n2675 vdd.n2674 0.151
R45660 vdd.n2674 vdd.n2673 0.151
R45661 vdd.n2673 vdd.n2672 0.151
R45662 vdd.n2672 vdd.n2671 0.151
R45663 vdd.n2671 vdd.n2670 0.151
R45664 vdd.n2879 vdd.n2868 0.151
R45665 vdd.n2868 vdd.n2867 0.151
R45666 vdd.n2867 vdd.n2866 0.151
R45667 vdd.n2866 vdd.n2865 0.151
R45668 vdd.n2865 vdd.n2864 0.151
R45669 vdd.n2864 vdd.n2863 0.151
R45670 vdd.n2863 vdd.n2862 0.151
R45671 vdd.n2862 vdd.n2861 0.151
R45672 vdd.n2861 vdd.n2860 0.151
R45673 vdd.n2860 vdd.n2859 0.151
R45674 vdd.n2859 vdd.n2858 0.151
R45675 vdd.n2858 vdd.n2857 0.151
R45676 vdd.n2857 vdd.n2856 0.151
R45677 vdd.n2856 vdd.n2855 0.151
R45678 vdd.n2855 vdd.n2854 0.151
R45679 vdd.n2854 vdd.n2853 0.151
R45680 vdd.n2853 vdd.n2852 0.151
R45681 vdd.n2852 vdd.n2851 0.151
R45682 vdd.n2851 vdd.n2850 0.151
R45683 vdd.n3059 vdd.n3048 0.151
R45684 vdd.n3048 vdd.n3047 0.151
R45685 vdd.n3047 vdd.n3046 0.151
R45686 vdd.n3046 vdd.n3045 0.151
R45687 vdd.n3045 vdd.n3044 0.151
R45688 vdd.n3044 vdd.n3043 0.151
R45689 vdd.n3043 vdd.n3042 0.151
R45690 vdd.n3042 vdd.n3041 0.151
R45691 vdd.n3041 vdd.n3040 0.151
R45692 vdd.n3040 vdd.n3039 0.151
R45693 vdd.n3039 vdd.n3038 0.151
R45694 vdd.n3038 vdd.n3037 0.151
R45695 vdd.n3037 vdd.n3036 0.151
R45696 vdd.n3036 vdd.n3035 0.151
R45697 vdd.n3035 vdd.n3034 0.151
R45698 vdd.n3034 vdd.n3033 0.151
R45699 vdd.n3033 vdd.n3032 0.151
R45700 vdd.n3032 vdd.n3031 0.151
R45701 vdd.n3031 vdd.n3030 0.151
R45702 vdd.n3239 vdd.n3228 0.151
R45703 vdd.n3228 vdd.n3227 0.151
R45704 vdd.n3227 vdd.n3226 0.151
R45705 vdd.n3226 vdd.n3225 0.151
R45706 vdd.n3225 vdd.n3224 0.151
R45707 vdd.n3224 vdd.n3223 0.151
R45708 vdd.n3223 vdd.n3222 0.151
R45709 vdd.n3222 vdd.n3221 0.151
R45710 vdd.n3221 vdd.n3220 0.151
R45711 vdd.n3220 vdd.n3219 0.151
R45712 vdd.n3219 vdd.n3218 0.151
R45713 vdd.n3218 vdd.n3217 0.151
R45714 vdd.n3217 vdd.n3216 0.151
R45715 vdd.n3216 vdd.n3215 0.151
R45716 vdd.n3215 vdd.n3214 0.151
R45717 vdd.n3214 vdd.n3213 0.151
R45718 vdd.n3213 vdd.n3212 0.151
R45719 vdd.n3212 vdd.n3211 0.151
R45720 vdd.n3211 vdd.n3210 0.151
R45721 vdd.n3419 vdd.n3408 0.151
R45722 vdd.n3408 vdd.n3407 0.151
R45723 vdd.n3407 vdd.n3406 0.151
R45724 vdd.n3406 vdd.n3405 0.151
R45725 vdd.n3405 vdd.n3404 0.151
R45726 vdd.n3404 vdd.n3403 0.151
R45727 vdd.n3403 vdd.n3402 0.151
R45728 vdd.n3402 vdd.n3401 0.151
R45729 vdd.n3401 vdd.n3400 0.151
R45730 vdd.n3400 vdd.n3399 0.151
R45731 vdd.n3399 vdd.n3398 0.151
R45732 vdd.n3398 vdd.n3397 0.151
R45733 vdd.n3397 vdd.n3396 0.151
R45734 vdd.n3396 vdd.n3395 0.151
R45735 vdd.n3395 vdd.n3394 0.151
R45736 vdd.n3394 vdd.n3393 0.151
R45737 vdd.n3393 vdd.n3392 0.151
R45738 vdd.n3392 vdd.n3391 0.151
R45739 vdd.n3391 vdd.n3390 0.151
R45740 vdd.n3599 vdd.n3588 0.151
R45741 vdd.n3588 vdd.n3587 0.151
R45742 vdd.n3587 vdd.n3586 0.151
R45743 vdd.n3586 vdd.n3585 0.151
R45744 vdd.n3585 vdd.n3584 0.151
R45745 vdd.n3584 vdd.n3583 0.151
R45746 vdd.n3583 vdd.n3582 0.151
R45747 vdd.n3582 vdd.n3581 0.151
R45748 vdd.n3581 vdd.n3580 0.151
R45749 vdd.n3580 vdd.n3579 0.151
R45750 vdd.n3579 vdd.n3578 0.151
R45751 vdd.n3578 vdd.n3577 0.151
R45752 vdd.n3577 vdd.n3576 0.151
R45753 vdd.n3576 vdd.n3575 0.151
R45754 vdd.n3575 vdd.n3574 0.151
R45755 vdd.n3574 vdd.n3573 0.151
R45756 vdd.n3573 vdd.n3572 0.151
R45757 vdd.n3572 vdd.n3571 0.151
R45758 vdd.n3571 vdd.n3570 0.151
R45759 vdd.n3779 vdd.n3768 0.151
R45760 vdd.n3768 vdd.n3767 0.151
R45761 vdd.n3767 vdd.n3766 0.151
R45762 vdd.n3766 vdd.n3765 0.151
R45763 vdd.n3765 vdd.n3764 0.151
R45764 vdd.n3764 vdd.n3763 0.151
R45765 vdd.n3763 vdd.n3762 0.151
R45766 vdd.n3762 vdd.n3761 0.151
R45767 vdd.n3761 vdd.n3760 0.151
R45768 vdd.n3760 vdd.n3759 0.151
R45769 vdd.n3759 vdd.n3758 0.151
R45770 vdd.n3758 vdd.n3757 0.151
R45771 vdd.n3757 vdd.n3756 0.151
R45772 vdd.n3756 vdd.n3755 0.151
R45773 vdd.n3755 vdd.n3754 0.151
R45774 vdd.n3754 vdd.n3753 0.151
R45775 vdd.n3753 vdd.n3752 0.151
R45776 vdd.n3752 vdd.n3751 0.151
R45777 vdd.n3751 vdd.n3750 0.151
R45778 vdd.n3959 vdd.n3948 0.151
R45779 vdd.n3948 vdd.n3947 0.151
R45780 vdd.n3947 vdd.n3946 0.151
R45781 vdd.n3946 vdd.n3945 0.151
R45782 vdd.n3945 vdd.n3944 0.151
R45783 vdd.n3944 vdd.n3943 0.151
R45784 vdd.n3943 vdd.n3942 0.151
R45785 vdd.n3942 vdd.n3941 0.151
R45786 vdd.n3941 vdd.n3940 0.151
R45787 vdd.n3940 vdd.n3939 0.151
R45788 vdd.n3939 vdd.n3938 0.151
R45789 vdd.n3938 vdd.n3937 0.151
R45790 vdd.n3937 vdd.n3936 0.151
R45791 vdd.n3936 vdd.n3935 0.151
R45792 vdd.n3935 vdd.n3934 0.151
R45793 vdd.n3934 vdd.n3933 0.151
R45794 vdd.n3933 vdd.n3932 0.151
R45795 vdd.n3932 vdd.n3931 0.151
R45796 vdd.n3931 vdd.n3930 0.151
R45797 vdd.n4139 vdd.n4128 0.151
R45798 vdd.n4128 vdd.n4127 0.151
R45799 vdd.n4127 vdd.n4126 0.151
R45800 vdd.n4126 vdd.n4125 0.151
R45801 vdd.n4125 vdd.n4124 0.151
R45802 vdd.n4124 vdd.n4123 0.151
R45803 vdd.n4123 vdd.n4122 0.151
R45804 vdd.n4122 vdd.n4121 0.151
R45805 vdd.n4121 vdd.n4120 0.151
R45806 vdd.n4120 vdd.n4119 0.151
R45807 vdd.n4119 vdd.n4118 0.151
R45808 vdd.n4118 vdd.n4117 0.151
R45809 vdd.n4117 vdd.n4116 0.151
R45810 vdd.n4116 vdd.n4115 0.151
R45811 vdd.n4115 vdd.n4114 0.151
R45812 vdd.n4114 vdd.n4113 0.151
R45813 vdd.n4113 vdd.n4112 0.151
R45814 vdd.n4112 vdd.n4111 0.151
R45815 vdd.n4111 vdd.n4110 0.151
R45816 vdd.n4319 vdd.n4308 0.151
R45817 vdd.n4308 vdd.n4307 0.151
R45818 vdd.n4307 vdd.n4306 0.151
R45819 vdd.n4306 vdd.n4305 0.151
R45820 vdd.n4305 vdd.n4304 0.151
R45821 vdd.n4304 vdd.n4303 0.151
R45822 vdd.n4303 vdd.n4302 0.151
R45823 vdd.n4302 vdd.n4301 0.151
R45824 vdd.n4301 vdd.n4300 0.151
R45825 vdd.n4300 vdd.n4299 0.151
R45826 vdd.n4299 vdd.n4298 0.151
R45827 vdd.n4298 vdd.n4297 0.151
R45828 vdd.n4297 vdd.n4296 0.151
R45829 vdd.n4296 vdd.n4295 0.151
R45830 vdd.n4295 vdd.n4294 0.151
R45831 vdd.n4294 vdd.n4293 0.151
R45832 vdd.n4293 vdd.n4292 0.151
R45833 vdd.n4292 vdd.n4291 0.151
R45834 vdd.n4291 vdd.n4290 0.151
R45835 vdd.n4499 vdd.n4488 0.151
R45836 vdd.n4488 vdd.n4487 0.151
R45837 vdd.n4487 vdd.n4486 0.151
R45838 vdd.n4486 vdd.n4485 0.151
R45839 vdd.n4485 vdd.n4484 0.151
R45840 vdd.n4484 vdd.n4483 0.151
R45841 vdd.n4483 vdd.n4482 0.151
R45842 vdd.n4482 vdd.n4481 0.151
R45843 vdd.n4481 vdd.n4480 0.151
R45844 vdd.n4480 vdd.n4479 0.151
R45845 vdd.n4479 vdd.n4478 0.151
R45846 vdd.n4478 vdd.n4477 0.151
R45847 vdd.n4477 vdd.n4476 0.151
R45848 vdd.n4476 vdd.n4475 0.151
R45849 vdd.n4475 vdd.n4474 0.151
R45850 vdd.n4474 vdd.n4473 0.151
R45851 vdd.n4473 vdd.n4472 0.151
R45852 vdd.n4472 vdd.n4471 0.151
R45853 vdd.n4471 vdd.n4470 0.151
R45854 vdd.n4679 vdd.n4668 0.151
R45855 vdd.n4668 vdd.n4667 0.151
R45856 vdd.n4667 vdd.n4666 0.151
R45857 vdd.n4666 vdd.n4665 0.151
R45858 vdd.n4665 vdd.n4664 0.151
R45859 vdd.n4664 vdd.n4663 0.151
R45860 vdd.n4663 vdd.n4662 0.151
R45861 vdd.n4662 vdd.n4661 0.151
R45862 vdd.n4661 vdd.n4660 0.151
R45863 vdd.n4660 vdd.n4659 0.151
R45864 vdd.n4659 vdd.n4658 0.151
R45865 vdd.n4658 vdd.n4657 0.151
R45866 vdd.n4657 vdd.n4656 0.151
R45867 vdd.n4656 vdd.n4655 0.151
R45868 vdd.n4655 vdd.n4654 0.151
R45869 vdd.n4654 vdd.n4653 0.151
R45870 vdd.n4653 vdd.n4652 0.151
R45871 vdd.n4652 vdd.n4651 0.151
R45872 vdd.n4651 vdd.n4650 0.151
R45873 vdd.n4859 vdd.n4848 0.151
R45874 vdd.n4848 vdd.n4847 0.151
R45875 vdd.n4847 vdd.n4846 0.151
R45876 vdd.n4846 vdd.n4845 0.151
R45877 vdd.n4845 vdd.n4844 0.151
R45878 vdd.n4844 vdd.n4843 0.151
R45879 vdd.n4843 vdd.n4842 0.151
R45880 vdd.n4842 vdd.n4841 0.151
R45881 vdd.n4841 vdd.n4840 0.151
R45882 vdd.n4840 vdd.n4839 0.151
R45883 vdd.n4839 vdd.n4838 0.151
R45884 vdd.n4838 vdd.n4837 0.151
R45885 vdd.n4837 vdd.n4836 0.151
R45886 vdd.n4836 vdd.n4835 0.151
R45887 vdd.n4835 vdd.n4834 0.151
R45888 vdd.n4834 vdd.n4833 0.151
R45889 vdd.n4833 vdd.n4832 0.151
R45890 vdd.n4832 vdd.n4831 0.151
R45891 vdd.n4831 vdd.n4830 0.151
R45892 vdd.n5039 vdd.n5028 0.151
R45893 vdd.n5028 vdd.n5027 0.151
R45894 vdd.n5027 vdd.n5026 0.151
R45895 vdd.n5026 vdd.n5025 0.151
R45896 vdd.n5025 vdd.n5024 0.151
R45897 vdd.n5024 vdd.n5023 0.151
R45898 vdd.n5023 vdd.n5022 0.151
R45899 vdd.n5022 vdd.n5021 0.151
R45900 vdd.n5021 vdd.n5020 0.151
R45901 vdd.n5020 vdd.n5019 0.151
R45902 vdd.n5019 vdd.n5018 0.151
R45903 vdd.n5018 vdd.n5017 0.151
R45904 vdd.n5017 vdd.n5016 0.151
R45905 vdd.n5016 vdd.n5015 0.151
R45906 vdd.n5015 vdd.n5014 0.151
R45907 vdd.n5014 vdd.n5013 0.151
R45908 vdd.n5013 vdd.n5012 0.151
R45909 vdd.n5012 vdd.n5011 0.151
R45910 vdd.n5011 vdd.n5010 0.151
R45911 vdd.n5219 vdd.n5208 0.151
R45912 vdd.n5208 vdd.n5207 0.151
R45913 vdd.n5207 vdd.n5206 0.151
R45914 vdd.n5206 vdd.n5205 0.151
R45915 vdd.n5205 vdd.n5204 0.151
R45916 vdd.n5204 vdd.n5203 0.151
R45917 vdd.n5203 vdd.n5202 0.151
R45918 vdd.n5202 vdd.n5201 0.151
R45919 vdd.n5201 vdd.n5200 0.151
R45920 vdd.n5200 vdd.n5199 0.151
R45921 vdd.n5199 vdd.n5198 0.151
R45922 vdd.n5198 vdd.n5197 0.151
R45923 vdd.n5197 vdd.n5196 0.151
R45924 vdd.n5196 vdd.n5195 0.151
R45925 vdd.n5195 vdd.n5194 0.151
R45926 vdd.n5194 vdd.n5193 0.151
R45927 vdd.n5193 vdd.n5192 0.151
R45928 vdd.n5192 vdd.n5191 0.151
R45929 vdd.n5191 vdd.n5190 0.151
R45930 vdd.n5399 vdd.n5388 0.151
R45931 vdd.n5388 vdd.n5387 0.151
R45932 vdd.n5387 vdd.n5386 0.151
R45933 vdd.n5386 vdd.n5385 0.151
R45934 vdd.n5385 vdd.n5384 0.151
R45935 vdd.n5384 vdd.n5383 0.151
R45936 vdd.n5383 vdd.n5382 0.151
R45937 vdd.n5382 vdd.n5381 0.151
R45938 vdd.n5381 vdd.n5380 0.151
R45939 vdd.n5380 vdd.n5379 0.151
R45940 vdd.n5379 vdd.n5378 0.151
R45941 vdd.n5378 vdd.n5377 0.151
R45942 vdd.n5377 vdd.n5376 0.151
R45943 vdd.n5376 vdd.n5375 0.151
R45944 vdd.n5375 vdd.n5374 0.151
R45945 vdd.n5374 vdd.n5373 0.151
R45946 vdd.n5373 vdd.n5372 0.151
R45947 vdd.n5372 vdd.n5371 0.151
R45948 vdd.n5371 vdd.n5370 0.151
R45949 vdd.n5579 vdd.n5568 0.151
R45950 vdd.n5568 vdd.n5567 0.151
R45951 vdd.n5567 vdd.n5566 0.151
R45952 vdd.n5566 vdd.n5565 0.151
R45953 vdd.n5565 vdd.n5564 0.151
R45954 vdd.n5564 vdd.n5563 0.151
R45955 vdd.n5563 vdd.n5562 0.151
R45956 vdd.n5562 vdd.n5561 0.151
R45957 vdd.n5561 vdd.n5560 0.151
R45958 vdd.n5560 vdd.n5559 0.151
R45959 vdd.n5559 vdd.n5558 0.151
R45960 vdd.n5558 vdd.n5557 0.151
R45961 vdd.n5557 vdd.n5556 0.151
R45962 vdd.n5556 vdd.n5555 0.151
R45963 vdd.n5555 vdd.n5554 0.151
R45964 vdd.n5554 vdd.n5553 0.151
R45965 vdd.n5553 vdd.n5552 0.151
R45966 vdd.n5552 vdd.n5551 0.151
R45967 vdd.n5551 vdd.n5550 0.151
R45968 vdd.n5759 vdd.n5748 0.151
R45969 vdd.n5748 vdd.n5747 0.151
R45970 vdd.n5747 vdd.n5746 0.151
R45971 vdd.n5746 vdd.n5745 0.151
R45972 vdd.n5745 vdd.n5744 0.151
R45973 vdd.n5744 vdd.n5743 0.151
R45974 vdd.n5743 vdd.n5742 0.151
R45975 vdd.n5742 vdd.n5741 0.151
R45976 vdd.n5741 vdd.n5740 0.151
R45977 vdd.n5740 vdd.n5739 0.151
R45978 vdd.n5739 vdd.n5738 0.151
R45979 vdd.n5738 vdd.n5737 0.151
R45980 vdd.n5737 vdd.n5736 0.151
R45981 vdd.n5736 vdd.n5735 0.151
R45982 vdd.n5735 vdd.n5734 0.151
R45983 vdd.n5734 vdd.n5733 0.151
R45984 vdd.n5733 vdd.n5732 0.151
R45985 vdd.n5732 vdd.n5731 0.151
R45986 vdd.n5731 vdd.n5730 0.151
R45987 vdd.n5939 vdd.n5928 0.151
R45988 vdd.n5928 vdd.n5927 0.151
R45989 vdd.n5927 vdd.n5926 0.151
R45990 vdd.n5926 vdd.n5925 0.151
R45991 vdd.n5925 vdd.n5924 0.151
R45992 vdd.n5924 vdd.n5923 0.151
R45993 vdd.n5923 vdd.n5922 0.151
R45994 vdd.n5922 vdd.n5921 0.151
R45995 vdd.n5921 vdd.n5920 0.151
R45996 vdd.n5920 vdd.n5919 0.151
R45997 vdd.n5919 vdd.n5918 0.151
R45998 vdd.n5918 vdd.n5917 0.151
R45999 vdd.n5917 vdd.n5916 0.151
R46000 vdd.n5916 vdd.n5915 0.151
R46001 vdd.n5915 vdd.n5914 0.151
R46002 vdd.n5914 vdd.n5913 0.151
R46003 vdd.n5913 vdd.n5912 0.151
R46004 vdd.n5912 vdd.n5911 0.151
R46005 vdd.n5911 vdd.n5910 0.151
R46006 vdd.n6119 vdd.n6108 0.151
R46007 vdd.n6108 vdd.n6107 0.151
R46008 vdd.n6107 vdd.n6106 0.151
R46009 vdd.n6106 vdd.n6105 0.151
R46010 vdd.n6105 vdd.n6104 0.151
R46011 vdd.n6104 vdd.n6103 0.151
R46012 vdd.n6103 vdd.n6102 0.151
R46013 vdd.n6102 vdd.n6101 0.151
R46014 vdd.n6101 vdd.n6100 0.151
R46015 vdd.n6100 vdd.n6099 0.151
R46016 vdd.n6099 vdd.n6098 0.151
R46017 vdd.n6098 vdd.n6097 0.151
R46018 vdd.n6097 vdd.n6096 0.151
R46019 vdd.n6096 vdd.n6095 0.151
R46020 vdd.n6095 vdd.n6094 0.151
R46021 vdd.n6094 vdd.n6093 0.151
R46022 vdd.n6093 vdd.n6092 0.151
R46023 vdd.n6092 vdd.n6091 0.151
R46024 vdd.n6091 vdd.n6090 0.151
R46025 vdd.n6299 vdd.n6288 0.151
R46026 vdd.n6288 vdd.n6287 0.151
R46027 vdd.n6287 vdd.n6286 0.151
R46028 vdd.n6286 vdd.n6285 0.151
R46029 vdd.n6285 vdd.n6284 0.151
R46030 vdd.n6284 vdd.n6283 0.151
R46031 vdd.n6283 vdd.n6282 0.151
R46032 vdd.n6282 vdd.n6281 0.151
R46033 vdd.n6281 vdd.n6280 0.151
R46034 vdd.n6280 vdd.n6279 0.151
R46035 vdd.n6279 vdd.n6278 0.151
R46036 vdd.n6278 vdd.n6277 0.151
R46037 vdd.n6277 vdd.n6276 0.151
R46038 vdd.n6276 vdd.n6275 0.151
R46039 vdd.n6275 vdd.n6274 0.151
R46040 vdd.n6274 vdd.n6273 0.151
R46041 vdd.n6273 vdd.n6272 0.151
R46042 vdd.n6272 vdd.n6271 0.151
R46043 vdd.n6271 vdd.n6270 0.151
R46044 vdd.n6479 vdd.n6468 0.151
R46045 vdd.n6468 vdd.n6467 0.151
R46046 vdd.n6467 vdd.n6466 0.151
R46047 vdd.n6466 vdd.n6465 0.151
R46048 vdd.n6465 vdd.n6464 0.151
R46049 vdd.n6464 vdd.n6463 0.151
R46050 vdd.n6463 vdd.n6462 0.151
R46051 vdd.n6462 vdd.n6461 0.151
R46052 vdd.n6461 vdd.n6460 0.151
R46053 vdd.n6460 vdd.n6459 0.151
R46054 vdd.n6459 vdd.n6458 0.151
R46055 vdd.n6458 vdd.n6457 0.151
R46056 vdd.n6457 vdd.n6456 0.151
R46057 vdd.n6456 vdd.n6455 0.151
R46058 vdd.n6455 vdd.n6454 0.151
R46059 vdd.n6454 vdd.n6453 0.151
R46060 vdd.n6453 vdd.n6452 0.151
R46061 vdd.n6452 vdd.n6451 0.151
R46062 vdd.n6451 vdd.n6450 0.151
R46063 vdd.n6659 vdd.n6648 0.151
R46064 vdd.n6648 vdd.n6647 0.151
R46065 vdd.n6647 vdd.n6646 0.151
R46066 vdd.n6646 vdd.n6645 0.151
R46067 vdd.n6645 vdd.n6644 0.151
R46068 vdd.n6644 vdd.n6643 0.151
R46069 vdd.n6643 vdd.n6642 0.151
R46070 vdd.n6642 vdd.n6641 0.151
R46071 vdd.n6641 vdd.n6640 0.151
R46072 vdd.n6640 vdd.n6639 0.151
R46073 vdd.n6639 vdd.n6638 0.151
R46074 vdd.n6638 vdd.n6637 0.151
R46075 vdd.n6637 vdd.n6636 0.151
R46076 vdd.n6636 vdd.n6635 0.151
R46077 vdd.n6635 vdd.n6634 0.151
R46078 vdd.n6634 vdd.n6633 0.151
R46079 vdd.n6633 vdd.n6632 0.151
R46080 vdd.n6632 vdd.n6631 0.151
R46081 vdd.n6631 vdd.n6630 0.151
R46082 vdd.n6839 vdd.n6828 0.151
R46083 vdd.n6828 vdd.n6827 0.151
R46084 vdd.n6827 vdd.n6826 0.151
R46085 vdd.n6826 vdd.n6825 0.151
R46086 vdd.n6825 vdd.n6824 0.151
R46087 vdd.n6824 vdd.n6823 0.151
R46088 vdd.n6823 vdd.n6822 0.151
R46089 vdd.n6822 vdd.n6821 0.151
R46090 vdd.n6821 vdd.n6820 0.151
R46091 vdd.n6820 vdd.n6819 0.151
R46092 vdd.n6819 vdd.n6818 0.151
R46093 vdd.n6818 vdd.n6817 0.151
R46094 vdd.n6817 vdd.n6816 0.151
R46095 vdd.n6816 vdd.n6815 0.151
R46096 vdd.n6815 vdd.n6814 0.151
R46097 vdd.n6814 vdd.n6813 0.151
R46098 vdd.n6813 vdd.n6812 0.151
R46099 vdd.n6812 vdd.n6811 0.151
R46100 vdd.n6811 vdd.n6810 0.151
R46101 vdd.n7019 vdd.n7008 0.151
R46102 vdd.n7008 vdd.n7007 0.151
R46103 vdd.n7007 vdd.n7006 0.151
R46104 vdd.n7006 vdd.n7005 0.151
R46105 vdd.n7005 vdd.n7004 0.151
R46106 vdd.n7004 vdd.n7003 0.151
R46107 vdd.n7003 vdd.n7002 0.151
R46108 vdd.n7002 vdd.n7001 0.151
R46109 vdd.n7001 vdd.n7000 0.151
R46110 vdd.n7000 vdd.n6999 0.151
R46111 vdd.n6999 vdd.n6998 0.151
R46112 vdd.n6998 vdd.n6997 0.151
R46113 vdd.n6997 vdd.n6996 0.151
R46114 vdd.n6996 vdd.n6995 0.151
R46115 vdd.n6995 vdd.n6994 0.151
R46116 vdd.n6994 vdd.n6993 0.151
R46117 vdd.n6993 vdd.n6992 0.151
R46118 vdd.n6992 vdd.n6991 0.151
R46119 vdd.n6991 vdd.n6990 0.151
R46120 vdd.n7199 vdd.n7188 0.151
R46121 vdd.n7188 vdd.n7187 0.151
R46122 vdd.n7187 vdd.n7186 0.151
R46123 vdd.n7186 vdd.n7185 0.151
R46124 vdd.n7185 vdd.n7184 0.151
R46125 vdd.n7184 vdd.n7183 0.151
R46126 vdd.n7183 vdd.n7182 0.151
R46127 vdd.n7182 vdd.n7181 0.151
R46128 vdd.n7181 vdd.n7180 0.151
R46129 vdd.n7180 vdd.n7179 0.151
R46130 vdd.n7179 vdd.n7178 0.151
R46131 vdd.n7178 vdd.n7177 0.151
R46132 vdd.n7177 vdd.n7176 0.151
R46133 vdd.n7176 vdd.n7175 0.151
R46134 vdd.n7175 vdd.n7174 0.151
R46135 vdd.n7174 vdd.n7173 0.151
R46136 vdd.n7173 vdd.n7172 0.151
R46137 vdd.n7172 vdd.n7171 0.151
R46138 vdd.n7171 vdd.n7170 0.151
R46139 vdd.n7379 vdd.n7368 0.151
R46140 vdd.n7368 vdd.n7367 0.151
R46141 vdd.n7367 vdd.n7366 0.151
R46142 vdd.n7366 vdd.n7365 0.151
R46143 vdd.n7365 vdd.n7364 0.151
R46144 vdd.n7364 vdd.n7363 0.151
R46145 vdd.n7363 vdd.n7362 0.151
R46146 vdd.n7362 vdd.n7361 0.151
R46147 vdd.n7361 vdd.n7360 0.151
R46148 vdd.n7360 vdd.n7359 0.151
R46149 vdd.n7359 vdd.n7358 0.151
R46150 vdd.n7358 vdd.n7357 0.151
R46151 vdd.n7357 vdd.n7356 0.151
R46152 vdd.n7356 vdd.n7355 0.151
R46153 vdd.n7355 vdd.n7354 0.151
R46154 vdd.n7354 vdd.n7353 0.151
R46155 vdd.n7353 vdd.n7352 0.151
R46156 vdd.n7352 vdd.n7351 0.151
R46157 vdd.n7351 vdd.n7350 0.151
R46158 vdd.n7559 vdd.n7548 0.151
R46159 vdd.n7548 vdd.n7547 0.151
R46160 vdd.n7547 vdd.n7546 0.151
R46161 vdd.n7546 vdd.n7545 0.151
R46162 vdd.n7545 vdd.n7544 0.151
R46163 vdd.n7544 vdd.n7543 0.151
R46164 vdd.n7543 vdd.n7542 0.151
R46165 vdd.n7542 vdd.n7541 0.151
R46166 vdd.n7541 vdd.n7540 0.151
R46167 vdd.n7540 vdd.n7539 0.151
R46168 vdd.n7539 vdd.n7538 0.151
R46169 vdd.n7538 vdd.n7537 0.151
R46170 vdd.n7537 vdd.n7536 0.151
R46171 vdd.n7536 vdd.n7535 0.151
R46172 vdd.n7535 vdd.n7534 0.151
R46173 vdd.n7534 vdd.n7533 0.151
R46174 vdd.n7533 vdd.n7532 0.151
R46175 vdd.n7532 vdd.n7531 0.151
R46176 vdd.n7531 vdd.n7530 0.151
R46177 vdd.n7739 vdd.n7728 0.151
R46178 vdd.n7728 vdd.n7727 0.151
R46179 vdd.n7727 vdd.n7726 0.151
R46180 vdd.n7726 vdd.n7725 0.151
R46181 vdd.n7725 vdd.n7724 0.151
R46182 vdd.n7724 vdd.n7723 0.151
R46183 vdd.n7723 vdd.n7722 0.151
R46184 vdd.n7722 vdd.n7721 0.151
R46185 vdd.n7721 vdd.n7720 0.151
R46186 vdd.n7720 vdd.n7719 0.151
R46187 vdd.n7719 vdd.n7718 0.151
R46188 vdd.n7718 vdd.n7717 0.151
R46189 vdd.n7717 vdd.n7716 0.151
R46190 vdd.n7716 vdd.n7715 0.151
R46191 vdd.n7715 vdd.n7714 0.151
R46192 vdd.n7714 vdd.n7713 0.151
R46193 vdd.n7713 vdd.n7712 0.151
R46194 vdd.n7712 vdd.n7711 0.151
R46195 vdd.n7711 vdd.n7710 0.151
R46196 vdd.n7919 vdd.n7908 0.151
R46197 vdd.n7908 vdd.n7907 0.151
R46198 vdd.n7907 vdd.n7906 0.151
R46199 vdd.n7906 vdd.n7905 0.151
R46200 vdd.n7905 vdd.n7904 0.151
R46201 vdd.n7904 vdd.n7903 0.151
R46202 vdd.n7903 vdd.n7902 0.151
R46203 vdd.n7902 vdd.n7901 0.151
R46204 vdd.n7901 vdd.n7900 0.151
R46205 vdd.n7900 vdd.n7899 0.151
R46206 vdd.n7899 vdd.n7898 0.151
R46207 vdd.n7898 vdd.n7897 0.151
R46208 vdd.n7897 vdd.n7896 0.151
R46209 vdd.n7896 vdd.n7895 0.151
R46210 vdd.n7895 vdd.n7894 0.151
R46211 vdd.n7894 vdd.n7893 0.151
R46212 vdd.n7893 vdd.n7892 0.151
R46213 vdd.n7892 vdd.n7891 0.151
R46214 vdd.n7891 vdd.n7890 0.151
R46215 vdd.n8099 vdd.n8088 0.151
R46216 vdd.n8088 vdd.n8087 0.151
R46217 vdd.n8087 vdd.n8086 0.151
R46218 vdd.n8086 vdd.n8085 0.151
R46219 vdd.n8085 vdd.n8084 0.151
R46220 vdd.n8084 vdd.n8083 0.151
R46221 vdd.n8083 vdd.n8082 0.151
R46222 vdd.n8082 vdd.n8081 0.151
R46223 vdd.n8081 vdd.n8080 0.151
R46224 vdd.n8080 vdd.n8079 0.151
R46225 vdd.n8079 vdd.n8078 0.151
R46226 vdd.n8078 vdd.n8077 0.151
R46227 vdd.n8077 vdd.n8076 0.151
R46228 vdd.n8076 vdd.n8075 0.151
R46229 vdd.n8075 vdd.n8074 0.151
R46230 vdd.n8074 vdd.n8073 0.151
R46231 vdd.n8073 vdd.n8072 0.151
R46232 vdd.n8072 vdd.n8071 0.151
R46233 vdd.n8071 vdd.n8070 0.151
R46234 vdd.n8279 vdd.n8268 0.151
R46235 vdd.n8268 vdd.n8267 0.151
R46236 vdd.n8267 vdd.n8266 0.151
R46237 vdd.n8266 vdd.n8265 0.151
R46238 vdd.n8265 vdd.n8264 0.151
R46239 vdd.n8264 vdd.n8263 0.151
R46240 vdd.n8263 vdd.n8262 0.151
R46241 vdd.n8262 vdd.n8261 0.151
R46242 vdd.n8261 vdd.n8260 0.151
R46243 vdd.n8260 vdd.n8259 0.151
R46244 vdd.n8259 vdd.n8258 0.151
R46245 vdd.n8258 vdd.n8257 0.151
R46246 vdd.n8257 vdd.n8256 0.151
R46247 vdd.n8256 vdd.n8255 0.151
R46248 vdd.n8255 vdd.n8254 0.151
R46249 vdd.n8254 vdd.n8253 0.151
R46250 vdd.n8253 vdd.n8252 0.151
R46251 vdd.n8252 vdd.n8251 0.151
R46252 vdd.n8251 vdd.n8250 0.151
R46253 vdd.n8459 vdd.n8448 0.151
R46254 vdd.n8448 vdd.n8447 0.151
R46255 vdd.n8447 vdd.n8446 0.151
R46256 vdd.n8446 vdd.n8445 0.151
R46257 vdd.n8445 vdd.n8444 0.151
R46258 vdd.n8444 vdd.n8443 0.151
R46259 vdd.n8443 vdd.n8442 0.151
R46260 vdd.n8442 vdd.n8441 0.151
R46261 vdd.n8441 vdd.n8440 0.151
R46262 vdd.n8440 vdd.n8439 0.151
R46263 vdd.n8439 vdd.n8438 0.151
R46264 vdd.n8438 vdd.n8437 0.151
R46265 vdd.n8437 vdd.n8436 0.151
R46266 vdd.n8436 vdd.n8435 0.151
R46267 vdd.n8435 vdd.n8434 0.151
R46268 vdd.n8434 vdd.n8433 0.151
R46269 vdd.n8433 vdd.n8432 0.151
R46270 vdd.n8432 vdd.n8431 0.151
R46271 vdd.n8431 vdd.n8430 0.151
R46272 vdd.n8639 vdd.n8628 0.151
R46273 vdd.n8628 vdd.n8627 0.151
R46274 vdd.n8627 vdd.n8626 0.151
R46275 vdd.n8626 vdd.n8625 0.151
R46276 vdd.n8625 vdd.n8624 0.151
R46277 vdd.n8624 vdd.n8623 0.151
R46278 vdd.n8623 vdd.n8622 0.151
R46279 vdd.n8622 vdd.n8621 0.151
R46280 vdd.n8621 vdd.n8620 0.151
R46281 vdd.n8620 vdd.n8619 0.151
R46282 vdd.n8619 vdd.n8618 0.151
R46283 vdd.n8618 vdd.n8617 0.151
R46284 vdd.n8617 vdd.n8616 0.151
R46285 vdd.n8616 vdd.n8615 0.151
R46286 vdd.n8615 vdd.n8614 0.151
R46287 vdd.n8614 vdd.n8613 0.151
R46288 vdd.n8613 vdd.n8612 0.151
R46289 vdd.n8612 vdd.n8611 0.151
R46290 vdd.n8611 vdd.n8610 0.151
R46291 vdd.n8819 vdd.n8808 0.151
R46292 vdd.n8808 vdd.n8807 0.151
R46293 vdd.n8807 vdd.n8806 0.151
R46294 vdd.n8806 vdd.n8805 0.151
R46295 vdd.n8805 vdd.n8804 0.151
R46296 vdd.n8804 vdd.n8803 0.151
R46297 vdd.n8803 vdd.n8802 0.151
R46298 vdd.n8802 vdd.n8801 0.151
R46299 vdd.n8801 vdd.n8800 0.151
R46300 vdd.n8800 vdd.n8799 0.151
R46301 vdd.n8799 vdd.n8798 0.151
R46302 vdd.n8798 vdd.n8797 0.151
R46303 vdd.n8797 vdd.n8796 0.151
R46304 vdd.n8796 vdd.n8795 0.151
R46305 vdd.n8795 vdd.n8794 0.151
R46306 vdd.n8794 vdd.n8793 0.151
R46307 vdd.n8793 vdd.n8792 0.151
R46308 vdd.n8792 vdd.n8791 0.151
R46309 vdd.n8791 vdd.n8790 0.151
R46310 vdd.n8999 vdd.n8988 0.151
R46311 vdd.n8988 vdd.n8987 0.151
R46312 vdd.n8987 vdd.n8986 0.151
R46313 vdd.n8986 vdd.n8985 0.151
R46314 vdd.n8985 vdd.n8984 0.151
R46315 vdd.n8984 vdd.n8983 0.151
R46316 vdd.n8983 vdd.n8982 0.151
R46317 vdd.n8982 vdd.n8981 0.151
R46318 vdd.n8981 vdd.n8980 0.151
R46319 vdd.n8980 vdd.n8979 0.151
R46320 vdd.n8979 vdd.n8978 0.151
R46321 vdd.n8978 vdd.n8977 0.151
R46322 vdd.n8977 vdd.n8976 0.151
R46323 vdd.n8976 vdd.n8975 0.151
R46324 vdd.n8975 vdd.n8974 0.151
R46325 vdd.n8974 vdd.n8973 0.151
R46326 vdd.n8973 vdd.n8972 0.151
R46327 vdd.n8972 vdd.n8971 0.151
R46328 vdd.n8971 vdd.n8970 0.151
R46329 vdd.n9179 vdd.n9168 0.151
R46330 vdd.n9168 vdd.n9167 0.151
R46331 vdd.n9167 vdd.n9166 0.151
R46332 vdd.n9166 vdd.n9165 0.151
R46333 vdd.n9165 vdd.n9164 0.151
R46334 vdd.n9164 vdd.n9163 0.151
R46335 vdd.n9163 vdd.n9162 0.151
R46336 vdd.n9162 vdd.n9161 0.151
R46337 vdd.n9161 vdd.n9160 0.151
R46338 vdd.n9160 vdd.n9159 0.151
R46339 vdd.n9159 vdd.n9158 0.151
R46340 vdd.n9158 vdd.n9157 0.151
R46341 vdd.n9157 vdd.n9156 0.151
R46342 vdd.n9156 vdd.n9155 0.151
R46343 vdd.n9155 vdd.n9154 0.151
R46344 vdd.n9154 vdd.n9153 0.151
R46345 vdd.n9153 vdd.n9152 0.151
R46346 vdd.n9152 vdd.n9151 0.151
R46347 vdd.n9151 vdd.n9150 0.151
R46348 vdd.n9359 vdd.n9348 0.151
R46349 vdd.n9348 vdd.n9347 0.151
R46350 vdd.n9347 vdd.n9346 0.151
R46351 vdd.n9346 vdd.n9345 0.151
R46352 vdd.n9345 vdd.n9344 0.151
R46353 vdd.n9344 vdd.n9343 0.151
R46354 vdd.n9343 vdd.n9342 0.151
R46355 vdd.n9342 vdd.n9341 0.151
R46356 vdd.n9341 vdd.n9340 0.151
R46357 vdd.n9340 vdd.n9339 0.151
R46358 vdd.n9339 vdd.n9338 0.151
R46359 vdd.n9338 vdd.n9337 0.151
R46360 vdd.n9337 vdd.n9336 0.151
R46361 vdd.n9336 vdd.n9335 0.151
R46362 vdd.n9335 vdd.n9334 0.151
R46363 vdd.n9334 vdd.n9333 0.151
R46364 vdd.n9333 vdd.n9332 0.151
R46365 vdd.n9332 vdd.n9331 0.151
R46366 vdd.n9331 vdd.n9330 0.151
R46367 vdd.n9539 vdd.n9528 0.151
R46368 vdd.n9528 vdd.n9527 0.151
R46369 vdd.n9527 vdd.n9526 0.151
R46370 vdd.n9526 vdd.n9525 0.151
R46371 vdd.n9525 vdd.n9524 0.151
R46372 vdd.n9524 vdd.n9523 0.151
R46373 vdd.n9523 vdd.n9522 0.151
R46374 vdd.n9522 vdd.n9521 0.151
R46375 vdd.n9521 vdd.n9520 0.151
R46376 vdd.n9520 vdd.n9519 0.151
R46377 vdd.n9519 vdd.n9518 0.151
R46378 vdd.n9518 vdd.n9517 0.151
R46379 vdd.n9517 vdd.n9516 0.151
R46380 vdd.n9516 vdd.n9515 0.151
R46381 vdd.n9515 vdd.n9514 0.151
R46382 vdd.n9514 vdd.n9513 0.151
R46383 vdd.n9513 vdd.n9512 0.151
R46384 vdd.n9512 vdd.n9511 0.151
R46385 vdd.n9511 vdd.n9510 0.151
R46386 vdd.n9719 vdd.n9708 0.151
R46387 vdd.n9708 vdd.n9707 0.151
R46388 vdd.n9707 vdd.n9706 0.151
R46389 vdd.n9706 vdd.n9705 0.151
R46390 vdd.n9705 vdd.n9704 0.151
R46391 vdd.n9704 vdd.n9703 0.151
R46392 vdd.n9703 vdd.n9702 0.151
R46393 vdd.n9702 vdd.n9701 0.151
R46394 vdd.n9701 vdd.n9700 0.151
R46395 vdd.n9700 vdd.n9699 0.151
R46396 vdd.n9699 vdd.n9698 0.151
R46397 vdd.n9698 vdd.n9697 0.151
R46398 vdd.n9697 vdd.n9696 0.151
R46399 vdd.n9696 vdd.n9695 0.151
R46400 vdd.n9695 vdd.n9694 0.151
R46401 vdd.n9694 vdd.n9693 0.151
R46402 vdd.n9693 vdd.n9692 0.151
R46403 vdd.n9692 vdd.n9691 0.151
R46404 vdd.n9691 vdd.n9690 0.151
R46405 vdd.n9899 vdd.n9888 0.151
R46406 vdd.n9888 vdd.n9887 0.151
R46407 vdd.n9887 vdd.n9886 0.151
R46408 vdd.n9886 vdd.n9885 0.151
R46409 vdd.n9885 vdd.n9884 0.151
R46410 vdd.n9884 vdd.n9883 0.151
R46411 vdd.n9883 vdd.n9882 0.151
R46412 vdd.n9882 vdd.n9881 0.151
R46413 vdd.n9881 vdd.n9880 0.151
R46414 vdd.n9880 vdd.n9879 0.151
R46415 vdd.n9879 vdd.n9878 0.151
R46416 vdd.n9878 vdd.n9877 0.151
R46417 vdd.n9877 vdd.n9876 0.151
R46418 vdd.n9876 vdd.n9875 0.151
R46419 vdd.n9875 vdd.n9874 0.151
R46420 vdd.n9874 vdd.n9873 0.151
R46421 vdd.n9873 vdd.n9872 0.151
R46422 vdd.n9872 vdd.n9871 0.151
R46423 vdd.n9871 vdd.n9870 0.151
R46424 vdd.n10079 vdd.n10068 0.151
R46425 vdd.n10068 vdd.n10067 0.151
R46426 vdd.n10067 vdd.n10066 0.151
R46427 vdd.n10066 vdd.n10065 0.151
R46428 vdd.n10065 vdd.n10064 0.151
R46429 vdd.n10064 vdd.n10063 0.151
R46430 vdd.n10063 vdd.n10062 0.151
R46431 vdd.n10062 vdd.n10061 0.151
R46432 vdd.n10061 vdd.n10060 0.151
R46433 vdd.n10060 vdd.n10059 0.151
R46434 vdd.n10059 vdd.n10058 0.151
R46435 vdd.n10058 vdd.n10057 0.151
R46436 vdd.n10057 vdd.n10056 0.151
R46437 vdd.n10056 vdd.n10055 0.151
R46438 vdd.n10055 vdd.n10054 0.151
R46439 vdd.n10054 vdd.n10053 0.151
R46440 vdd.n10053 vdd.n10052 0.151
R46441 vdd.n10052 vdd.n10051 0.151
R46442 vdd.n10051 vdd.n10050 0.151
R46443 vdd.n10259 vdd.n10248 0.151
R46444 vdd.n10248 vdd.n10247 0.151
R46445 vdd.n10247 vdd.n10246 0.151
R46446 vdd.n10246 vdd.n10245 0.151
R46447 vdd.n10245 vdd.n10244 0.151
R46448 vdd.n10244 vdd.n10243 0.151
R46449 vdd.n10243 vdd.n10242 0.151
R46450 vdd.n10242 vdd.n10241 0.151
R46451 vdd.n10241 vdd.n10240 0.151
R46452 vdd.n10240 vdd.n10239 0.151
R46453 vdd.n10239 vdd.n10238 0.151
R46454 vdd.n10238 vdd.n10237 0.151
R46455 vdd.n10237 vdd.n10236 0.151
R46456 vdd.n10236 vdd.n10235 0.151
R46457 vdd.n10235 vdd.n10234 0.151
R46458 vdd.n10234 vdd.n10233 0.151
R46459 vdd.n10233 vdd.n10232 0.151
R46460 vdd.n10232 vdd.n10231 0.151
R46461 vdd.n10231 vdd.n10230 0.151
R46462 vdd.n10439 vdd.n10428 0.151
R46463 vdd.n10428 vdd.n10427 0.151
R46464 vdd.n10427 vdd.n10426 0.151
R46465 vdd.n10426 vdd.n10425 0.151
R46466 vdd.n10425 vdd.n10424 0.151
R46467 vdd.n10424 vdd.n10423 0.151
R46468 vdd.n10423 vdd.n10422 0.151
R46469 vdd.n10422 vdd.n10421 0.151
R46470 vdd.n10421 vdd.n10420 0.151
R46471 vdd.n10420 vdd.n10419 0.151
R46472 vdd.n10419 vdd.n10418 0.151
R46473 vdd.n10418 vdd.n10417 0.151
R46474 vdd.n10417 vdd.n10416 0.151
R46475 vdd.n10416 vdd.n10415 0.151
R46476 vdd.n10415 vdd.n10414 0.151
R46477 vdd.n10414 vdd.n10413 0.151
R46478 vdd.n10413 vdd.n10412 0.151
R46479 vdd.n10412 vdd.n10411 0.151
R46480 vdd.n10411 vdd.n10410 0.151
R46481 vdd.n10619 vdd.n10608 0.151
R46482 vdd.n10608 vdd.n10607 0.151
R46483 vdd.n10607 vdd.n10606 0.151
R46484 vdd.n10606 vdd.n10605 0.151
R46485 vdd.n10605 vdd.n10604 0.151
R46486 vdd.n10604 vdd.n10603 0.151
R46487 vdd.n10603 vdd.n10602 0.151
R46488 vdd.n10602 vdd.n10601 0.151
R46489 vdd.n10601 vdd.n10600 0.151
R46490 vdd.n10600 vdd.n10599 0.151
R46491 vdd.n10599 vdd.n10598 0.151
R46492 vdd.n10598 vdd.n10597 0.151
R46493 vdd.n10597 vdd.n10596 0.151
R46494 vdd.n10596 vdd.n10595 0.151
R46495 vdd.n10595 vdd.n10594 0.151
R46496 vdd.n10594 vdd.n10593 0.151
R46497 vdd.n10593 vdd.n10592 0.151
R46498 vdd.n10592 vdd.n10591 0.151
R46499 vdd.n10591 vdd.n10590 0.151
R46500 vdd.n10799 vdd.n10788 0.151
R46501 vdd.n10788 vdd.n10787 0.151
R46502 vdd.n10787 vdd.n10786 0.151
R46503 vdd.n10786 vdd.n10785 0.151
R46504 vdd.n10785 vdd.n10784 0.151
R46505 vdd.n10784 vdd.n10783 0.151
R46506 vdd.n10783 vdd.n10782 0.151
R46507 vdd.n10782 vdd.n10781 0.151
R46508 vdd.n10781 vdd.n10780 0.151
R46509 vdd.n10780 vdd.n10779 0.151
R46510 vdd.n10779 vdd.n10778 0.151
R46511 vdd.n10778 vdd.n10777 0.151
R46512 vdd.n10777 vdd.n10776 0.151
R46513 vdd.n10776 vdd.n10775 0.151
R46514 vdd.n10775 vdd.n10774 0.151
R46515 vdd.n10774 vdd.n10773 0.151
R46516 vdd.n10773 vdd.n10772 0.151
R46517 vdd.n10772 vdd.n10771 0.151
R46518 vdd.n10771 vdd.n10770 0.151
R46519 vdd.n10979 vdd.n10968 0.151
R46520 vdd.n10968 vdd.n10967 0.151
R46521 vdd.n10967 vdd.n10966 0.151
R46522 vdd.n10966 vdd.n10965 0.151
R46523 vdd.n10965 vdd.n10964 0.151
R46524 vdd.n10964 vdd.n10963 0.151
R46525 vdd.n10963 vdd.n10962 0.151
R46526 vdd.n10962 vdd.n10961 0.151
R46527 vdd.n10961 vdd.n10960 0.151
R46528 vdd.n10960 vdd.n10959 0.151
R46529 vdd.n10959 vdd.n10958 0.151
R46530 vdd.n10958 vdd.n10957 0.151
R46531 vdd.n10957 vdd.n10956 0.151
R46532 vdd.n10956 vdd.n10955 0.151
R46533 vdd.n10955 vdd.n10954 0.151
R46534 vdd.n10954 vdd.n10953 0.151
R46535 vdd.n10953 vdd.n10952 0.151
R46536 vdd.n10952 vdd.n10951 0.151
R46537 vdd.n10951 vdd.n10950 0.151
R46538 vdd.n11159 vdd.n11148 0.151
R46539 vdd.n11148 vdd.n11147 0.151
R46540 vdd.n11147 vdd.n11146 0.151
R46541 vdd.n11146 vdd.n11145 0.151
R46542 vdd.n11145 vdd.n11144 0.151
R46543 vdd.n11144 vdd.n11143 0.151
R46544 vdd.n11143 vdd.n11142 0.151
R46545 vdd.n11142 vdd.n11141 0.151
R46546 vdd.n11141 vdd.n11140 0.151
R46547 vdd.n11140 vdd.n11139 0.151
R46548 vdd.n11139 vdd.n11138 0.151
R46549 vdd.n11138 vdd.n11137 0.151
R46550 vdd.n11137 vdd.n11136 0.151
R46551 vdd.n11136 vdd.n11135 0.151
R46552 vdd.n11135 vdd.n11134 0.151
R46553 vdd.n11134 vdd.n11133 0.151
R46554 vdd.n11133 vdd.n11132 0.151
R46555 vdd.n11132 vdd.n11131 0.151
R46556 vdd.n11131 vdd.n11130 0.151
R46557 vdd.n11339 vdd.n11328 0.151
R46558 vdd.n11328 vdd.n11327 0.151
R46559 vdd.n11327 vdd.n11326 0.151
R46560 vdd.n11326 vdd.n11325 0.151
R46561 vdd.n11325 vdd.n11324 0.151
R46562 vdd.n11324 vdd.n11323 0.151
R46563 vdd.n11323 vdd.n11322 0.151
R46564 vdd.n11322 vdd.n11321 0.151
R46565 vdd.n11321 vdd.n11320 0.151
R46566 vdd.n11320 vdd.n11319 0.151
R46567 vdd.n11319 vdd.n11318 0.151
R46568 vdd.n11318 vdd.n11317 0.151
R46569 vdd.n11317 vdd.n11316 0.151
R46570 vdd.n11316 vdd.n11315 0.151
R46571 vdd.n11315 vdd.n11314 0.151
R46572 vdd.n11314 vdd.n11313 0.151
R46573 vdd.n11313 vdd.n11312 0.151
R46574 vdd.n11312 vdd.n11311 0.151
R46575 vdd.n11311 vdd.n11310 0.151
R46576 vdd.n11362 vdd.n11360 0.131
R46577 vdd.n11365 vdd.n11363 0.131
R46578 vdd.n11368 vdd.n11366 0.131
R46579 vdd.n11371 vdd.n11369 0.131
R46580 vdd.n11374 vdd.n11372 0.131
R46581 vdd.n11377 vdd.n11375 0.131
R46582 vdd.n11380 vdd.n11378 0.131
R46583 vdd.n11383 vdd.n11381 0.131
R46584 vdd.n11386 vdd.n11384 0.131
R46585 vdd.n11390 vdd.n11388 0.131
R46586 vdd.n11393 vdd.n11391 0.131
R46587 vdd.n11396 vdd.n11394 0.131
R46588 vdd.n11399 vdd.n11397 0.131
R46589 vdd.n11402 vdd.n11400 0.131
R46590 vdd.n11405 vdd.n11403 0.131
R46591 vdd.n11408 vdd.n11406 0.131
R46592 vdd.n11411 vdd.n11409 0.131
R46593 vdd.n11413 vdd.n11411 0.131
R46594 vdd.n11415 vdd.n11413 0.131
R46595 vdd.n11409 vdd.n11408 0.131
R46596 vdd.n11406 vdd.n11405 0.131
R46597 vdd.n11403 vdd.n11402 0.131
R46598 vdd.n11400 vdd.n11399 0.131
R46599 vdd.n11397 vdd.n11396 0.131
R46600 vdd.n11394 vdd.n11393 0.131
R46601 vdd.n11391 vdd.n11390 0.131
R46602 vdd.n11388 vdd.n11387 0.131
R46603 vdd.n11384 vdd.n11383 0.131
R46604 vdd.n11381 vdd.n11380 0.131
R46605 vdd.n11378 vdd.n11377 0.131
R46606 vdd.n11375 vdd.n11374 0.131
R46607 vdd.n11372 vdd.n11371 0.131
R46608 vdd.n11369 vdd.n11368 0.131
R46609 vdd.n11366 vdd.n11365 0.131
R46610 vdd.n11363 vdd.n11362 0.131
R46611 vdd.n11360 vdd.n11359 0.131
R46612 vdd.n13484 vdd.n13482 0.131
R46613 vdd.n13487 vdd.n13485 0.131
R46614 vdd.n13490 vdd.n13488 0.131
R46615 vdd.n13493 vdd.n13491 0.131
R46616 vdd.n13496 vdd.n13494 0.131
R46617 vdd.n13499 vdd.n13497 0.131
R46618 vdd.n13502 vdd.n13500 0.131
R46619 vdd.n13505 vdd.n13503 0.131
R46620 vdd.n13509 vdd.n13507 0.131
R46621 vdd.n13512 vdd.n13510 0.131
R46622 vdd.n13515 vdd.n13513 0.131
R46623 vdd.n13518 vdd.n13516 0.131
R46624 vdd.n13521 vdd.n13519 0.131
R46625 vdd.n13524 vdd.n13522 0.131
R46626 vdd.n13527 vdd.n13525 0.131
R46627 vdd.n13530 vdd.n13528 0.131
R46628 vdd.n13532 vdd.n13530 0.131
R46629 vdd.n13479 vdd.n13478 0.131
R46630 vdd.n13534 vdd.n13532 0.131
R46631 vdd.n13528 vdd.n13527 0.131
R46632 vdd.n13525 vdd.n13524 0.131
R46633 vdd.n13522 vdd.n13521 0.131
R46634 vdd.n13519 vdd.n13518 0.131
R46635 vdd.n13516 vdd.n13515 0.131
R46636 vdd.n13513 vdd.n13512 0.131
R46637 vdd.n13510 vdd.n13509 0.131
R46638 vdd.n13507 vdd.n13506 0.131
R46639 vdd.n13503 vdd.n13502 0.131
R46640 vdd.n13500 vdd.n13499 0.131
R46641 vdd.n13497 vdd.n13496 0.131
R46642 vdd.n13494 vdd.n13493 0.131
R46643 vdd.n13491 vdd.n13490 0.131
R46644 vdd.n13488 vdd.n13487 0.131
R46645 vdd.n13485 vdd.n13484 0.131
R46646 vdd.n13482 vdd.n13481 0.131
R46647 vdd.n13481 vdd.n13479 0.131
R46648 vdd.n13535 vdd.n13458 0.123
R46649 vdd.n13536 vdd.n13278 0.123
R46650 vdd.n13537 vdd.n13098 0.123
R46651 vdd.n13538 vdd.n12918 0.123
R46652 vdd.n13539 vdd.n12738 0.123
R46653 vdd.n13540 vdd.n12558 0.123
R46654 vdd.n13541 vdd.n12378 0.123
R46655 vdd.n13542 vdd.n12198 0.123
R46656 vdd.n13543 vdd.n12018 0.123
R46657 vdd.n13544 vdd.n11838 0.123
R46658 vdd.n13545 vdd.n11658 0.123
R46659 vdd.n11478 vdd.n179 0.123
R46660 vdd.n11477 vdd.n359 0.123
R46661 vdd.n11476 vdd.n539 0.123
R46662 vdd.n11475 vdd.n719 0.123
R46663 vdd.n11474 vdd.n899 0.123
R46664 vdd.n11473 vdd.n1079 0.123
R46665 vdd.n11472 vdd.n1259 0.123
R46666 vdd.n11471 vdd.n1439 0.123
R46667 vdd.n11470 vdd.n1619 0.123
R46668 vdd.n11469 vdd.n1799 0.123
R46669 vdd.n11468 vdd.n1979 0.123
R46670 vdd.n11467 vdd.n2159 0.123
R46671 vdd.n11466 vdd.n2339 0.123
R46672 vdd.n11465 vdd.n2519 0.123
R46673 vdd.n11464 vdd.n2699 0.123
R46674 vdd.n11463 vdd.n2879 0.123
R46675 vdd.n11462 vdd.n3059 0.123
R46676 vdd.n11461 vdd.n3239 0.123
R46677 vdd.n11460 vdd.n3419 0.123
R46678 vdd.n11459 vdd.n3599 0.123
R46679 vdd.n11458 vdd.n3779 0.123
R46680 vdd.n11457 vdd.n3959 0.123
R46681 vdd.n11456 vdd.n4139 0.123
R46682 vdd.n11455 vdd.n4319 0.123
R46683 vdd.n11454 vdd.n4499 0.123
R46684 vdd.n11453 vdd.n4679 0.123
R46685 vdd.n11452 vdd.n4859 0.123
R46686 vdd.n11451 vdd.n5039 0.123
R46687 vdd.n11450 vdd.n5219 0.123
R46688 vdd.n11449 vdd.n5399 0.123
R46689 vdd.n11448 vdd.n5579 0.123
R46690 vdd.n11447 vdd.n5759 0.123
R46691 vdd.n11446 vdd.n5939 0.123
R46692 vdd.n11445 vdd.n6119 0.123
R46693 vdd.n11444 vdd.n6299 0.123
R46694 vdd.n11443 vdd.n6479 0.123
R46695 vdd.n11442 vdd.n6659 0.123
R46696 vdd.n11441 vdd.n6839 0.123
R46697 vdd.n11440 vdd.n7019 0.123
R46698 vdd.n11439 vdd.n7199 0.123
R46699 vdd.n11438 vdd.n7379 0.123
R46700 vdd.n11437 vdd.n7559 0.123
R46701 vdd.n11436 vdd.n7739 0.123
R46702 vdd.n11435 vdd.n7919 0.123
R46703 vdd.n11434 vdd.n8099 0.123
R46704 vdd.n11433 vdd.n8279 0.123
R46705 vdd.n11432 vdd.n8459 0.123
R46706 vdd.n11431 vdd.n8639 0.123
R46707 vdd.n11430 vdd.n8819 0.123
R46708 vdd.n11429 vdd.n8999 0.123
R46709 vdd.n11428 vdd.n9179 0.123
R46710 vdd.n11427 vdd.n9359 0.123
R46711 vdd.n11426 vdd.n9539 0.123
R46712 vdd.n11425 vdd.n9719 0.123
R46713 vdd.n11424 vdd.n9899 0.123
R46714 vdd.n11423 vdd.n10079 0.123
R46715 vdd.n11422 vdd.n10259 0.123
R46716 vdd.n11421 vdd.n10439 0.123
R46717 vdd.n11420 vdd.n10619 0.123
R46718 vdd.n11419 vdd.n10799 0.123
R46719 vdd.n11418 vdd.n10979 0.123
R46720 vdd.n11417 vdd.n11159 0.123
R46721 vdd.n11416 vdd.n11339 0.123
R46722 vdd.n13484 vdd.n13483 0.01
R46723 vdd.n13487 vdd.n13486 0.01
R46724 vdd.n13490 vdd.n13489 0.01
R46725 vdd.n13493 vdd.n13492 0.01
R46726 vdd.n13496 vdd.n13495 0.01
R46727 vdd.n13499 vdd.n13498 0.01
R46728 vdd.n13502 vdd.n13501 0.01
R46729 vdd.n13509 vdd.n13508 0.01
R46730 vdd.n13512 vdd.n13511 0.01
R46731 vdd.n13515 vdd.n13514 0.01
R46732 vdd.n13518 vdd.n13517 0.01
R46733 vdd.n13521 vdd.n13520 0.01
R46734 vdd.n13524 vdd.n13523 0.01
R46735 vdd.n13527 vdd.n13526 0.01
R46736 vdd.n13530 vdd.n13529 0.01
R46737 vdd.n13481 vdd.n13480 0.01
R46738 vdd.n13429 vdd.n13427 0.01
R46739 vdd.n13429 vdd.n13423 0.01
R46740 vdd.n13430 vdd.n13416 0.01
R46741 vdd.n13430 vdd.n13422 0.01
R46742 vdd.n13431 vdd.n13408 0.01
R46743 vdd.n13431 vdd.n13414 0.01
R46744 vdd.n13432 vdd.n13400 0.01
R46745 vdd.n13432 vdd.n13406 0.01
R46746 vdd.n13433 vdd.n13392 0.01
R46747 vdd.n13433 vdd.n13398 0.01
R46748 vdd.n13434 vdd.n13384 0.01
R46749 vdd.n13434 vdd.n13390 0.01
R46750 vdd.n13435 vdd.n13376 0.01
R46751 vdd.n13435 vdd.n13382 0.01
R46752 vdd.n13436 vdd.n13368 0.01
R46753 vdd.n13436 vdd.n13374 0.01
R46754 vdd.n13437 vdd.n13360 0.01
R46755 vdd.n13437 vdd.n13366 0.01
R46756 vdd.n13438 vdd.n13352 0.01
R46757 vdd.n13438 vdd.n13358 0.01
R46758 vdd.n13439 vdd.n13344 0.01
R46759 vdd.n13439 vdd.n13348 0.01
R46760 vdd.n13440 vdd.n13336 0.01
R46761 vdd.n13440 vdd.n13342 0.01
R46762 vdd.n13441 vdd.n13328 0.01
R46763 vdd.n13441 vdd.n13334 0.01
R46764 vdd.n13442 vdd.n13320 0.01
R46765 vdd.n13442 vdd.n13326 0.01
R46766 vdd.n13443 vdd.n13312 0.01
R46767 vdd.n13443 vdd.n13318 0.01
R46768 vdd.n13444 vdd.n13304 0.01
R46769 vdd.n13444 vdd.n13310 0.01
R46770 vdd.n13445 vdd.n13296 0.01
R46771 vdd.n13445 vdd.n13302 0.01
R46772 vdd.n13446 vdd.n13288 0.01
R46773 vdd.n13446 vdd.n13294 0.01
R46774 vdd.n13447 vdd.n13280 0.01
R46775 vdd.n13447 vdd.n13286 0.01
R46776 vdd.n13458 vdd.n13453 0.01
R46777 vdd.n13458 vdd.n13454 0.01
R46778 vdd.n13249 vdd.n13247 0.01
R46779 vdd.n13249 vdd.n13243 0.01
R46780 vdd.n13250 vdd.n13236 0.01
R46781 vdd.n13250 vdd.n13242 0.01
R46782 vdd.n13251 vdd.n13228 0.01
R46783 vdd.n13251 vdd.n13234 0.01
R46784 vdd.n13252 vdd.n13220 0.01
R46785 vdd.n13252 vdd.n13226 0.01
R46786 vdd.n13253 vdd.n13212 0.01
R46787 vdd.n13253 vdd.n13218 0.01
R46788 vdd.n13254 vdd.n13204 0.01
R46789 vdd.n13254 vdd.n13210 0.01
R46790 vdd.n13255 vdd.n13196 0.01
R46791 vdd.n13255 vdd.n13202 0.01
R46792 vdd.n13256 vdd.n13188 0.01
R46793 vdd.n13256 vdd.n13194 0.01
R46794 vdd.n13257 vdd.n13180 0.01
R46795 vdd.n13257 vdd.n13186 0.01
R46796 vdd.n13258 vdd.n13172 0.01
R46797 vdd.n13258 vdd.n13178 0.01
R46798 vdd.n13259 vdd.n13164 0.01
R46799 vdd.n13259 vdd.n13168 0.01
R46800 vdd.n13260 vdd.n13156 0.01
R46801 vdd.n13260 vdd.n13162 0.01
R46802 vdd.n13261 vdd.n13148 0.01
R46803 vdd.n13261 vdd.n13154 0.01
R46804 vdd.n13262 vdd.n13140 0.01
R46805 vdd.n13262 vdd.n13146 0.01
R46806 vdd.n13263 vdd.n13132 0.01
R46807 vdd.n13263 vdd.n13138 0.01
R46808 vdd.n13264 vdd.n13124 0.01
R46809 vdd.n13264 vdd.n13130 0.01
R46810 vdd.n13265 vdd.n13116 0.01
R46811 vdd.n13265 vdd.n13122 0.01
R46812 vdd.n13266 vdd.n13108 0.01
R46813 vdd.n13266 vdd.n13114 0.01
R46814 vdd.n13267 vdd.n13100 0.01
R46815 vdd.n13267 vdd.n13106 0.01
R46816 vdd.n13278 vdd.n13273 0.01
R46817 vdd.n13278 vdd.n13274 0.01
R46818 vdd.n13069 vdd.n13067 0.01
R46819 vdd.n13069 vdd.n13063 0.01
R46820 vdd.n13070 vdd.n13056 0.01
R46821 vdd.n13070 vdd.n13062 0.01
R46822 vdd.n13071 vdd.n13048 0.01
R46823 vdd.n13071 vdd.n13054 0.01
R46824 vdd.n13072 vdd.n13040 0.01
R46825 vdd.n13072 vdd.n13046 0.01
R46826 vdd.n13073 vdd.n13032 0.01
R46827 vdd.n13073 vdd.n13038 0.01
R46828 vdd.n13074 vdd.n13024 0.01
R46829 vdd.n13074 vdd.n13030 0.01
R46830 vdd.n13075 vdd.n13016 0.01
R46831 vdd.n13075 vdd.n13022 0.01
R46832 vdd.n13076 vdd.n13008 0.01
R46833 vdd.n13076 vdd.n13014 0.01
R46834 vdd.n13077 vdd.n13000 0.01
R46835 vdd.n13077 vdd.n13006 0.01
R46836 vdd.n13078 vdd.n12992 0.01
R46837 vdd.n13078 vdd.n12998 0.01
R46838 vdd.n13079 vdd.n12984 0.01
R46839 vdd.n13079 vdd.n12988 0.01
R46840 vdd.n13080 vdd.n12976 0.01
R46841 vdd.n13080 vdd.n12982 0.01
R46842 vdd.n13081 vdd.n12968 0.01
R46843 vdd.n13081 vdd.n12974 0.01
R46844 vdd.n13082 vdd.n12960 0.01
R46845 vdd.n13082 vdd.n12966 0.01
R46846 vdd.n13083 vdd.n12952 0.01
R46847 vdd.n13083 vdd.n12958 0.01
R46848 vdd.n13084 vdd.n12944 0.01
R46849 vdd.n13084 vdd.n12950 0.01
R46850 vdd.n13085 vdd.n12936 0.01
R46851 vdd.n13085 vdd.n12942 0.01
R46852 vdd.n13086 vdd.n12928 0.01
R46853 vdd.n13086 vdd.n12934 0.01
R46854 vdd.n13087 vdd.n12920 0.01
R46855 vdd.n13087 vdd.n12926 0.01
R46856 vdd.n13098 vdd.n13093 0.01
R46857 vdd.n13098 vdd.n13094 0.01
R46858 vdd.n12889 vdd.n12887 0.01
R46859 vdd.n12889 vdd.n12883 0.01
R46860 vdd.n12890 vdd.n12876 0.01
R46861 vdd.n12890 vdd.n12882 0.01
R46862 vdd.n12891 vdd.n12868 0.01
R46863 vdd.n12891 vdd.n12874 0.01
R46864 vdd.n12892 vdd.n12860 0.01
R46865 vdd.n12892 vdd.n12866 0.01
R46866 vdd.n12893 vdd.n12852 0.01
R46867 vdd.n12893 vdd.n12858 0.01
R46868 vdd.n12894 vdd.n12844 0.01
R46869 vdd.n12894 vdd.n12850 0.01
R46870 vdd.n12895 vdd.n12836 0.01
R46871 vdd.n12895 vdd.n12842 0.01
R46872 vdd.n12896 vdd.n12828 0.01
R46873 vdd.n12896 vdd.n12834 0.01
R46874 vdd.n12897 vdd.n12820 0.01
R46875 vdd.n12897 vdd.n12826 0.01
R46876 vdd.n12898 vdd.n12812 0.01
R46877 vdd.n12898 vdd.n12818 0.01
R46878 vdd.n12899 vdd.n12804 0.01
R46879 vdd.n12899 vdd.n12808 0.01
R46880 vdd.n12900 vdd.n12796 0.01
R46881 vdd.n12900 vdd.n12802 0.01
R46882 vdd.n12901 vdd.n12788 0.01
R46883 vdd.n12901 vdd.n12794 0.01
R46884 vdd.n12902 vdd.n12780 0.01
R46885 vdd.n12902 vdd.n12786 0.01
R46886 vdd.n12903 vdd.n12772 0.01
R46887 vdd.n12903 vdd.n12778 0.01
R46888 vdd.n12904 vdd.n12764 0.01
R46889 vdd.n12904 vdd.n12770 0.01
R46890 vdd.n12905 vdd.n12756 0.01
R46891 vdd.n12905 vdd.n12762 0.01
R46892 vdd.n12906 vdd.n12748 0.01
R46893 vdd.n12906 vdd.n12754 0.01
R46894 vdd.n12907 vdd.n12740 0.01
R46895 vdd.n12907 vdd.n12746 0.01
R46896 vdd.n12918 vdd.n12913 0.01
R46897 vdd.n12918 vdd.n12914 0.01
R46898 vdd.n12709 vdd.n12707 0.01
R46899 vdd.n12709 vdd.n12703 0.01
R46900 vdd.n12710 vdd.n12696 0.01
R46901 vdd.n12710 vdd.n12702 0.01
R46902 vdd.n12711 vdd.n12688 0.01
R46903 vdd.n12711 vdd.n12694 0.01
R46904 vdd.n12712 vdd.n12680 0.01
R46905 vdd.n12712 vdd.n12686 0.01
R46906 vdd.n12713 vdd.n12672 0.01
R46907 vdd.n12713 vdd.n12678 0.01
R46908 vdd.n12714 vdd.n12664 0.01
R46909 vdd.n12714 vdd.n12670 0.01
R46910 vdd.n12715 vdd.n12656 0.01
R46911 vdd.n12715 vdd.n12662 0.01
R46912 vdd.n12716 vdd.n12648 0.01
R46913 vdd.n12716 vdd.n12654 0.01
R46914 vdd.n12717 vdd.n12640 0.01
R46915 vdd.n12717 vdd.n12646 0.01
R46916 vdd.n12718 vdd.n12632 0.01
R46917 vdd.n12718 vdd.n12638 0.01
R46918 vdd.n12719 vdd.n12624 0.01
R46919 vdd.n12719 vdd.n12628 0.01
R46920 vdd.n12720 vdd.n12616 0.01
R46921 vdd.n12720 vdd.n12622 0.01
R46922 vdd.n12721 vdd.n12608 0.01
R46923 vdd.n12721 vdd.n12614 0.01
R46924 vdd.n12722 vdd.n12600 0.01
R46925 vdd.n12722 vdd.n12606 0.01
R46926 vdd.n12723 vdd.n12592 0.01
R46927 vdd.n12723 vdd.n12598 0.01
R46928 vdd.n12724 vdd.n12584 0.01
R46929 vdd.n12724 vdd.n12590 0.01
R46930 vdd.n12725 vdd.n12576 0.01
R46931 vdd.n12725 vdd.n12582 0.01
R46932 vdd.n12726 vdd.n12568 0.01
R46933 vdd.n12726 vdd.n12574 0.01
R46934 vdd.n12727 vdd.n12560 0.01
R46935 vdd.n12727 vdd.n12566 0.01
R46936 vdd.n12738 vdd.n12733 0.01
R46937 vdd.n12738 vdd.n12734 0.01
R46938 vdd.n12529 vdd.n12527 0.01
R46939 vdd.n12529 vdd.n12523 0.01
R46940 vdd.n12530 vdd.n12516 0.01
R46941 vdd.n12530 vdd.n12522 0.01
R46942 vdd.n12531 vdd.n12508 0.01
R46943 vdd.n12531 vdd.n12514 0.01
R46944 vdd.n12532 vdd.n12500 0.01
R46945 vdd.n12532 vdd.n12506 0.01
R46946 vdd.n12533 vdd.n12492 0.01
R46947 vdd.n12533 vdd.n12498 0.01
R46948 vdd.n12534 vdd.n12484 0.01
R46949 vdd.n12534 vdd.n12490 0.01
R46950 vdd.n12535 vdd.n12476 0.01
R46951 vdd.n12535 vdd.n12482 0.01
R46952 vdd.n12536 vdd.n12468 0.01
R46953 vdd.n12536 vdd.n12474 0.01
R46954 vdd.n12537 vdd.n12460 0.01
R46955 vdd.n12537 vdd.n12466 0.01
R46956 vdd.n12538 vdd.n12452 0.01
R46957 vdd.n12538 vdd.n12458 0.01
R46958 vdd.n12539 vdd.n12444 0.01
R46959 vdd.n12539 vdd.n12448 0.01
R46960 vdd.n12540 vdd.n12436 0.01
R46961 vdd.n12540 vdd.n12442 0.01
R46962 vdd.n12541 vdd.n12428 0.01
R46963 vdd.n12541 vdd.n12434 0.01
R46964 vdd.n12542 vdd.n12420 0.01
R46965 vdd.n12542 vdd.n12426 0.01
R46966 vdd.n12543 vdd.n12412 0.01
R46967 vdd.n12543 vdd.n12418 0.01
R46968 vdd.n12544 vdd.n12404 0.01
R46969 vdd.n12544 vdd.n12410 0.01
R46970 vdd.n12545 vdd.n12396 0.01
R46971 vdd.n12545 vdd.n12402 0.01
R46972 vdd.n12546 vdd.n12388 0.01
R46973 vdd.n12546 vdd.n12394 0.01
R46974 vdd.n12547 vdd.n12380 0.01
R46975 vdd.n12547 vdd.n12386 0.01
R46976 vdd.n12558 vdd.n12553 0.01
R46977 vdd.n12558 vdd.n12554 0.01
R46978 vdd.n12349 vdd.n12347 0.01
R46979 vdd.n12349 vdd.n12343 0.01
R46980 vdd.n12350 vdd.n12336 0.01
R46981 vdd.n12350 vdd.n12342 0.01
R46982 vdd.n12351 vdd.n12328 0.01
R46983 vdd.n12351 vdd.n12334 0.01
R46984 vdd.n12352 vdd.n12320 0.01
R46985 vdd.n12352 vdd.n12326 0.01
R46986 vdd.n12353 vdd.n12312 0.01
R46987 vdd.n12353 vdd.n12318 0.01
R46988 vdd.n12354 vdd.n12304 0.01
R46989 vdd.n12354 vdd.n12310 0.01
R46990 vdd.n12355 vdd.n12296 0.01
R46991 vdd.n12355 vdd.n12302 0.01
R46992 vdd.n12356 vdd.n12288 0.01
R46993 vdd.n12356 vdd.n12294 0.01
R46994 vdd.n12357 vdd.n12280 0.01
R46995 vdd.n12357 vdd.n12286 0.01
R46996 vdd.n12358 vdd.n12272 0.01
R46997 vdd.n12358 vdd.n12278 0.01
R46998 vdd.n12359 vdd.n12264 0.01
R46999 vdd.n12359 vdd.n12268 0.01
R47000 vdd.n12360 vdd.n12256 0.01
R47001 vdd.n12360 vdd.n12262 0.01
R47002 vdd.n12361 vdd.n12248 0.01
R47003 vdd.n12361 vdd.n12254 0.01
R47004 vdd.n12362 vdd.n12240 0.01
R47005 vdd.n12362 vdd.n12246 0.01
R47006 vdd.n12363 vdd.n12232 0.01
R47007 vdd.n12363 vdd.n12238 0.01
R47008 vdd.n12364 vdd.n12224 0.01
R47009 vdd.n12364 vdd.n12230 0.01
R47010 vdd.n12365 vdd.n12216 0.01
R47011 vdd.n12365 vdd.n12222 0.01
R47012 vdd.n12366 vdd.n12208 0.01
R47013 vdd.n12366 vdd.n12214 0.01
R47014 vdd.n12367 vdd.n12200 0.01
R47015 vdd.n12367 vdd.n12206 0.01
R47016 vdd.n12378 vdd.n12373 0.01
R47017 vdd.n12378 vdd.n12374 0.01
R47018 vdd.n12169 vdd.n12167 0.01
R47019 vdd.n12169 vdd.n12163 0.01
R47020 vdd.n12170 vdd.n12156 0.01
R47021 vdd.n12170 vdd.n12162 0.01
R47022 vdd.n12171 vdd.n12148 0.01
R47023 vdd.n12171 vdd.n12154 0.01
R47024 vdd.n12172 vdd.n12140 0.01
R47025 vdd.n12172 vdd.n12146 0.01
R47026 vdd.n12173 vdd.n12132 0.01
R47027 vdd.n12173 vdd.n12138 0.01
R47028 vdd.n12174 vdd.n12124 0.01
R47029 vdd.n12174 vdd.n12130 0.01
R47030 vdd.n12175 vdd.n12116 0.01
R47031 vdd.n12175 vdd.n12122 0.01
R47032 vdd.n12176 vdd.n12108 0.01
R47033 vdd.n12176 vdd.n12114 0.01
R47034 vdd.n12177 vdd.n12100 0.01
R47035 vdd.n12177 vdd.n12106 0.01
R47036 vdd.n12178 vdd.n12092 0.01
R47037 vdd.n12178 vdd.n12098 0.01
R47038 vdd.n12179 vdd.n12084 0.01
R47039 vdd.n12179 vdd.n12088 0.01
R47040 vdd.n12180 vdd.n12076 0.01
R47041 vdd.n12180 vdd.n12082 0.01
R47042 vdd.n12181 vdd.n12068 0.01
R47043 vdd.n12181 vdd.n12074 0.01
R47044 vdd.n12182 vdd.n12060 0.01
R47045 vdd.n12182 vdd.n12066 0.01
R47046 vdd.n12183 vdd.n12052 0.01
R47047 vdd.n12183 vdd.n12058 0.01
R47048 vdd.n12184 vdd.n12044 0.01
R47049 vdd.n12184 vdd.n12050 0.01
R47050 vdd.n12185 vdd.n12036 0.01
R47051 vdd.n12185 vdd.n12042 0.01
R47052 vdd.n12186 vdd.n12028 0.01
R47053 vdd.n12186 vdd.n12034 0.01
R47054 vdd.n12187 vdd.n12020 0.01
R47055 vdd.n12187 vdd.n12026 0.01
R47056 vdd.n12198 vdd.n12193 0.01
R47057 vdd.n12198 vdd.n12194 0.01
R47058 vdd.n11989 vdd.n11987 0.01
R47059 vdd.n11989 vdd.n11983 0.01
R47060 vdd.n11990 vdd.n11976 0.01
R47061 vdd.n11990 vdd.n11982 0.01
R47062 vdd.n11991 vdd.n11968 0.01
R47063 vdd.n11991 vdd.n11974 0.01
R47064 vdd.n11992 vdd.n11960 0.01
R47065 vdd.n11992 vdd.n11966 0.01
R47066 vdd.n11993 vdd.n11952 0.01
R47067 vdd.n11993 vdd.n11958 0.01
R47068 vdd.n11994 vdd.n11944 0.01
R47069 vdd.n11994 vdd.n11950 0.01
R47070 vdd.n11995 vdd.n11936 0.01
R47071 vdd.n11995 vdd.n11942 0.01
R47072 vdd.n11996 vdd.n11928 0.01
R47073 vdd.n11996 vdd.n11934 0.01
R47074 vdd.n11997 vdd.n11920 0.01
R47075 vdd.n11997 vdd.n11926 0.01
R47076 vdd.n11998 vdd.n11912 0.01
R47077 vdd.n11998 vdd.n11918 0.01
R47078 vdd.n11999 vdd.n11904 0.01
R47079 vdd.n11999 vdd.n11908 0.01
R47080 vdd.n12000 vdd.n11896 0.01
R47081 vdd.n12000 vdd.n11902 0.01
R47082 vdd.n12001 vdd.n11888 0.01
R47083 vdd.n12001 vdd.n11894 0.01
R47084 vdd.n12002 vdd.n11880 0.01
R47085 vdd.n12002 vdd.n11886 0.01
R47086 vdd.n12003 vdd.n11872 0.01
R47087 vdd.n12003 vdd.n11878 0.01
R47088 vdd.n12004 vdd.n11864 0.01
R47089 vdd.n12004 vdd.n11870 0.01
R47090 vdd.n12005 vdd.n11856 0.01
R47091 vdd.n12005 vdd.n11862 0.01
R47092 vdd.n12006 vdd.n11848 0.01
R47093 vdd.n12006 vdd.n11854 0.01
R47094 vdd.n12007 vdd.n11840 0.01
R47095 vdd.n12007 vdd.n11846 0.01
R47096 vdd.n12018 vdd.n12013 0.01
R47097 vdd.n12018 vdd.n12014 0.01
R47098 vdd.n11809 vdd.n11807 0.01
R47099 vdd.n11809 vdd.n11803 0.01
R47100 vdd.n11810 vdd.n11796 0.01
R47101 vdd.n11810 vdd.n11802 0.01
R47102 vdd.n11811 vdd.n11788 0.01
R47103 vdd.n11811 vdd.n11794 0.01
R47104 vdd.n11812 vdd.n11780 0.01
R47105 vdd.n11812 vdd.n11786 0.01
R47106 vdd.n11813 vdd.n11772 0.01
R47107 vdd.n11813 vdd.n11778 0.01
R47108 vdd.n11814 vdd.n11764 0.01
R47109 vdd.n11814 vdd.n11770 0.01
R47110 vdd.n11815 vdd.n11756 0.01
R47111 vdd.n11815 vdd.n11762 0.01
R47112 vdd.n11816 vdd.n11748 0.01
R47113 vdd.n11816 vdd.n11754 0.01
R47114 vdd.n11817 vdd.n11740 0.01
R47115 vdd.n11817 vdd.n11746 0.01
R47116 vdd.n11818 vdd.n11732 0.01
R47117 vdd.n11818 vdd.n11738 0.01
R47118 vdd.n11819 vdd.n11724 0.01
R47119 vdd.n11819 vdd.n11728 0.01
R47120 vdd.n11820 vdd.n11716 0.01
R47121 vdd.n11820 vdd.n11722 0.01
R47122 vdd.n11821 vdd.n11708 0.01
R47123 vdd.n11821 vdd.n11714 0.01
R47124 vdd.n11822 vdd.n11700 0.01
R47125 vdd.n11822 vdd.n11706 0.01
R47126 vdd.n11823 vdd.n11692 0.01
R47127 vdd.n11823 vdd.n11698 0.01
R47128 vdd.n11824 vdd.n11684 0.01
R47129 vdd.n11824 vdd.n11690 0.01
R47130 vdd.n11825 vdd.n11676 0.01
R47131 vdd.n11825 vdd.n11682 0.01
R47132 vdd.n11826 vdd.n11668 0.01
R47133 vdd.n11826 vdd.n11674 0.01
R47134 vdd.n11827 vdd.n11660 0.01
R47135 vdd.n11827 vdd.n11666 0.01
R47136 vdd.n11838 vdd.n11833 0.01
R47137 vdd.n11838 vdd.n11834 0.01
R47138 vdd.n11629 vdd.n11627 0.01
R47139 vdd.n11629 vdd.n11623 0.01
R47140 vdd.n11630 vdd.n11616 0.01
R47141 vdd.n11630 vdd.n11622 0.01
R47142 vdd.n11631 vdd.n11608 0.01
R47143 vdd.n11631 vdd.n11614 0.01
R47144 vdd.n11632 vdd.n11600 0.01
R47145 vdd.n11632 vdd.n11606 0.01
R47146 vdd.n11633 vdd.n11592 0.01
R47147 vdd.n11633 vdd.n11598 0.01
R47148 vdd.n11634 vdd.n11584 0.01
R47149 vdd.n11634 vdd.n11590 0.01
R47150 vdd.n11635 vdd.n11576 0.01
R47151 vdd.n11635 vdd.n11582 0.01
R47152 vdd.n11636 vdd.n11568 0.01
R47153 vdd.n11636 vdd.n11574 0.01
R47154 vdd.n11637 vdd.n11560 0.01
R47155 vdd.n11637 vdd.n11566 0.01
R47156 vdd.n11638 vdd.n11552 0.01
R47157 vdd.n11638 vdd.n11558 0.01
R47158 vdd.n11639 vdd.n11544 0.01
R47159 vdd.n11639 vdd.n11548 0.01
R47160 vdd.n11640 vdd.n11536 0.01
R47161 vdd.n11640 vdd.n11542 0.01
R47162 vdd.n11641 vdd.n11528 0.01
R47163 vdd.n11641 vdd.n11534 0.01
R47164 vdd.n11642 vdd.n11520 0.01
R47165 vdd.n11642 vdd.n11526 0.01
R47166 vdd.n11643 vdd.n11512 0.01
R47167 vdd.n11643 vdd.n11518 0.01
R47168 vdd.n11644 vdd.n11504 0.01
R47169 vdd.n11644 vdd.n11510 0.01
R47170 vdd.n11645 vdd.n11496 0.01
R47171 vdd.n11645 vdd.n11502 0.01
R47172 vdd.n11646 vdd.n11488 0.01
R47173 vdd.n11646 vdd.n11494 0.01
R47174 vdd.n11647 vdd.n11480 0.01
R47175 vdd.n11647 vdd.n11486 0.01
R47176 vdd.n11658 vdd.n11653 0.01
R47177 vdd.n11658 vdd.n11654 0.01
R47178 vdd.n150 vdd.n148 0.01
R47179 vdd.n150 vdd.n144 0.01
R47180 vdd.n151 vdd.n137 0.01
R47181 vdd.n151 vdd.n143 0.01
R47182 vdd.n152 vdd.n129 0.01
R47183 vdd.n152 vdd.n135 0.01
R47184 vdd.n153 vdd.n121 0.01
R47185 vdd.n153 vdd.n127 0.01
R47186 vdd.n154 vdd.n113 0.01
R47187 vdd.n154 vdd.n119 0.01
R47188 vdd.n155 vdd.n105 0.01
R47189 vdd.n155 vdd.n111 0.01
R47190 vdd.n156 vdd.n97 0.01
R47191 vdd.n156 vdd.n103 0.01
R47192 vdd.n157 vdd.n89 0.01
R47193 vdd.n157 vdd.n95 0.01
R47194 vdd.n158 vdd.n81 0.01
R47195 vdd.n158 vdd.n87 0.01
R47196 vdd.n159 vdd.n73 0.01
R47197 vdd.n159 vdd.n79 0.01
R47198 vdd.n160 vdd.n65 0.01
R47199 vdd.n160 vdd.n69 0.01
R47200 vdd.n161 vdd.n57 0.01
R47201 vdd.n161 vdd.n63 0.01
R47202 vdd.n162 vdd.n49 0.01
R47203 vdd.n162 vdd.n55 0.01
R47204 vdd.n163 vdd.n41 0.01
R47205 vdd.n163 vdd.n47 0.01
R47206 vdd.n164 vdd.n33 0.01
R47207 vdd.n164 vdd.n39 0.01
R47208 vdd.n165 vdd.n25 0.01
R47209 vdd.n165 vdd.n31 0.01
R47210 vdd.n166 vdd.n17 0.01
R47211 vdd.n166 vdd.n23 0.01
R47212 vdd.n167 vdd.n9 0.01
R47213 vdd.n167 vdd.n15 0.01
R47214 vdd.n168 vdd.n1 0.01
R47215 vdd.n168 vdd.n7 0.01
R47216 vdd.n179 vdd.n174 0.01
R47217 vdd.n179 vdd.n175 0.01
R47218 vdd.n330 vdd.n328 0.01
R47219 vdd.n330 vdd.n324 0.01
R47220 vdd.n331 vdd.n317 0.01
R47221 vdd.n331 vdd.n323 0.01
R47222 vdd.n332 vdd.n309 0.01
R47223 vdd.n332 vdd.n315 0.01
R47224 vdd.n333 vdd.n301 0.01
R47225 vdd.n333 vdd.n307 0.01
R47226 vdd.n334 vdd.n293 0.01
R47227 vdd.n334 vdd.n299 0.01
R47228 vdd.n335 vdd.n285 0.01
R47229 vdd.n335 vdd.n291 0.01
R47230 vdd.n336 vdd.n277 0.01
R47231 vdd.n336 vdd.n283 0.01
R47232 vdd.n337 vdd.n269 0.01
R47233 vdd.n337 vdd.n275 0.01
R47234 vdd.n338 vdd.n261 0.01
R47235 vdd.n338 vdd.n267 0.01
R47236 vdd.n339 vdd.n253 0.01
R47237 vdd.n339 vdd.n259 0.01
R47238 vdd.n340 vdd.n245 0.01
R47239 vdd.n340 vdd.n249 0.01
R47240 vdd.n341 vdd.n237 0.01
R47241 vdd.n341 vdd.n243 0.01
R47242 vdd.n342 vdd.n229 0.01
R47243 vdd.n342 vdd.n235 0.01
R47244 vdd.n343 vdd.n221 0.01
R47245 vdd.n343 vdd.n227 0.01
R47246 vdd.n344 vdd.n213 0.01
R47247 vdd.n344 vdd.n219 0.01
R47248 vdd.n345 vdd.n205 0.01
R47249 vdd.n345 vdd.n211 0.01
R47250 vdd.n346 vdd.n197 0.01
R47251 vdd.n346 vdd.n203 0.01
R47252 vdd.n347 vdd.n189 0.01
R47253 vdd.n347 vdd.n195 0.01
R47254 vdd.n348 vdd.n181 0.01
R47255 vdd.n348 vdd.n187 0.01
R47256 vdd.n359 vdd.n354 0.01
R47257 vdd.n359 vdd.n355 0.01
R47258 vdd.n510 vdd.n508 0.01
R47259 vdd.n510 vdd.n504 0.01
R47260 vdd.n511 vdd.n497 0.01
R47261 vdd.n511 vdd.n503 0.01
R47262 vdd.n512 vdd.n489 0.01
R47263 vdd.n512 vdd.n495 0.01
R47264 vdd.n513 vdd.n481 0.01
R47265 vdd.n513 vdd.n487 0.01
R47266 vdd.n514 vdd.n473 0.01
R47267 vdd.n514 vdd.n479 0.01
R47268 vdd.n515 vdd.n465 0.01
R47269 vdd.n515 vdd.n471 0.01
R47270 vdd.n516 vdd.n457 0.01
R47271 vdd.n516 vdd.n463 0.01
R47272 vdd.n517 vdd.n449 0.01
R47273 vdd.n517 vdd.n455 0.01
R47274 vdd.n518 vdd.n441 0.01
R47275 vdd.n518 vdd.n447 0.01
R47276 vdd.n519 vdd.n433 0.01
R47277 vdd.n519 vdd.n439 0.01
R47278 vdd.n520 vdd.n425 0.01
R47279 vdd.n520 vdd.n429 0.01
R47280 vdd.n521 vdd.n417 0.01
R47281 vdd.n521 vdd.n423 0.01
R47282 vdd.n522 vdd.n409 0.01
R47283 vdd.n522 vdd.n415 0.01
R47284 vdd.n523 vdd.n401 0.01
R47285 vdd.n523 vdd.n407 0.01
R47286 vdd.n524 vdd.n393 0.01
R47287 vdd.n524 vdd.n399 0.01
R47288 vdd.n525 vdd.n385 0.01
R47289 vdd.n525 vdd.n391 0.01
R47290 vdd.n526 vdd.n377 0.01
R47291 vdd.n526 vdd.n383 0.01
R47292 vdd.n527 vdd.n369 0.01
R47293 vdd.n527 vdd.n375 0.01
R47294 vdd.n528 vdd.n361 0.01
R47295 vdd.n528 vdd.n367 0.01
R47296 vdd.n539 vdd.n534 0.01
R47297 vdd.n539 vdd.n535 0.01
R47298 vdd.n690 vdd.n688 0.01
R47299 vdd.n690 vdd.n684 0.01
R47300 vdd.n691 vdd.n677 0.01
R47301 vdd.n691 vdd.n683 0.01
R47302 vdd.n692 vdd.n669 0.01
R47303 vdd.n692 vdd.n675 0.01
R47304 vdd.n693 vdd.n661 0.01
R47305 vdd.n693 vdd.n667 0.01
R47306 vdd.n694 vdd.n653 0.01
R47307 vdd.n694 vdd.n659 0.01
R47308 vdd.n695 vdd.n645 0.01
R47309 vdd.n695 vdd.n651 0.01
R47310 vdd.n696 vdd.n637 0.01
R47311 vdd.n696 vdd.n643 0.01
R47312 vdd.n697 vdd.n629 0.01
R47313 vdd.n697 vdd.n635 0.01
R47314 vdd.n698 vdd.n621 0.01
R47315 vdd.n698 vdd.n627 0.01
R47316 vdd.n699 vdd.n613 0.01
R47317 vdd.n699 vdd.n619 0.01
R47318 vdd.n700 vdd.n605 0.01
R47319 vdd.n700 vdd.n609 0.01
R47320 vdd.n701 vdd.n597 0.01
R47321 vdd.n701 vdd.n603 0.01
R47322 vdd.n702 vdd.n589 0.01
R47323 vdd.n702 vdd.n595 0.01
R47324 vdd.n703 vdd.n581 0.01
R47325 vdd.n703 vdd.n587 0.01
R47326 vdd.n704 vdd.n573 0.01
R47327 vdd.n704 vdd.n579 0.01
R47328 vdd.n705 vdd.n565 0.01
R47329 vdd.n705 vdd.n571 0.01
R47330 vdd.n706 vdd.n557 0.01
R47331 vdd.n706 vdd.n563 0.01
R47332 vdd.n707 vdd.n549 0.01
R47333 vdd.n707 vdd.n555 0.01
R47334 vdd.n708 vdd.n541 0.01
R47335 vdd.n708 vdd.n547 0.01
R47336 vdd.n719 vdd.n714 0.01
R47337 vdd.n719 vdd.n715 0.01
R47338 vdd.n870 vdd.n868 0.01
R47339 vdd.n870 vdd.n864 0.01
R47340 vdd.n871 vdd.n857 0.01
R47341 vdd.n871 vdd.n863 0.01
R47342 vdd.n872 vdd.n849 0.01
R47343 vdd.n872 vdd.n855 0.01
R47344 vdd.n873 vdd.n841 0.01
R47345 vdd.n873 vdd.n847 0.01
R47346 vdd.n874 vdd.n833 0.01
R47347 vdd.n874 vdd.n839 0.01
R47348 vdd.n875 vdd.n825 0.01
R47349 vdd.n875 vdd.n831 0.01
R47350 vdd.n876 vdd.n817 0.01
R47351 vdd.n876 vdd.n823 0.01
R47352 vdd.n877 vdd.n809 0.01
R47353 vdd.n877 vdd.n815 0.01
R47354 vdd.n878 vdd.n801 0.01
R47355 vdd.n878 vdd.n807 0.01
R47356 vdd.n879 vdd.n793 0.01
R47357 vdd.n879 vdd.n799 0.01
R47358 vdd.n880 vdd.n785 0.01
R47359 vdd.n880 vdd.n789 0.01
R47360 vdd.n881 vdd.n777 0.01
R47361 vdd.n881 vdd.n783 0.01
R47362 vdd.n882 vdd.n769 0.01
R47363 vdd.n882 vdd.n775 0.01
R47364 vdd.n883 vdd.n761 0.01
R47365 vdd.n883 vdd.n767 0.01
R47366 vdd.n884 vdd.n753 0.01
R47367 vdd.n884 vdd.n759 0.01
R47368 vdd.n885 vdd.n745 0.01
R47369 vdd.n885 vdd.n751 0.01
R47370 vdd.n886 vdd.n737 0.01
R47371 vdd.n886 vdd.n743 0.01
R47372 vdd.n887 vdd.n729 0.01
R47373 vdd.n887 vdd.n735 0.01
R47374 vdd.n888 vdd.n721 0.01
R47375 vdd.n888 vdd.n727 0.01
R47376 vdd.n899 vdd.n894 0.01
R47377 vdd.n899 vdd.n895 0.01
R47378 vdd.n1050 vdd.n1048 0.01
R47379 vdd.n1050 vdd.n1044 0.01
R47380 vdd.n1051 vdd.n1037 0.01
R47381 vdd.n1051 vdd.n1043 0.01
R47382 vdd.n1052 vdd.n1029 0.01
R47383 vdd.n1052 vdd.n1035 0.01
R47384 vdd.n1053 vdd.n1021 0.01
R47385 vdd.n1053 vdd.n1027 0.01
R47386 vdd.n1054 vdd.n1013 0.01
R47387 vdd.n1054 vdd.n1019 0.01
R47388 vdd.n1055 vdd.n1005 0.01
R47389 vdd.n1055 vdd.n1011 0.01
R47390 vdd.n1056 vdd.n997 0.01
R47391 vdd.n1056 vdd.n1003 0.01
R47392 vdd.n1057 vdd.n989 0.01
R47393 vdd.n1057 vdd.n995 0.01
R47394 vdd.n1058 vdd.n981 0.01
R47395 vdd.n1058 vdd.n987 0.01
R47396 vdd.n1059 vdd.n973 0.01
R47397 vdd.n1059 vdd.n979 0.01
R47398 vdd.n1060 vdd.n965 0.01
R47399 vdd.n1060 vdd.n969 0.01
R47400 vdd.n1061 vdd.n957 0.01
R47401 vdd.n1061 vdd.n963 0.01
R47402 vdd.n1062 vdd.n949 0.01
R47403 vdd.n1062 vdd.n955 0.01
R47404 vdd.n1063 vdd.n941 0.01
R47405 vdd.n1063 vdd.n947 0.01
R47406 vdd.n1064 vdd.n933 0.01
R47407 vdd.n1064 vdd.n939 0.01
R47408 vdd.n1065 vdd.n925 0.01
R47409 vdd.n1065 vdd.n931 0.01
R47410 vdd.n1066 vdd.n917 0.01
R47411 vdd.n1066 vdd.n923 0.01
R47412 vdd.n1067 vdd.n909 0.01
R47413 vdd.n1067 vdd.n915 0.01
R47414 vdd.n1068 vdd.n901 0.01
R47415 vdd.n1068 vdd.n907 0.01
R47416 vdd.n1079 vdd.n1074 0.01
R47417 vdd.n1079 vdd.n1075 0.01
R47418 vdd.n1230 vdd.n1228 0.01
R47419 vdd.n1230 vdd.n1224 0.01
R47420 vdd.n1231 vdd.n1217 0.01
R47421 vdd.n1231 vdd.n1223 0.01
R47422 vdd.n1232 vdd.n1209 0.01
R47423 vdd.n1232 vdd.n1215 0.01
R47424 vdd.n1233 vdd.n1201 0.01
R47425 vdd.n1233 vdd.n1207 0.01
R47426 vdd.n1234 vdd.n1193 0.01
R47427 vdd.n1234 vdd.n1199 0.01
R47428 vdd.n1235 vdd.n1185 0.01
R47429 vdd.n1235 vdd.n1191 0.01
R47430 vdd.n1236 vdd.n1177 0.01
R47431 vdd.n1236 vdd.n1183 0.01
R47432 vdd.n1237 vdd.n1169 0.01
R47433 vdd.n1237 vdd.n1175 0.01
R47434 vdd.n1238 vdd.n1161 0.01
R47435 vdd.n1238 vdd.n1167 0.01
R47436 vdd.n1239 vdd.n1153 0.01
R47437 vdd.n1239 vdd.n1159 0.01
R47438 vdd.n1240 vdd.n1145 0.01
R47439 vdd.n1240 vdd.n1149 0.01
R47440 vdd.n1241 vdd.n1137 0.01
R47441 vdd.n1241 vdd.n1143 0.01
R47442 vdd.n1242 vdd.n1129 0.01
R47443 vdd.n1242 vdd.n1135 0.01
R47444 vdd.n1243 vdd.n1121 0.01
R47445 vdd.n1243 vdd.n1127 0.01
R47446 vdd.n1244 vdd.n1113 0.01
R47447 vdd.n1244 vdd.n1119 0.01
R47448 vdd.n1245 vdd.n1105 0.01
R47449 vdd.n1245 vdd.n1111 0.01
R47450 vdd.n1246 vdd.n1097 0.01
R47451 vdd.n1246 vdd.n1103 0.01
R47452 vdd.n1247 vdd.n1089 0.01
R47453 vdd.n1247 vdd.n1095 0.01
R47454 vdd.n1248 vdd.n1081 0.01
R47455 vdd.n1248 vdd.n1087 0.01
R47456 vdd.n1259 vdd.n1254 0.01
R47457 vdd.n1259 vdd.n1255 0.01
R47458 vdd.n1410 vdd.n1408 0.01
R47459 vdd.n1410 vdd.n1404 0.01
R47460 vdd.n1411 vdd.n1397 0.01
R47461 vdd.n1411 vdd.n1403 0.01
R47462 vdd.n1412 vdd.n1389 0.01
R47463 vdd.n1412 vdd.n1395 0.01
R47464 vdd.n1413 vdd.n1381 0.01
R47465 vdd.n1413 vdd.n1387 0.01
R47466 vdd.n1414 vdd.n1373 0.01
R47467 vdd.n1414 vdd.n1379 0.01
R47468 vdd.n1415 vdd.n1365 0.01
R47469 vdd.n1415 vdd.n1371 0.01
R47470 vdd.n1416 vdd.n1357 0.01
R47471 vdd.n1416 vdd.n1363 0.01
R47472 vdd.n1417 vdd.n1349 0.01
R47473 vdd.n1417 vdd.n1355 0.01
R47474 vdd.n1418 vdd.n1341 0.01
R47475 vdd.n1418 vdd.n1347 0.01
R47476 vdd.n1419 vdd.n1333 0.01
R47477 vdd.n1419 vdd.n1339 0.01
R47478 vdd.n1420 vdd.n1325 0.01
R47479 vdd.n1420 vdd.n1329 0.01
R47480 vdd.n1421 vdd.n1317 0.01
R47481 vdd.n1421 vdd.n1323 0.01
R47482 vdd.n1422 vdd.n1309 0.01
R47483 vdd.n1422 vdd.n1315 0.01
R47484 vdd.n1423 vdd.n1301 0.01
R47485 vdd.n1423 vdd.n1307 0.01
R47486 vdd.n1424 vdd.n1293 0.01
R47487 vdd.n1424 vdd.n1299 0.01
R47488 vdd.n1425 vdd.n1285 0.01
R47489 vdd.n1425 vdd.n1291 0.01
R47490 vdd.n1426 vdd.n1277 0.01
R47491 vdd.n1426 vdd.n1283 0.01
R47492 vdd.n1427 vdd.n1269 0.01
R47493 vdd.n1427 vdd.n1275 0.01
R47494 vdd.n1428 vdd.n1261 0.01
R47495 vdd.n1428 vdd.n1267 0.01
R47496 vdd.n1439 vdd.n1434 0.01
R47497 vdd.n1439 vdd.n1435 0.01
R47498 vdd.n1590 vdd.n1588 0.01
R47499 vdd.n1590 vdd.n1584 0.01
R47500 vdd.n1591 vdd.n1577 0.01
R47501 vdd.n1591 vdd.n1583 0.01
R47502 vdd.n1592 vdd.n1569 0.01
R47503 vdd.n1592 vdd.n1575 0.01
R47504 vdd.n1593 vdd.n1561 0.01
R47505 vdd.n1593 vdd.n1567 0.01
R47506 vdd.n1594 vdd.n1553 0.01
R47507 vdd.n1594 vdd.n1559 0.01
R47508 vdd.n1595 vdd.n1545 0.01
R47509 vdd.n1595 vdd.n1551 0.01
R47510 vdd.n1596 vdd.n1537 0.01
R47511 vdd.n1596 vdd.n1543 0.01
R47512 vdd.n1597 vdd.n1529 0.01
R47513 vdd.n1597 vdd.n1535 0.01
R47514 vdd.n1598 vdd.n1521 0.01
R47515 vdd.n1598 vdd.n1527 0.01
R47516 vdd.n1599 vdd.n1513 0.01
R47517 vdd.n1599 vdd.n1519 0.01
R47518 vdd.n1600 vdd.n1505 0.01
R47519 vdd.n1600 vdd.n1509 0.01
R47520 vdd.n1601 vdd.n1497 0.01
R47521 vdd.n1601 vdd.n1503 0.01
R47522 vdd.n1602 vdd.n1489 0.01
R47523 vdd.n1602 vdd.n1495 0.01
R47524 vdd.n1603 vdd.n1481 0.01
R47525 vdd.n1603 vdd.n1487 0.01
R47526 vdd.n1604 vdd.n1473 0.01
R47527 vdd.n1604 vdd.n1479 0.01
R47528 vdd.n1605 vdd.n1465 0.01
R47529 vdd.n1605 vdd.n1471 0.01
R47530 vdd.n1606 vdd.n1457 0.01
R47531 vdd.n1606 vdd.n1463 0.01
R47532 vdd.n1607 vdd.n1449 0.01
R47533 vdd.n1607 vdd.n1455 0.01
R47534 vdd.n1608 vdd.n1441 0.01
R47535 vdd.n1608 vdd.n1447 0.01
R47536 vdd.n1619 vdd.n1614 0.01
R47537 vdd.n1619 vdd.n1615 0.01
R47538 vdd.n1770 vdd.n1768 0.01
R47539 vdd.n1770 vdd.n1764 0.01
R47540 vdd.n1771 vdd.n1757 0.01
R47541 vdd.n1771 vdd.n1763 0.01
R47542 vdd.n1772 vdd.n1749 0.01
R47543 vdd.n1772 vdd.n1755 0.01
R47544 vdd.n1773 vdd.n1741 0.01
R47545 vdd.n1773 vdd.n1747 0.01
R47546 vdd.n1774 vdd.n1733 0.01
R47547 vdd.n1774 vdd.n1739 0.01
R47548 vdd.n1775 vdd.n1725 0.01
R47549 vdd.n1775 vdd.n1731 0.01
R47550 vdd.n1776 vdd.n1717 0.01
R47551 vdd.n1776 vdd.n1723 0.01
R47552 vdd.n1777 vdd.n1709 0.01
R47553 vdd.n1777 vdd.n1715 0.01
R47554 vdd.n1778 vdd.n1701 0.01
R47555 vdd.n1778 vdd.n1707 0.01
R47556 vdd.n1779 vdd.n1693 0.01
R47557 vdd.n1779 vdd.n1699 0.01
R47558 vdd.n1780 vdd.n1685 0.01
R47559 vdd.n1780 vdd.n1689 0.01
R47560 vdd.n1781 vdd.n1677 0.01
R47561 vdd.n1781 vdd.n1683 0.01
R47562 vdd.n1782 vdd.n1669 0.01
R47563 vdd.n1782 vdd.n1675 0.01
R47564 vdd.n1783 vdd.n1661 0.01
R47565 vdd.n1783 vdd.n1667 0.01
R47566 vdd.n1784 vdd.n1653 0.01
R47567 vdd.n1784 vdd.n1659 0.01
R47568 vdd.n1785 vdd.n1645 0.01
R47569 vdd.n1785 vdd.n1651 0.01
R47570 vdd.n1786 vdd.n1637 0.01
R47571 vdd.n1786 vdd.n1643 0.01
R47572 vdd.n1787 vdd.n1629 0.01
R47573 vdd.n1787 vdd.n1635 0.01
R47574 vdd.n1788 vdd.n1621 0.01
R47575 vdd.n1788 vdd.n1627 0.01
R47576 vdd.n1799 vdd.n1794 0.01
R47577 vdd.n1799 vdd.n1795 0.01
R47578 vdd.n1950 vdd.n1948 0.01
R47579 vdd.n1950 vdd.n1944 0.01
R47580 vdd.n1951 vdd.n1937 0.01
R47581 vdd.n1951 vdd.n1943 0.01
R47582 vdd.n1952 vdd.n1929 0.01
R47583 vdd.n1952 vdd.n1935 0.01
R47584 vdd.n1953 vdd.n1921 0.01
R47585 vdd.n1953 vdd.n1927 0.01
R47586 vdd.n1954 vdd.n1913 0.01
R47587 vdd.n1954 vdd.n1919 0.01
R47588 vdd.n1955 vdd.n1905 0.01
R47589 vdd.n1955 vdd.n1911 0.01
R47590 vdd.n1956 vdd.n1897 0.01
R47591 vdd.n1956 vdd.n1903 0.01
R47592 vdd.n1957 vdd.n1889 0.01
R47593 vdd.n1957 vdd.n1895 0.01
R47594 vdd.n1958 vdd.n1881 0.01
R47595 vdd.n1958 vdd.n1887 0.01
R47596 vdd.n1959 vdd.n1873 0.01
R47597 vdd.n1959 vdd.n1879 0.01
R47598 vdd.n1960 vdd.n1865 0.01
R47599 vdd.n1960 vdd.n1869 0.01
R47600 vdd.n1961 vdd.n1857 0.01
R47601 vdd.n1961 vdd.n1863 0.01
R47602 vdd.n1962 vdd.n1849 0.01
R47603 vdd.n1962 vdd.n1855 0.01
R47604 vdd.n1963 vdd.n1841 0.01
R47605 vdd.n1963 vdd.n1847 0.01
R47606 vdd.n1964 vdd.n1833 0.01
R47607 vdd.n1964 vdd.n1839 0.01
R47608 vdd.n1965 vdd.n1825 0.01
R47609 vdd.n1965 vdd.n1831 0.01
R47610 vdd.n1966 vdd.n1817 0.01
R47611 vdd.n1966 vdd.n1823 0.01
R47612 vdd.n1967 vdd.n1809 0.01
R47613 vdd.n1967 vdd.n1815 0.01
R47614 vdd.n1968 vdd.n1801 0.01
R47615 vdd.n1968 vdd.n1807 0.01
R47616 vdd.n1979 vdd.n1974 0.01
R47617 vdd.n1979 vdd.n1975 0.01
R47618 vdd.n2130 vdd.n2128 0.01
R47619 vdd.n2130 vdd.n2124 0.01
R47620 vdd.n2131 vdd.n2117 0.01
R47621 vdd.n2131 vdd.n2123 0.01
R47622 vdd.n2132 vdd.n2109 0.01
R47623 vdd.n2132 vdd.n2115 0.01
R47624 vdd.n2133 vdd.n2101 0.01
R47625 vdd.n2133 vdd.n2107 0.01
R47626 vdd.n2134 vdd.n2093 0.01
R47627 vdd.n2134 vdd.n2099 0.01
R47628 vdd.n2135 vdd.n2085 0.01
R47629 vdd.n2135 vdd.n2091 0.01
R47630 vdd.n2136 vdd.n2077 0.01
R47631 vdd.n2136 vdd.n2083 0.01
R47632 vdd.n2137 vdd.n2069 0.01
R47633 vdd.n2137 vdd.n2075 0.01
R47634 vdd.n2138 vdd.n2061 0.01
R47635 vdd.n2138 vdd.n2067 0.01
R47636 vdd.n2139 vdd.n2053 0.01
R47637 vdd.n2139 vdd.n2059 0.01
R47638 vdd.n2140 vdd.n2045 0.01
R47639 vdd.n2140 vdd.n2049 0.01
R47640 vdd.n2141 vdd.n2037 0.01
R47641 vdd.n2141 vdd.n2043 0.01
R47642 vdd.n2142 vdd.n2029 0.01
R47643 vdd.n2142 vdd.n2035 0.01
R47644 vdd.n2143 vdd.n2021 0.01
R47645 vdd.n2143 vdd.n2027 0.01
R47646 vdd.n2144 vdd.n2013 0.01
R47647 vdd.n2144 vdd.n2019 0.01
R47648 vdd.n2145 vdd.n2005 0.01
R47649 vdd.n2145 vdd.n2011 0.01
R47650 vdd.n2146 vdd.n1997 0.01
R47651 vdd.n2146 vdd.n2003 0.01
R47652 vdd.n2147 vdd.n1989 0.01
R47653 vdd.n2147 vdd.n1995 0.01
R47654 vdd.n2148 vdd.n1981 0.01
R47655 vdd.n2148 vdd.n1987 0.01
R47656 vdd.n2159 vdd.n2154 0.01
R47657 vdd.n2159 vdd.n2155 0.01
R47658 vdd.n2310 vdd.n2308 0.01
R47659 vdd.n2310 vdd.n2304 0.01
R47660 vdd.n2311 vdd.n2297 0.01
R47661 vdd.n2311 vdd.n2303 0.01
R47662 vdd.n2312 vdd.n2289 0.01
R47663 vdd.n2312 vdd.n2295 0.01
R47664 vdd.n2313 vdd.n2281 0.01
R47665 vdd.n2313 vdd.n2287 0.01
R47666 vdd.n2314 vdd.n2273 0.01
R47667 vdd.n2314 vdd.n2279 0.01
R47668 vdd.n2315 vdd.n2265 0.01
R47669 vdd.n2315 vdd.n2271 0.01
R47670 vdd.n2316 vdd.n2257 0.01
R47671 vdd.n2316 vdd.n2263 0.01
R47672 vdd.n2317 vdd.n2249 0.01
R47673 vdd.n2317 vdd.n2255 0.01
R47674 vdd.n2318 vdd.n2241 0.01
R47675 vdd.n2318 vdd.n2247 0.01
R47676 vdd.n2319 vdd.n2233 0.01
R47677 vdd.n2319 vdd.n2239 0.01
R47678 vdd.n2320 vdd.n2225 0.01
R47679 vdd.n2320 vdd.n2229 0.01
R47680 vdd.n2321 vdd.n2217 0.01
R47681 vdd.n2321 vdd.n2223 0.01
R47682 vdd.n2322 vdd.n2209 0.01
R47683 vdd.n2322 vdd.n2215 0.01
R47684 vdd.n2323 vdd.n2201 0.01
R47685 vdd.n2323 vdd.n2207 0.01
R47686 vdd.n2324 vdd.n2193 0.01
R47687 vdd.n2324 vdd.n2199 0.01
R47688 vdd.n2325 vdd.n2185 0.01
R47689 vdd.n2325 vdd.n2191 0.01
R47690 vdd.n2326 vdd.n2177 0.01
R47691 vdd.n2326 vdd.n2183 0.01
R47692 vdd.n2327 vdd.n2169 0.01
R47693 vdd.n2327 vdd.n2175 0.01
R47694 vdd.n2328 vdd.n2161 0.01
R47695 vdd.n2328 vdd.n2167 0.01
R47696 vdd.n2339 vdd.n2334 0.01
R47697 vdd.n2339 vdd.n2335 0.01
R47698 vdd.n2490 vdd.n2488 0.01
R47699 vdd.n2490 vdd.n2484 0.01
R47700 vdd.n2491 vdd.n2477 0.01
R47701 vdd.n2491 vdd.n2483 0.01
R47702 vdd.n2492 vdd.n2469 0.01
R47703 vdd.n2492 vdd.n2475 0.01
R47704 vdd.n2493 vdd.n2461 0.01
R47705 vdd.n2493 vdd.n2467 0.01
R47706 vdd.n2494 vdd.n2453 0.01
R47707 vdd.n2494 vdd.n2459 0.01
R47708 vdd.n2495 vdd.n2445 0.01
R47709 vdd.n2495 vdd.n2451 0.01
R47710 vdd.n2496 vdd.n2437 0.01
R47711 vdd.n2496 vdd.n2443 0.01
R47712 vdd.n2497 vdd.n2429 0.01
R47713 vdd.n2497 vdd.n2435 0.01
R47714 vdd.n2498 vdd.n2421 0.01
R47715 vdd.n2498 vdd.n2427 0.01
R47716 vdd.n2499 vdd.n2413 0.01
R47717 vdd.n2499 vdd.n2419 0.01
R47718 vdd.n2500 vdd.n2405 0.01
R47719 vdd.n2500 vdd.n2409 0.01
R47720 vdd.n2501 vdd.n2397 0.01
R47721 vdd.n2501 vdd.n2403 0.01
R47722 vdd.n2502 vdd.n2389 0.01
R47723 vdd.n2502 vdd.n2395 0.01
R47724 vdd.n2503 vdd.n2381 0.01
R47725 vdd.n2503 vdd.n2387 0.01
R47726 vdd.n2504 vdd.n2373 0.01
R47727 vdd.n2504 vdd.n2379 0.01
R47728 vdd.n2505 vdd.n2365 0.01
R47729 vdd.n2505 vdd.n2371 0.01
R47730 vdd.n2506 vdd.n2357 0.01
R47731 vdd.n2506 vdd.n2363 0.01
R47732 vdd.n2507 vdd.n2349 0.01
R47733 vdd.n2507 vdd.n2355 0.01
R47734 vdd.n2508 vdd.n2341 0.01
R47735 vdd.n2508 vdd.n2347 0.01
R47736 vdd.n2519 vdd.n2514 0.01
R47737 vdd.n2519 vdd.n2515 0.01
R47738 vdd.n2670 vdd.n2668 0.01
R47739 vdd.n2670 vdd.n2664 0.01
R47740 vdd.n2671 vdd.n2657 0.01
R47741 vdd.n2671 vdd.n2663 0.01
R47742 vdd.n2672 vdd.n2649 0.01
R47743 vdd.n2672 vdd.n2655 0.01
R47744 vdd.n2673 vdd.n2641 0.01
R47745 vdd.n2673 vdd.n2647 0.01
R47746 vdd.n2674 vdd.n2633 0.01
R47747 vdd.n2674 vdd.n2639 0.01
R47748 vdd.n2675 vdd.n2625 0.01
R47749 vdd.n2675 vdd.n2631 0.01
R47750 vdd.n2676 vdd.n2617 0.01
R47751 vdd.n2676 vdd.n2623 0.01
R47752 vdd.n2677 vdd.n2609 0.01
R47753 vdd.n2677 vdd.n2615 0.01
R47754 vdd.n2678 vdd.n2601 0.01
R47755 vdd.n2678 vdd.n2607 0.01
R47756 vdd.n2679 vdd.n2593 0.01
R47757 vdd.n2679 vdd.n2599 0.01
R47758 vdd.n2680 vdd.n2585 0.01
R47759 vdd.n2680 vdd.n2589 0.01
R47760 vdd.n2681 vdd.n2577 0.01
R47761 vdd.n2681 vdd.n2583 0.01
R47762 vdd.n2682 vdd.n2569 0.01
R47763 vdd.n2682 vdd.n2575 0.01
R47764 vdd.n2683 vdd.n2561 0.01
R47765 vdd.n2683 vdd.n2567 0.01
R47766 vdd.n2684 vdd.n2553 0.01
R47767 vdd.n2684 vdd.n2559 0.01
R47768 vdd.n2685 vdd.n2545 0.01
R47769 vdd.n2685 vdd.n2551 0.01
R47770 vdd.n2686 vdd.n2537 0.01
R47771 vdd.n2686 vdd.n2543 0.01
R47772 vdd.n2687 vdd.n2529 0.01
R47773 vdd.n2687 vdd.n2535 0.01
R47774 vdd.n2688 vdd.n2521 0.01
R47775 vdd.n2688 vdd.n2527 0.01
R47776 vdd.n2699 vdd.n2694 0.01
R47777 vdd.n2699 vdd.n2695 0.01
R47778 vdd.n2850 vdd.n2848 0.01
R47779 vdd.n2850 vdd.n2844 0.01
R47780 vdd.n2851 vdd.n2837 0.01
R47781 vdd.n2851 vdd.n2843 0.01
R47782 vdd.n2852 vdd.n2829 0.01
R47783 vdd.n2852 vdd.n2835 0.01
R47784 vdd.n2853 vdd.n2821 0.01
R47785 vdd.n2853 vdd.n2827 0.01
R47786 vdd.n2854 vdd.n2813 0.01
R47787 vdd.n2854 vdd.n2819 0.01
R47788 vdd.n2855 vdd.n2805 0.01
R47789 vdd.n2855 vdd.n2811 0.01
R47790 vdd.n2856 vdd.n2797 0.01
R47791 vdd.n2856 vdd.n2803 0.01
R47792 vdd.n2857 vdd.n2789 0.01
R47793 vdd.n2857 vdd.n2795 0.01
R47794 vdd.n2858 vdd.n2781 0.01
R47795 vdd.n2858 vdd.n2787 0.01
R47796 vdd.n2859 vdd.n2773 0.01
R47797 vdd.n2859 vdd.n2779 0.01
R47798 vdd.n2860 vdd.n2765 0.01
R47799 vdd.n2860 vdd.n2769 0.01
R47800 vdd.n2861 vdd.n2757 0.01
R47801 vdd.n2861 vdd.n2763 0.01
R47802 vdd.n2862 vdd.n2749 0.01
R47803 vdd.n2862 vdd.n2755 0.01
R47804 vdd.n2863 vdd.n2741 0.01
R47805 vdd.n2863 vdd.n2747 0.01
R47806 vdd.n2864 vdd.n2733 0.01
R47807 vdd.n2864 vdd.n2739 0.01
R47808 vdd.n2865 vdd.n2725 0.01
R47809 vdd.n2865 vdd.n2731 0.01
R47810 vdd.n2866 vdd.n2717 0.01
R47811 vdd.n2866 vdd.n2723 0.01
R47812 vdd.n2867 vdd.n2709 0.01
R47813 vdd.n2867 vdd.n2715 0.01
R47814 vdd.n2868 vdd.n2701 0.01
R47815 vdd.n2868 vdd.n2707 0.01
R47816 vdd.n2879 vdd.n2874 0.01
R47817 vdd.n2879 vdd.n2875 0.01
R47818 vdd.n3030 vdd.n3028 0.01
R47819 vdd.n3030 vdd.n3024 0.01
R47820 vdd.n3031 vdd.n3017 0.01
R47821 vdd.n3031 vdd.n3023 0.01
R47822 vdd.n3032 vdd.n3009 0.01
R47823 vdd.n3032 vdd.n3015 0.01
R47824 vdd.n3033 vdd.n3001 0.01
R47825 vdd.n3033 vdd.n3007 0.01
R47826 vdd.n3034 vdd.n2993 0.01
R47827 vdd.n3034 vdd.n2999 0.01
R47828 vdd.n3035 vdd.n2985 0.01
R47829 vdd.n3035 vdd.n2991 0.01
R47830 vdd.n3036 vdd.n2977 0.01
R47831 vdd.n3036 vdd.n2983 0.01
R47832 vdd.n3037 vdd.n2969 0.01
R47833 vdd.n3037 vdd.n2975 0.01
R47834 vdd.n3038 vdd.n2961 0.01
R47835 vdd.n3038 vdd.n2967 0.01
R47836 vdd.n3039 vdd.n2953 0.01
R47837 vdd.n3039 vdd.n2959 0.01
R47838 vdd.n3040 vdd.n2945 0.01
R47839 vdd.n3040 vdd.n2949 0.01
R47840 vdd.n3041 vdd.n2937 0.01
R47841 vdd.n3041 vdd.n2943 0.01
R47842 vdd.n3042 vdd.n2929 0.01
R47843 vdd.n3042 vdd.n2935 0.01
R47844 vdd.n3043 vdd.n2921 0.01
R47845 vdd.n3043 vdd.n2927 0.01
R47846 vdd.n3044 vdd.n2913 0.01
R47847 vdd.n3044 vdd.n2919 0.01
R47848 vdd.n3045 vdd.n2905 0.01
R47849 vdd.n3045 vdd.n2911 0.01
R47850 vdd.n3046 vdd.n2897 0.01
R47851 vdd.n3046 vdd.n2903 0.01
R47852 vdd.n3047 vdd.n2889 0.01
R47853 vdd.n3047 vdd.n2895 0.01
R47854 vdd.n3048 vdd.n2881 0.01
R47855 vdd.n3048 vdd.n2887 0.01
R47856 vdd.n3059 vdd.n3054 0.01
R47857 vdd.n3059 vdd.n3055 0.01
R47858 vdd.n3210 vdd.n3208 0.01
R47859 vdd.n3210 vdd.n3204 0.01
R47860 vdd.n3211 vdd.n3197 0.01
R47861 vdd.n3211 vdd.n3203 0.01
R47862 vdd.n3212 vdd.n3189 0.01
R47863 vdd.n3212 vdd.n3195 0.01
R47864 vdd.n3213 vdd.n3181 0.01
R47865 vdd.n3213 vdd.n3187 0.01
R47866 vdd.n3214 vdd.n3173 0.01
R47867 vdd.n3214 vdd.n3179 0.01
R47868 vdd.n3215 vdd.n3165 0.01
R47869 vdd.n3215 vdd.n3171 0.01
R47870 vdd.n3216 vdd.n3157 0.01
R47871 vdd.n3216 vdd.n3163 0.01
R47872 vdd.n3217 vdd.n3149 0.01
R47873 vdd.n3217 vdd.n3155 0.01
R47874 vdd.n3218 vdd.n3141 0.01
R47875 vdd.n3218 vdd.n3147 0.01
R47876 vdd.n3219 vdd.n3133 0.01
R47877 vdd.n3219 vdd.n3139 0.01
R47878 vdd.n3220 vdd.n3125 0.01
R47879 vdd.n3220 vdd.n3129 0.01
R47880 vdd.n3221 vdd.n3117 0.01
R47881 vdd.n3221 vdd.n3123 0.01
R47882 vdd.n3222 vdd.n3109 0.01
R47883 vdd.n3222 vdd.n3115 0.01
R47884 vdd.n3223 vdd.n3101 0.01
R47885 vdd.n3223 vdd.n3107 0.01
R47886 vdd.n3224 vdd.n3093 0.01
R47887 vdd.n3224 vdd.n3099 0.01
R47888 vdd.n3225 vdd.n3085 0.01
R47889 vdd.n3225 vdd.n3091 0.01
R47890 vdd.n3226 vdd.n3077 0.01
R47891 vdd.n3226 vdd.n3083 0.01
R47892 vdd.n3227 vdd.n3069 0.01
R47893 vdd.n3227 vdd.n3075 0.01
R47894 vdd.n3228 vdd.n3061 0.01
R47895 vdd.n3228 vdd.n3067 0.01
R47896 vdd.n3239 vdd.n3234 0.01
R47897 vdd.n3239 vdd.n3235 0.01
R47898 vdd.n3390 vdd.n3388 0.01
R47899 vdd.n3390 vdd.n3384 0.01
R47900 vdd.n3391 vdd.n3377 0.01
R47901 vdd.n3391 vdd.n3383 0.01
R47902 vdd.n3392 vdd.n3369 0.01
R47903 vdd.n3392 vdd.n3375 0.01
R47904 vdd.n3393 vdd.n3361 0.01
R47905 vdd.n3393 vdd.n3367 0.01
R47906 vdd.n3394 vdd.n3353 0.01
R47907 vdd.n3394 vdd.n3359 0.01
R47908 vdd.n3395 vdd.n3345 0.01
R47909 vdd.n3395 vdd.n3351 0.01
R47910 vdd.n3396 vdd.n3337 0.01
R47911 vdd.n3396 vdd.n3343 0.01
R47912 vdd.n3397 vdd.n3329 0.01
R47913 vdd.n3397 vdd.n3335 0.01
R47914 vdd.n3398 vdd.n3321 0.01
R47915 vdd.n3398 vdd.n3327 0.01
R47916 vdd.n3399 vdd.n3313 0.01
R47917 vdd.n3399 vdd.n3319 0.01
R47918 vdd.n3400 vdd.n3305 0.01
R47919 vdd.n3400 vdd.n3309 0.01
R47920 vdd.n3401 vdd.n3297 0.01
R47921 vdd.n3401 vdd.n3303 0.01
R47922 vdd.n3402 vdd.n3289 0.01
R47923 vdd.n3402 vdd.n3295 0.01
R47924 vdd.n3403 vdd.n3281 0.01
R47925 vdd.n3403 vdd.n3287 0.01
R47926 vdd.n3404 vdd.n3273 0.01
R47927 vdd.n3404 vdd.n3279 0.01
R47928 vdd.n3405 vdd.n3265 0.01
R47929 vdd.n3405 vdd.n3271 0.01
R47930 vdd.n3406 vdd.n3257 0.01
R47931 vdd.n3406 vdd.n3263 0.01
R47932 vdd.n3407 vdd.n3249 0.01
R47933 vdd.n3407 vdd.n3255 0.01
R47934 vdd.n3408 vdd.n3241 0.01
R47935 vdd.n3408 vdd.n3247 0.01
R47936 vdd.n3419 vdd.n3414 0.01
R47937 vdd.n3419 vdd.n3415 0.01
R47938 vdd.n3570 vdd.n3568 0.01
R47939 vdd.n3570 vdd.n3564 0.01
R47940 vdd.n3571 vdd.n3557 0.01
R47941 vdd.n3571 vdd.n3563 0.01
R47942 vdd.n3572 vdd.n3549 0.01
R47943 vdd.n3572 vdd.n3555 0.01
R47944 vdd.n3573 vdd.n3541 0.01
R47945 vdd.n3573 vdd.n3547 0.01
R47946 vdd.n3574 vdd.n3533 0.01
R47947 vdd.n3574 vdd.n3539 0.01
R47948 vdd.n3575 vdd.n3525 0.01
R47949 vdd.n3575 vdd.n3531 0.01
R47950 vdd.n3576 vdd.n3517 0.01
R47951 vdd.n3576 vdd.n3523 0.01
R47952 vdd.n3577 vdd.n3509 0.01
R47953 vdd.n3577 vdd.n3515 0.01
R47954 vdd.n3578 vdd.n3501 0.01
R47955 vdd.n3578 vdd.n3507 0.01
R47956 vdd.n3579 vdd.n3493 0.01
R47957 vdd.n3579 vdd.n3499 0.01
R47958 vdd.n3580 vdd.n3485 0.01
R47959 vdd.n3580 vdd.n3489 0.01
R47960 vdd.n3581 vdd.n3477 0.01
R47961 vdd.n3581 vdd.n3483 0.01
R47962 vdd.n3582 vdd.n3469 0.01
R47963 vdd.n3582 vdd.n3475 0.01
R47964 vdd.n3583 vdd.n3461 0.01
R47965 vdd.n3583 vdd.n3467 0.01
R47966 vdd.n3584 vdd.n3453 0.01
R47967 vdd.n3584 vdd.n3459 0.01
R47968 vdd.n3585 vdd.n3445 0.01
R47969 vdd.n3585 vdd.n3451 0.01
R47970 vdd.n3586 vdd.n3437 0.01
R47971 vdd.n3586 vdd.n3443 0.01
R47972 vdd.n3587 vdd.n3429 0.01
R47973 vdd.n3587 vdd.n3435 0.01
R47974 vdd.n3588 vdd.n3421 0.01
R47975 vdd.n3588 vdd.n3427 0.01
R47976 vdd.n3599 vdd.n3594 0.01
R47977 vdd.n3599 vdd.n3595 0.01
R47978 vdd.n3750 vdd.n3748 0.01
R47979 vdd.n3750 vdd.n3744 0.01
R47980 vdd.n3751 vdd.n3737 0.01
R47981 vdd.n3751 vdd.n3743 0.01
R47982 vdd.n3752 vdd.n3729 0.01
R47983 vdd.n3752 vdd.n3735 0.01
R47984 vdd.n3753 vdd.n3721 0.01
R47985 vdd.n3753 vdd.n3727 0.01
R47986 vdd.n3754 vdd.n3713 0.01
R47987 vdd.n3754 vdd.n3719 0.01
R47988 vdd.n3755 vdd.n3705 0.01
R47989 vdd.n3755 vdd.n3711 0.01
R47990 vdd.n3756 vdd.n3697 0.01
R47991 vdd.n3756 vdd.n3703 0.01
R47992 vdd.n3757 vdd.n3689 0.01
R47993 vdd.n3757 vdd.n3695 0.01
R47994 vdd.n3758 vdd.n3681 0.01
R47995 vdd.n3758 vdd.n3687 0.01
R47996 vdd.n3759 vdd.n3673 0.01
R47997 vdd.n3759 vdd.n3679 0.01
R47998 vdd.n3760 vdd.n3665 0.01
R47999 vdd.n3760 vdd.n3669 0.01
R48000 vdd.n3761 vdd.n3657 0.01
R48001 vdd.n3761 vdd.n3663 0.01
R48002 vdd.n3762 vdd.n3649 0.01
R48003 vdd.n3762 vdd.n3655 0.01
R48004 vdd.n3763 vdd.n3641 0.01
R48005 vdd.n3763 vdd.n3647 0.01
R48006 vdd.n3764 vdd.n3633 0.01
R48007 vdd.n3764 vdd.n3639 0.01
R48008 vdd.n3765 vdd.n3625 0.01
R48009 vdd.n3765 vdd.n3631 0.01
R48010 vdd.n3766 vdd.n3617 0.01
R48011 vdd.n3766 vdd.n3623 0.01
R48012 vdd.n3767 vdd.n3609 0.01
R48013 vdd.n3767 vdd.n3615 0.01
R48014 vdd.n3768 vdd.n3601 0.01
R48015 vdd.n3768 vdd.n3607 0.01
R48016 vdd.n3779 vdd.n3774 0.01
R48017 vdd.n3779 vdd.n3775 0.01
R48018 vdd.n3930 vdd.n3928 0.01
R48019 vdd.n3930 vdd.n3924 0.01
R48020 vdd.n3931 vdd.n3917 0.01
R48021 vdd.n3931 vdd.n3923 0.01
R48022 vdd.n3932 vdd.n3909 0.01
R48023 vdd.n3932 vdd.n3915 0.01
R48024 vdd.n3933 vdd.n3901 0.01
R48025 vdd.n3933 vdd.n3907 0.01
R48026 vdd.n3934 vdd.n3893 0.01
R48027 vdd.n3934 vdd.n3899 0.01
R48028 vdd.n3935 vdd.n3885 0.01
R48029 vdd.n3935 vdd.n3891 0.01
R48030 vdd.n3936 vdd.n3877 0.01
R48031 vdd.n3936 vdd.n3883 0.01
R48032 vdd.n3937 vdd.n3869 0.01
R48033 vdd.n3937 vdd.n3875 0.01
R48034 vdd.n3938 vdd.n3861 0.01
R48035 vdd.n3938 vdd.n3867 0.01
R48036 vdd.n3939 vdd.n3853 0.01
R48037 vdd.n3939 vdd.n3859 0.01
R48038 vdd.n3940 vdd.n3845 0.01
R48039 vdd.n3940 vdd.n3849 0.01
R48040 vdd.n3941 vdd.n3837 0.01
R48041 vdd.n3941 vdd.n3843 0.01
R48042 vdd.n3942 vdd.n3829 0.01
R48043 vdd.n3942 vdd.n3835 0.01
R48044 vdd.n3943 vdd.n3821 0.01
R48045 vdd.n3943 vdd.n3827 0.01
R48046 vdd.n3944 vdd.n3813 0.01
R48047 vdd.n3944 vdd.n3819 0.01
R48048 vdd.n3945 vdd.n3805 0.01
R48049 vdd.n3945 vdd.n3811 0.01
R48050 vdd.n3946 vdd.n3797 0.01
R48051 vdd.n3946 vdd.n3803 0.01
R48052 vdd.n3947 vdd.n3789 0.01
R48053 vdd.n3947 vdd.n3795 0.01
R48054 vdd.n3948 vdd.n3781 0.01
R48055 vdd.n3948 vdd.n3787 0.01
R48056 vdd.n3959 vdd.n3954 0.01
R48057 vdd.n3959 vdd.n3955 0.01
R48058 vdd.n4110 vdd.n4108 0.01
R48059 vdd.n4110 vdd.n4104 0.01
R48060 vdd.n4111 vdd.n4097 0.01
R48061 vdd.n4111 vdd.n4103 0.01
R48062 vdd.n4112 vdd.n4089 0.01
R48063 vdd.n4112 vdd.n4095 0.01
R48064 vdd.n4113 vdd.n4081 0.01
R48065 vdd.n4113 vdd.n4087 0.01
R48066 vdd.n4114 vdd.n4073 0.01
R48067 vdd.n4114 vdd.n4079 0.01
R48068 vdd.n4115 vdd.n4065 0.01
R48069 vdd.n4115 vdd.n4071 0.01
R48070 vdd.n4116 vdd.n4057 0.01
R48071 vdd.n4116 vdd.n4063 0.01
R48072 vdd.n4117 vdd.n4049 0.01
R48073 vdd.n4117 vdd.n4055 0.01
R48074 vdd.n4118 vdd.n4041 0.01
R48075 vdd.n4118 vdd.n4047 0.01
R48076 vdd.n4119 vdd.n4033 0.01
R48077 vdd.n4119 vdd.n4039 0.01
R48078 vdd.n4120 vdd.n4025 0.01
R48079 vdd.n4120 vdd.n4029 0.01
R48080 vdd.n4121 vdd.n4017 0.01
R48081 vdd.n4121 vdd.n4023 0.01
R48082 vdd.n4122 vdd.n4009 0.01
R48083 vdd.n4122 vdd.n4015 0.01
R48084 vdd.n4123 vdd.n4001 0.01
R48085 vdd.n4123 vdd.n4007 0.01
R48086 vdd.n4124 vdd.n3993 0.01
R48087 vdd.n4124 vdd.n3999 0.01
R48088 vdd.n4125 vdd.n3985 0.01
R48089 vdd.n4125 vdd.n3991 0.01
R48090 vdd.n4126 vdd.n3977 0.01
R48091 vdd.n4126 vdd.n3983 0.01
R48092 vdd.n4127 vdd.n3969 0.01
R48093 vdd.n4127 vdd.n3975 0.01
R48094 vdd.n4128 vdd.n3961 0.01
R48095 vdd.n4128 vdd.n3967 0.01
R48096 vdd.n4139 vdd.n4134 0.01
R48097 vdd.n4139 vdd.n4135 0.01
R48098 vdd.n4290 vdd.n4288 0.01
R48099 vdd.n4290 vdd.n4284 0.01
R48100 vdd.n4291 vdd.n4277 0.01
R48101 vdd.n4291 vdd.n4283 0.01
R48102 vdd.n4292 vdd.n4269 0.01
R48103 vdd.n4292 vdd.n4275 0.01
R48104 vdd.n4293 vdd.n4261 0.01
R48105 vdd.n4293 vdd.n4267 0.01
R48106 vdd.n4294 vdd.n4253 0.01
R48107 vdd.n4294 vdd.n4259 0.01
R48108 vdd.n4295 vdd.n4245 0.01
R48109 vdd.n4295 vdd.n4251 0.01
R48110 vdd.n4296 vdd.n4237 0.01
R48111 vdd.n4296 vdd.n4243 0.01
R48112 vdd.n4297 vdd.n4229 0.01
R48113 vdd.n4297 vdd.n4235 0.01
R48114 vdd.n4298 vdd.n4221 0.01
R48115 vdd.n4298 vdd.n4227 0.01
R48116 vdd.n4299 vdd.n4213 0.01
R48117 vdd.n4299 vdd.n4219 0.01
R48118 vdd.n4300 vdd.n4205 0.01
R48119 vdd.n4300 vdd.n4209 0.01
R48120 vdd.n4301 vdd.n4197 0.01
R48121 vdd.n4301 vdd.n4203 0.01
R48122 vdd.n4302 vdd.n4189 0.01
R48123 vdd.n4302 vdd.n4195 0.01
R48124 vdd.n4303 vdd.n4181 0.01
R48125 vdd.n4303 vdd.n4187 0.01
R48126 vdd.n4304 vdd.n4173 0.01
R48127 vdd.n4304 vdd.n4179 0.01
R48128 vdd.n4305 vdd.n4165 0.01
R48129 vdd.n4305 vdd.n4171 0.01
R48130 vdd.n4306 vdd.n4157 0.01
R48131 vdd.n4306 vdd.n4163 0.01
R48132 vdd.n4307 vdd.n4149 0.01
R48133 vdd.n4307 vdd.n4155 0.01
R48134 vdd.n4308 vdd.n4141 0.01
R48135 vdd.n4308 vdd.n4147 0.01
R48136 vdd.n4319 vdd.n4314 0.01
R48137 vdd.n4319 vdd.n4315 0.01
R48138 vdd.n4470 vdd.n4468 0.01
R48139 vdd.n4470 vdd.n4464 0.01
R48140 vdd.n4471 vdd.n4457 0.01
R48141 vdd.n4471 vdd.n4463 0.01
R48142 vdd.n4472 vdd.n4449 0.01
R48143 vdd.n4472 vdd.n4455 0.01
R48144 vdd.n4473 vdd.n4441 0.01
R48145 vdd.n4473 vdd.n4447 0.01
R48146 vdd.n4474 vdd.n4433 0.01
R48147 vdd.n4474 vdd.n4439 0.01
R48148 vdd.n4475 vdd.n4425 0.01
R48149 vdd.n4475 vdd.n4431 0.01
R48150 vdd.n4476 vdd.n4417 0.01
R48151 vdd.n4476 vdd.n4423 0.01
R48152 vdd.n4477 vdd.n4409 0.01
R48153 vdd.n4477 vdd.n4415 0.01
R48154 vdd.n4478 vdd.n4401 0.01
R48155 vdd.n4478 vdd.n4407 0.01
R48156 vdd.n4479 vdd.n4393 0.01
R48157 vdd.n4479 vdd.n4399 0.01
R48158 vdd.n4480 vdd.n4385 0.01
R48159 vdd.n4480 vdd.n4389 0.01
R48160 vdd.n4481 vdd.n4377 0.01
R48161 vdd.n4481 vdd.n4383 0.01
R48162 vdd.n4482 vdd.n4369 0.01
R48163 vdd.n4482 vdd.n4375 0.01
R48164 vdd.n4483 vdd.n4361 0.01
R48165 vdd.n4483 vdd.n4367 0.01
R48166 vdd.n4484 vdd.n4353 0.01
R48167 vdd.n4484 vdd.n4359 0.01
R48168 vdd.n4485 vdd.n4345 0.01
R48169 vdd.n4485 vdd.n4351 0.01
R48170 vdd.n4486 vdd.n4337 0.01
R48171 vdd.n4486 vdd.n4343 0.01
R48172 vdd.n4487 vdd.n4329 0.01
R48173 vdd.n4487 vdd.n4335 0.01
R48174 vdd.n4488 vdd.n4321 0.01
R48175 vdd.n4488 vdd.n4327 0.01
R48176 vdd.n4499 vdd.n4494 0.01
R48177 vdd.n4499 vdd.n4495 0.01
R48178 vdd.n4650 vdd.n4648 0.01
R48179 vdd.n4650 vdd.n4644 0.01
R48180 vdd.n4651 vdd.n4637 0.01
R48181 vdd.n4651 vdd.n4643 0.01
R48182 vdd.n4652 vdd.n4629 0.01
R48183 vdd.n4652 vdd.n4635 0.01
R48184 vdd.n4653 vdd.n4621 0.01
R48185 vdd.n4653 vdd.n4627 0.01
R48186 vdd.n4654 vdd.n4613 0.01
R48187 vdd.n4654 vdd.n4619 0.01
R48188 vdd.n4655 vdd.n4605 0.01
R48189 vdd.n4655 vdd.n4611 0.01
R48190 vdd.n4656 vdd.n4597 0.01
R48191 vdd.n4656 vdd.n4603 0.01
R48192 vdd.n4657 vdd.n4589 0.01
R48193 vdd.n4657 vdd.n4595 0.01
R48194 vdd.n4658 vdd.n4581 0.01
R48195 vdd.n4658 vdd.n4587 0.01
R48196 vdd.n4659 vdd.n4573 0.01
R48197 vdd.n4659 vdd.n4579 0.01
R48198 vdd.n4660 vdd.n4565 0.01
R48199 vdd.n4660 vdd.n4569 0.01
R48200 vdd.n4661 vdd.n4557 0.01
R48201 vdd.n4661 vdd.n4563 0.01
R48202 vdd.n4662 vdd.n4549 0.01
R48203 vdd.n4662 vdd.n4555 0.01
R48204 vdd.n4663 vdd.n4541 0.01
R48205 vdd.n4663 vdd.n4547 0.01
R48206 vdd.n4664 vdd.n4533 0.01
R48207 vdd.n4664 vdd.n4539 0.01
R48208 vdd.n4665 vdd.n4525 0.01
R48209 vdd.n4665 vdd.n4531 0.01
R48210 vdd.n4666 vdd.n4517 0.01
R48211 vdd.n4666 vdd.n4523 0.01
R48212 vdd.n4667 vdd.n4509 0.01
R48213 vdd.n4667 vdd.n4515 0.01
R48214 vdd.n4668 vdd.n4501 0.01
R48215 vdd.n4668 vdd.n4507 0.01
R48216 vdd.n4679 vdd.n4674 0.01
R48217 vdd.n4679 vdd.n4675 0.01
R48218 vdd.n4830 vdd.n4828 0.01
R48219 vdd.n4830 vdd.n4824 0.01
R48220 vdd.n4831 vdd.n4817 0.01
R48221 vdd.n4831 vdd.n4823 0.01
R48222 vdd.n4832 vdd.n4809 0.01
R48223 vdd.n4832 vdd.n4815 0.01
R48224 vdd.n4833 vdd.n4801 0.01
R48225 vdd.n4833 vdd.n4807 0.01
R48226 vdd.n4834 vdd.n4793 0.01
R48227 vdd.n4834 vdd.n4799 0.01
R48228 vdd.n4835 vdd.n4785 0.01
R48229 vdd.n4835 vdd.n4791 0.01
R48230 vdd.n4836 vdd.n4777 0.01
R48231 vdd.n4836 vdd.n4783 0.01
R48232 vdd.n4837 vdd.n4769 0.01
R48233 vdd.n4837 vdd.n4775 0.01
R48234 vdd.n4838 vdd.n4761 0.01
R48235 vdd.n4838 vdd.n4767 0.01
R48236 vdd.n4839 vdd.n4753 0.01
R48237 vdd.n4839 vdd.n4759 0.01
R48238 vdd.n4840 vdd.n4745 0.01
R48239 vdd.n4840 vdd.n4749 0.01
R48240 vdd.n4841 vdd.n4737 0.01
R48241 vdd.n4841 vdd.n4743 0.01
R48242 vdd.n4842 vdd.n4729 0.01
R48243 vdd.n4842 vdd.n4735 0.01
R48244 vdd.n4843 vdd.n4721 0.01
R48245 vdd.n4843 vdd.n4727 0.01
R48246 vdd.n4844 vdd.n4713 0.01
R48247 vdd.n4844 vdd.n4719 0.01
R48248 vdd.n4845 vdd.n4705 0.01
R48249 vdd.n4845 vdd.n4711 0.01
R48250 vdd.n4846 vdd.n4697 0.01
R48251 vdd.n4846 vdd.n4703 0.01
R48252 vdd.n4847 vdd.n4689 0.01
R48253 vdd.n4847 vdd.n4695 0.01
R48254 vdd.n4848 vdd.n4681 0.01
R48255 vdd.n4848 vdd.n4687 0.01
R48256 vdd.n4859 vdd.n4854 0.01
R48257 vdd.n4859 vdd.n4855 0.01
R48258 vdd.n5010 vdd.n5008 0.01
R48259 vdd.n5010 vdd.n5004 0.01
R48260 vdd.n5011 vdd.n4997 0.01
R48261 vdd.n5011 vdd.n5003 0.01
R48262 vdd.n5012 vdd.n4989 0.01
R48263 vdd.n5012 vdd.n4995 0.01
R48264 vdd.n5013 vdd.n4981 0.01
R48265 vdd.n5013 vdd.n4987 0.01
R48266 vdd.n5014 vdd.n4973 0.01
R48267 vdd.n5014 vdd.n4979 0.01
R48268 vdd.n5015 vdd.n4965 0.01
R48269 vdd.n5015 vdd.n4971 0.01
R48270 vdd.n5016 vdd.n4957 0.01
R48271 vdd.n5016 vdd.n4963 0.01
R48272 vdd.n5017 vdd.n4949 0.01
R48273 vdd.n5017 vdd.n4955 0.01
R48274 vdd.n5018 vdd.n4941 0.01
R48275 vdd.n5018 vdd.n4947 0.01
R48276 vdd.n5019 vdd.n4933 0.01
R48277 vdd.n5019 vdd.n4939 0.01
R48278 vdd.n5020 vdd.n4925 0.01
R48279 vdd.n5020 vdd.n4929 0.01
R48280 vdd.n5021 vdd.n4917 0.01
R48281 vdd.n5021 vdd.n4923 0.01
R48282 vdd.n5022 vdd.n4909 0.01
R48283 vdd.n5022 vdd.n4915 0.01
R48284 vdd.n5023 vdd.n4901 0.01
R48285 vdd.n5023 vdd.n4907 0.01
R48286 vdd.n5024 vdd.n4893 0.01
R48287 vdd.n5024 vdd.n4899 0.01
R48288 vdd.n5025 vdd.n4885 0.01
R48289 vdd.n5025 vdd.n4891 0.01
R48290 vdd.n5026 vdd.n4877 0.01
R48291 vdd.n5026 vdd.n4883 0.01
R48292 vdd.n5027 vdd.n4869 0.01
R48293 vdd.n5027 vdd.n4875 0.01
R48294 vdd.n5028 vdd.n4861 0.01
R48295 vdd.n5028 vdd.n4867 0.01
R48296 vdd.n5039 vdd.n5034 0.01
R48297 vdd.n5039 vdd.n5035 0.01
R48298 vdd.n5190 vdd.n5188 0.01
R48299 vdd.n5190 vdd.n5184 0.01
R48300 vdd.n5191 vdd.n5177 0.01
R48301 vdd.n5191 vdd.n5183 0.01
R48302 vdd.n5192 vdd.n5169 0.01
R48303 vdd.n5192 vdd.n5175 0.01
R48304 vdd.n5193 vdd.n5161 0.01
R48305 vdd.n5193 vdd.n5167 0.01
R48306 vdd.n5194 vdd.n5153 0.01
R48307 vdd.n5194 vdd.n5159 0.01
R48308 vdd.n5195 vdd.n5145 0.01
R48309 vdd.n5195 vdd.n5151 0.01
R48310 vdd.n5196 vdd.n5137 0.01
R48311 vdd.n5196 vdd.n5143 0.01
R48312 vdd.n5197 vdd.n5129 0.01
R48313 vdd.n5197 vdd.n5135 0.01
R48314 vdd.n5198 vdd.n5121 0.01
R48315 vdd.n5198 vdd.n5127 0.01
R48316 vdd.n5199 vdd.n5113 0.01
R48317 vdd.n5199 vdd.n5119 0.01
R48318 vdd.n5200 vdd.n5105 0.01
R48319 vdd.n5200 vdd.n5109 0.01
R48320 vdd.n5201 vdd.n5097 0.01
R48321 vdd.n5201 vdd.n5103 0.01
R48322 vdd.n5202 vdd.n5089 0.01
R48323 vdd.n5202 vdd.n5095 0.01
R48324 vdd.n5203 vdd.n5081 0.01
R48325 vdd.n5203 vdd.n5087 0.01
R48326 vdd.n5204 vdd.n5073 0.01
R48327 vdd.n5204 vdd.n5079 0.01
R48328 vdd.n5205 vdd.n5065 0.01
R48329 vdd.n5205 vdd.n5071 0.01
R48330 vdd.n5206 vdd.n5057 0.01
R48331 vdd.n5206 vdd.n5063 0.01
R48332 vdd.n5207 vdd.n5049 0.01
R48333 vdd.n5207 vdd.n5055 0.01
R48334 vdd.n5208 vdd.n5041 0.01
R48335 vdd.n5208 vdd.n5047 0.01
R48336 vdd.n5219 vdd.n5214 0.01
R48337 vdd.n5219 vdd.n5215 0.01
R48338 vdd.n5370 vdd.n5368 0.01
R48339 vdd.n5370 vdd.n5364 0.01
R48340 vdd.n5371 vdd.n5357 0.01
R48341 vdd.n5371 vdd.n5363 0.01
R48342 vdd.n5372 vdd.n5349 0.01
R48343 vdd.n5372 vdd.n5355 0.01
R48344 vdd.n5373 vdd.n5341 0.01
R48345 vdd.n5373 vdd.n5347 0.01
R48346 vdd.n5374 vdd.n5333 0.01
R48347 vdd.n5374 vdd.n5339 0.01
R48348 vdd.n5375 vdd.n5325 0.01
R48349 vdd.n5375 vdd.n5331 0.01
R48350 vdd.n5376 vdd.n5317 0.01
R48351 vdd.n5376 vdd.n5323 0.01
R48352 vdd.n5377 vdd.n5309 0.01
R48353 vdd.n5377 vdd.n5315 0.01
R48354 vdd.n5378 vdd.n5301 0.01
R48355 vdd.n5378 vdd.n5307 0.01
R48356 vdd.n5379 vdd.n5293 0.01
R48357 vdd.n5379 vdd.n5299 0.01
R48358 vdd.n5380 vdd.n5285 0.01
R48359 vdd.n5380 vdd.n5289 0.01
R48360 vdd.n5381 vdd.n5277 0.01
R48361 vdd.n5381 vdd.n5283 0.01
R48362 vdd.n5382 vdd.n5269 0.01
R48363 vdd.n5382 vdd.n5275 0.01
R48364 vdd.n5383 vdd.n5261 0.01
R48365 vdd.n5383 vdd.n5267 0.01
R48366 vdd.n5384 vdd.n5253 0.01
R48367 vdd.n5384 vdd.n5259 0.01
R48368 vdd.n5385 vdd.n5245 0.01
R48369 vdd.n5385 vdd.n5251 0.01
R48370 vdd.n5386 vdd.n5237 0.01
R48371 vdd.n5386 vdd.n5243 0.01
R48372 vdd.n5387 vdd.n5229 0.01
R48373 vdd.n5387 vdd.n5235 0.01
R48374 vdd.n5388 vdd.n5221 0.01
R48375 vdd.n5388 vdd.n5227 0.01
R48376 vdd.n5399 vdd.n5394 0.01
R48377 vdd.n5399 vdd.n5395 0.01
R48378 vdd.n5550 vdd.n5548 0.01
R48379 vdd.n5550 vdd.n5544 0.01
R48380 vdd.n5551 vdd.n5537 0.01
R48381 vdd.n5551 vdd.n5543 0.01
R48382 vdd.n5552 vdd.n5529 0.01
R48383 vdd.n5552 vdd.n5535 0.01
R48384 vdd.n5553 vdd.n5521 0.01
R48385 vdd.n5553 vdd.n5527 0.01
R48386 vdd.n5554 vdd.n5513 0.01
R48387 vdd.n5554 vdd.n5519 0.01
R48388 vdd.n5555 vdd.n5505 0.01
R48389 vdd.n5555 vdd.n5511 0.01
R48390 vdd.n5556 vdd.n5497 0.01
R48391 vdd.n5556 vdd.n5503 0.01
R48392 vdd.n5557 vdd.n5489 0.01
R48393 vdd.n5557 vdd.n5495 0.01
R48394 vdd.n5558 vdd.n5481 0.01
R48395 vdd.n5558 vdd.n5487 0.01
R48396 vdd.n5559 vdd.n5473 0.01
R48397 vdd.n5559 vdd.n5479 0.01
R48398 vdd.n5560 vdd.n5465 0.01
R48399 vdd.n5560 vdd.n5469 0.01
R48400 vdd.n5561 vdd.n5457 0.01
R48401 vdd.n5561 vdd.n5463 0.01
R48402 vdd.n5562 vdd.n5449 0.01
R48403 vdd.n5562 vdd.n5455 0.01
R48404 vdd.n5563 vdd.n5441 0.01
R48405 vdd.n5563 vdd.n5447 0.01
R48406 vdd.n5564 vdd.n5433 0.01
R48407 vdd.n5564 vdd.n5439 0.01
R48408 vdd.n5565 vdd.n5425 0.01
R48409 vdd.n5565 vdd.n5431 0.01
R48410 vdd.n5566 vdd.n5417 0.01
R48411 vdd.n5566 vdd.n5423 0.01
R48412 vdd.n5567 vdd.n5409 0.01
R48413 vdd.n5567 vdd.n5415 0.01
R48414 vdd.n5568 vdd.n5401 0.01
R48415 vdd.n5568 vdd.n5407 0.01
R48416 vdd.n5579 vdd.n5574 0.01
R48417 vdd.n5579 vdd.n5575 0.01
R48418 vdd.n5730 vdd.n5728 0.01
R48419 vdd.n5730 vdd.n5724 0.01
R48420 vdd.n5731 vdd.n5717 0.01
R48421 vdd.n5731 vdd.n5723 0.01
R48422 vdd.n5732 vdd.n5709 0.01
R48423 vdd.n5732 vdd.n5715 0.01
R48424 vdd.n5733 vdd.n5701 0.01
R48425 vdd.n5733 vdd.n5707 0.01
R48426 vdd.n5734 vdd.n5693 0.01
R48427 vdd.n5734 vdd.n5699 0.01
R48428 vdd.n5735 vdd.n5685 0.01
R48429 vdd.n5735 vdd.n5691 0.01
R48430 vdd.n5736 vdd.n5677 0.01
R48431 vdd.n5736 vdd.n5683 0.01
R48432 vdd.n5737 vdd.n5669 0.01
R48433 vdd.n5737 vdd.n5675 0.01
R48434 vdd.n5738 vdd.n5661 0.01
R48435 vdd.n5738 vdd.n5667 0.01
R48436 vdd.n5739 vdd.n5653 0.01
R48437 vdd.n5739 vdd.n5659 0.01
R48438 vdd.n5740 vdd.n5645 0.01
R48439 vdd.n5740 vdd.n5649 0.01
R48440 vdd.n5741 vdd.n5637 0.01
R48441 vdd.n5741 vdd.n5643 0.01
R48442 vdd.n5742 vdd.n5629 0.01
R48443 vdd.n5742 vdd.n5635 0.01
R48444 vdd.n5743 vdd.n5621 0.01
R48445 vdd.n5743 vdd.n5627 0.01
R48446 vdd.n5744 vdd.n5613 0.01
R48447 vdd.n5744 vdd.n5619 0.01
R48448 vdd.n5745 vdd.n5605 0.01
R48449 vdd.n5745 vdd.n5611 0.01
R48450 vdd.n5746 vdd.n5597 0.01
R48451 vdd.n5746 vdd.n5603 0.01
R48452 vdd.n5747 vdd.n5589 0.01
R48453 vdd.n5747 vdd.n5595 0.01
R48454 vdd.n5748 vdd.n5581 0.01
R48455 vdd.n5748 vdd.n5587 0.01
R48456 vdd.n5759 vdd.n5754 0.01
R48457 vdd.n5759 vdd.n5755 0.01
R48458 vdd.n5910 vdd.n5908 0.01
R48459 vdd.n5910 vdd.n5904 0.01
R48460 vdd.n5911 vdd.n5897 0.01
R48461 vdd.n5911 vdd.n5903 0.01
R48462 vdd.n5912 vdd.n5889 0.01
R48463 vdd.n5912 vdd.n5895 0.01
R48464 vdd.n5913 vdd.n5881 0.01
R48465 vdd.n5913 vdd.n5887 0.01
R48466 vdd.n5914 vdd.n5873 0.01
R48467 vdd.n5914 vdd.n5879 0.01
R48468 vdd.n5915 vdd.n5865 0.01
R48469 vdd.n5915 vdd.n5871 0.01
R48470 vdd.n5916 vdd.n5857 0.01
R48471 vdd.n5916 vdd.n5863 0.01
R48472 vdd.n5917 vdd.n5849 0.01
R48473 vdd.n5917 vdd.n5855 0.01
R48474 vdd.n5918 vdd.n5841 0.01
R48475 vdd.n5918 vdd.n5847 0.01
R48476 vdd.n5919 vdd.n5833 0.01
R48477 vdd.n5919 vdd.n5839 0.01
R48478 vdd.n5920 vdd.n5825 0.01
R48479 vdd.n5920 vdd.n5829 0.01
R48480 vdd.n5921 vdd.n5817 0.01
R48481 vdd.n5921 vdd.n5823 0.01
R48482 vdd.n5922 vdd.n5809 0.01
R48483 vdd.n5922 vdd.n5815 0.01
R48484 vdd.n5923 vdd.n5801 0.01
R48485 vdd.n5923 vdd.n5807 0.01
R48486 vdd.n5924 vdd.n5793 0.01
R48487 vdd.n5924 vdd.n5799 0.01
R48488 vdd.n5925 vdd.n5785 0.01
R48489 vdd.n5925 vdd.n5791 0.01
R48490 vdd.n5926 vdd.n5777 0.01
R48491 vdd.n5926 vdd.n5783 0.01
R48492 vdd.n5927 vdd.n5769 0.01
R48493 vdd.n5927 vdd.n5775 0.01
R48494 vdd.n5928 vdd.n5761 0.01
R48495 vdd.n5928 vdd.n5767 0.01
R48496 vdd.n5939 vdd.n5934 0.01
R48497 vdd.n5939 vdd.n5935 0.01
R48498 vdd.n6090 vdd.n6088 0.01
R48499 vdd.n6090 vdd.n6084 0.01
R48500 vdd.n6091 vdd.n6077 0.01
R48501 vdd.n6091 vdd.n6083 0.01
R48502 vdd.n6092 vdd.n6069 0.01
R48503 vdd.n6092 vdd.n6075 0.01
R48504 vdd.n6093 vdd.n6061 0.01
R48505 vdd.n6093 vdd.n6067 0.01
R48506 vdd.n6094 vdd.n6053 0.01
R48507 vdd.n6094 vdd.n6059 0.01
R48508 vdd.n6095 vdd.n6045 0.01
R48509 vdd.n6095 vdd.n6051 0.01
R48510 vdd.n6096 vdd.n6037 0.01
R48511 vdd.n6096 vdd.n6043 0.01
R48512 vdd.n6097 vdd.n6029 0.01
R48513 vdd.n6097 vdd.n6035 0.01
R48514 vdd.n6098 vdd.n6021 0.01
R48515 vdd.n6098 vdd.n6027 0.01
R48516 vdd.n6099 vdd.n6013 0.01
R48517 vdd.n6099 vdd.n6019 0.01
R48518 vdd.n6100 vdd.n6005 0.01
R48519 vdd.n6100 vdd.n6009 0.01
R48520 vdd.n6101 vdd.n5997 0.01
R48521 vdd.n6101 vdd.n6003 0.01
R48522 vdd.n6102 vdd.n5989 0.01
R48523 vdd.n6102 vdd.n5995 0.01
R48524 vdd.n6103 vdd.n5981 0.01
R48525 vdd.n6103 vdd.n5987 0.01
R48526 vdd.n6104 vdd.n5973 0.01
R48527 vdd.n6104 vdd.n5979 0.01
R48528 vdd.n6105 vdd.n5965 0.01
R48529 vdd.n6105 vdd.n5971 0.01
R48530 vdd.n6106 vdd.n5957 0.01
R48531 vdd.n6106 vdd.n5963 0.01
R48532 vdd.n6107 vdd.n5949 0.01
R48533 vdd.n6107 vdd.n5955 0.01
R48534 vdd.n6108 vdd.n5941 0.01
R48535 vdd.n6108 vdd.n5947 0.01
R48536 vdd.n6119 vdd.n6114 0.01
R48537 vdd.n6119 vdd.n6115 0.01
R48538 vdd.n6270 vdd.n6268 0.01
R48539 vdd.n6270 vdd.n6264 0.01
R48540 vdd.n6271 vdd.n6257 0.01
R48541 vdd.n6271 vdd.n6263 0.01
R48542 vdd.n6272 vdd.n6249 0.01
R48543 vdd.n6272 vdd.n6255 0.01
R48544 vdd.n6273 vdd.n6241 0.01
R48545 vdd.n6273 vdd.n6247 0.01
R48546 vdd.n6274 vdd.n6233 0.01
R48547 vdd.n6274 vdd.n6239 0.01
R48548 vdd.n6275 vdd.n6225 0.01
R48549 vdd.n6275 vdd.n6231 0.01
R48550 vdd.n6276 vdd.n6217 0.01
R48551 vdd.n6276 vdd.n6223 0.01
R48552 vdd.n6277 vdd.n6209 0.01
R48553 vdd.n6277 vdd.n6215 0.01
R48554 vdd.n6278 vdd.n6201 0.01
R48555 vdd.n6278 vdd.n6207 0.01
R48556 vdd.n6279 vdd.n6193 0.01
R48557 vdd.n6279 vdd.n6199 0.01
R48558 vdd.n6280 vdd.n6185 0.01
R48559 vdd.n6280 vdd.n6189 0.01
R48560 vdd.n6281 vdd.n6177 0.01
R48561 vdd.n6281 vdd.n6183 0.01
R48562 vdd.n6282 vdd.n6169 0.01
R48563 vdd.n6282 vdd.n6175 0.01
R48564 vdd.n6283 vdd.n6161 0.01
R48565 vdd.n6283 vdd.n6167 0.01
R48566 vdd.n6284 vdd.n6153 0.01
R48567 vdd.n6284 vdd.n6159 0.01
R48568 vdd.n6285 vdd.n6145 0.01
R48569 vdd.n6285 vdd.n6151 0.01
R48570 vdd.n6286 vdd.n6137 0.01
R48571 vdd.n6286 vdd.n6143 0.01
R48572 vdd.n6287 vdd.n6129 0.01
R48573 vdd.n6287 vdd.n6135 0.01
R48574 vdd.n6288 vdd.n6121 0.01
R48575 vdd.n6288 vdd.n6127 0.01
R48576 vdd.n6299 vdd.n6294 0.01
R48577 vdd.n6299 vdd.n6295 0.01
R48578 vdd.n6450 vdd.n6448 0.01
R48579 vdd.n6450 vdd.n6444 0.01
R48580 vdd.n6451 vdd.n6437 0.01
R48581 vdd.n6451 vdd.n6443 0.01
R48582 vdd.n6452 vdd.n6429 0.01
R48583 vdd.n6452 vdd.n6435 0.01
R48584 vdd.n6453 vdd.n6421 0.01
R48585 vdd.n6453 vdd.n6427 0.01
R48586 vdd.n6454 vdd.n6413 0.01
R48587 vdd.n6454 vdd.n6419 0.01
R48588 vdd.n6455 vdd.n6405 0.01
R48589 vdd.n6455 vdd.n6411 0.01
R48590 vdd.n6456 vdd.n6397 0.01
R48591 vdd.n6456 vdd.n6403 0.01
R48592 vdd.n6457 vdd.n6389 0.01
R48593 vdd.n6457 vdd.n6395 0.01
R48594 vdd.n6458 vdd.n6381 0.01
R48595 vdd.n6458 vdd.n6387 0.01
R48596 vdd.n6459 vdd.n6373 0.01
R48597 vdd.n6459 vdd.n6379 0.01
R48598 vdd.n6460 vdd.n6365 0.01
R48599 vdd.n6460 vdd.n6369 0.01
R48600 vdd.n6461 vdd.n6357 0.01
R48601 vdd.n6461 vdd.n6363 0.01
R48602 vdd.n6462 vdd.n6349 0.01
R48603 vdd.n6462 vdd.n6355 0.01
R48604 vdd.n6463 vdd.n6341 0.01
R48605 vdd.n6463 vdd.n6347 0.01
R48606 vdd.n6464 vdd.n6333 0.01
R48607 vdd.n6464 vdd.n6339 0.01
R48608 vdd.n6465 vdd.n6325 0.01
R48609 vdd.n6465 vdd.n6331 0.01
R48610 vdd.n6466 vdd.n6317 0.01
R48611 vdd.n6466 vdd.n6323 0.01
R48612 vdd.n6467 vdd.n6309 0.01
R48613 vdd.n6467 vdd.n6315 0.01
R48614 vdd.n6468 vdd.n6301 0.01
R48615 vdd.n6468 vdd.n6307 0.01
R48616 vdd.n6479 vdd.n6474 0.01
R48617 vdd.n6479 vdd.n6475 0.01
R48618 vdd.n6630 vdd.n6628 0.01
R48619 vdd.n6630 vdd.n6624 0.01
R48620 vdd.n6631 vdd.n6617 0.01
R48621 vdd.n6631 vdd.n6623 0.01
R48622 vdd.n6632 vdd.n6609 0.01
R48623 vdd.n6632 vdd.n6615 0.01
R48624 vdd.n6633 vdd.n6601 0.01
R48625 vdd.n6633 vdd.n6607 0.01
R48626 vdd.n6634 vdd.n6593 0.01
R48627 vdd.n6634 vdd.n6599 0.01
R48628 vdd.n6635 vdd.n6585 0.01
R48629 vdd.n6635 vdd.n6591 0.01
R48630 vdd.n6636 vdd.n6577 0.01
R48631 vdd.n6636 vdd.n6583 0.01
R48632 vdd.n6637 vdd.n6569 0.01
R48633 vdd.n6637 vdd.n6575 0.01
R48634 vdd.n6638 vdd.n6561 0.01
R48635 vdd.n6638 vdd.n6567 0.01
R48636 vdd.n6639 vdd.n6553 0.01
R48637 vdd.n6639 vdd.n6559 0.01
R48638 vdd.n6640 vdd.n6545 0.01
R48639 vdd.n6640 vdd.n6549 0.01
R48640 vdd.n6641 vdd.n6537 0.01
R48641 vdd.n6641 vdd.n6543 0.01
R48642 vdd.n6642 vdd.n6529 0.01
R48643 vdd.n6642 vdd.n6535 0.01
R48644 vdd.n6643 vdd.n6521 0.01
R48645 vdd.n6643 vdd.n6527 0.01
R48646 vdd.n6644 vdd.n6513 0.01
R48647 vdd.n6644 vdd.n6519 0.01
R48648 vdd.n6645 vdd.n6505 0.01
R48649 vdd.n6645 vdd.n6511 0.01
R48650 vdd.n6646 vdd.n6497 0.01
R48651 vdd.n6646 vdd.n6503 0.01
R48652 vdd.n6647 vdd.n6489 0.01
R48653 vdd.n6647 vdd.n6495 0.01
R48654 vdd.n6648 vdd.n6481 0.01
R48655 vdd.n6648 vdd.n6487 0.01
R48656 vdd.n6659 vdd.n6654 0.01
R48657 vdd.n6659 vdd.n6655 0.01
R48658 vdd.n6810 vdd.n6808 0.01
R48659 vdd.n6810 vdd.n6804 0.01
R48660 vdd.n6811 vdd.n6797 0.01
R48661 vdd.n6811 vdd.n6803 0.01
R48662 vdd.n6812 vdd.n6789 0.01
R48663 vdd.n6812 vdd.n6795 0.01
R48664 vdd.n6813 vdd.n6781 0.01
R48665 vdd.n6813 vdd.n6787 0.01
R48666 vdd.n6814 vdd.n6773 0.01
R48667 vdd.n6814 vdd.n6779 0.01
R48668 vdd.n6815 vdd.n6765 0.01
R48669 vdd.n6815 vdd.n6771 0.01
R48670 vdd.n6816 vdd.n6757 0.01
R48671 vdd.n6816 vdd.n6763 0.01
R48672 vdd.n6817 vdd.n6749 0.01
R48673 vdd.n6817 vdd.n6755 0.01
R48674 vdd.n6818 vdd.n6741 0.01
R48675 vdd.n6818 vdd.n6747 0.01
R48676 vdd.n6819 vdd.n6733 0.01
R48677 vdd.n6819 vdd.n6739 0.01
R48678 vdd.n6820 vdd.n6725 0.01
R48679 vdd.n6820 vdd.n6729 0.01
R48680 vdd.n6821 vdd.n6717 0.01
R48681 vdd.n6821 vdd.n6723 0.01
R48682 vdd.n6822 vdd.n6709 0.01
R48683 vdd.n6822 vdd.n6715 0.01
R48684 vdd.n6823 vdd.n6701 0.01
R48685 vdd.n6823 vdd.n6707 0.01
R48686 vdd.n6824 vdd.n6693 0.01
R48687 vdd.n6824 vdd.n6699 0.01
R48688 vdd.n6825 vdd.n6685 0.01
R48689 vdd.n6825 vdd.n6691 0.01
R48690 vdd.n6826 vdd.n6677 0.01
R48691 vdd.n6826 vdd.n6683 0.01
R48692 vdd.n6827 vdd.n6669 0.01
R48693 vdd.n6827 vdd.n6675 0.01
R48694 vdd.n6828 vdd.n6661 0.01
R48695 vdd.n6828 vdd.n6667 0.01
R48696 vdd.n6839 vdd.n6834 0.01
R48697 vdd.n6839 vdd.n6835 0.01
R48698 vdd.n6990 vdd.n6988 0.01
R48699 vdd.n6990 vdd.n6984 0.01
R48700 vdd.n6991 vdd.n6977 0.01
R48701 vdd.n6991 vdd.n6983 0.01
R48702 vdd.n6992 vdd.n6969 0.01
R48703 vdd.n6992 vdd.n6975 0.01
R48704 vdd.n6993 vdd.n6961 0.01
R48705 vdd.n6993 vdd.n6967 0.01
R48706 vdd.n6994 vdd.n6953 0.01
R48707 vdd.n6994 vdd.n6959 0.01
R48708 vdd.n6995 vdd.n6945 0.01
R48709 vdd.n6995 vdd.n6951 0.01
R48710 vdd.n6996 vdd.n6937 0.01
R48711 vdd.n6996 vdd.n6943 0.01
R48712 vdd.n6997 vdd.n6929 0.01
R48713 vdd.n6997 vdd.n6935 0.01
R48714 vdd.n6998 vdd.n6921 0.01
R48715 vdd.n6998 vdd.n6927 0.01
R48716 vdd.n6999 vdd.n6913 0.01
R48717 vdd.n6999 vdd.n6919 0.01
R48718 vdd.n7000 vdd.n6905 0.01
R48719 vdd.n7000 vdd.n6909 0.01
R48720 vdd.n7001 vdd.n6897 0.01
R48721 vdd.n7001 vdd.n6903 0.01
R48722 vdd.n7002 vdd.n6889 0.01
R48723 vdd.n7002 vdd.n6895 0.01
R48724 vdd.n7003 vdd.n6881 0.01
R48725 vdd.n7003 vdd.n6887 0.01
R48726 vdd.n7004 vdd.n6873 0.01
R48727 vdd.n7004 vdd.n6879 0.01
R48728 vdd.n7005 vdd.n6865 0.01
R48729 vdd.n7005 vdd.n6871 0.01
R48730 vdd.n7006 vdd.n6857 0.01
R48731 vdd.n7006 vdd.n6863 0.01
R48732 vdd.n7007 vdd.n6849 0.01
R48733 vdd.n7007 vdd.n6855 0.01
R48734 vdd.n7008 vdd.n6841 0.01
R48735 vdd.n7008 vdd.n6847 0.01
R48736 vdd.n7019 vdd.n7014 0.01
R48737 vdd.n7019 vdd.n7015 0.01
R48738 vdd.n7170 vdd.n7168 0.01
R48739 vdd.n7170 vdd.n7164 0.01
R48740 vdd.n7171 vdd.n7157 0.01
R48741 vdd.n7171 vdd.n7163 0.01
R48742 vdd.n7172 vdd.n7149 0.01
R48743 vdd.n7172 vdd.n7155 0.01
R48744 vdd.n7173 vdd.n7141 0.01
R48745 vdd.n7173 vdd.n7147 0.01
R48746 vdd.n7174 vdd.n7133 0.01
R48747 vdd.n7174 vdd.n7139 0.01
R48748 vdd.n7175 vdd.n7125 0.01
R48749 vdd.n7175 vdd.n7131 0.01
R48750 vdd.n7176 vdd.n7117 0.01
R48751 vdd.n7176 vdd.n7123 0.01
R48752 vdd.n7177 vdd.n7109 0.01
R48753 vdd.n7177 vdd.n7115 0.01
R48754 vdd.n7178 vdd.n7101 0.01
R48755 vdd.n7178 vdd.n7107 0.01
R48756 vdd.n7179 vdd.n7093 0.01
R48757 vdd.n7179 vdd.n7099 0.01
R48758 vdd.n7180 vdd.n7085 0.01
R48759 vdd.n7180 vdd.n7089 0.01
R48760 vdd.n7181 vdd.n7077 0.01
R48761 vdd.n7181 vdd.n7083 0.01
R48762 vdd.n7182 vdd.n7069 0.01
R48763 vdd.n7182 vdd.n7075 0.01
R48764 vdd.n7183 vdd.n7061 0.01
R48765 vdd.n7183 vdd.n7067 0.01
R48766 vdd.n7184 vdd.n7053 0.01
R48767 vdd.n7184 vdd.n7059 0.01
R48768 vdd.n7185 vdd.n7045 0.01
R48769 vdd.n7185 vdd.n7051 0.01
R48770 vdd.n7186 vdd.n7037 0.01
R48771 vdd.n7186 vdd.n7043 0.01
R48772 vdd.n7187 vdd.n7029 0.01
R48773 vdd.n7187 vdd.n7035 0.01
R48774 vdd.n7188 vdd.n7021 0.01
R48775 vdd.n7188 vdd.n7027 0.01
R48776 vdd.n7199 vdd.n7194 0.01
R48777 vdd.n7199 vdd.n7195 0.01
R48778 vdd.n7350 vdd.n7348 0.01
R48779 vdd.n7350 vdd.n7344 0.01
R48780 vdd.n7351 vdd.n7337 0.01
R48781 vdd.n7351 vdd.n7343 0.01
R48782 vdd.n7352 vdd.n7329 0.01
R48783 vdd.n7352 vdd.n7335 0.01
R48784 vdd.n7353 vdd.n7321 0.01
R48785 vdd.n7353 vdd.n7327 0.01
R48786 vdd.n7354 vdd.n7313 0.01
R48787 vdd.n7354 vdd.n7319 0.01
R48788 vdd.n7355 vdd.n7305 0.01
R48789 vdd.n7355 vdd.n7311 0.01
R48790 vdd.n7356 vdd.n7297 0.01
R48791 vdd.n7356 vdd.n7303 0.01
R48792 vdd.n7357 vdd.n7289 0.01
R48793 vdd.n7357 vdd.n7295 0.01
R48794 vdd.n7358 vdd.n7281 0.01
R48795 vdd.n7358 vdd.n7287 0.01
R48796 vdd.n7359 vdd.n7273 0.01
R48797 vdd.n7359 vdd.n7279 0.01
R48798 vdd.n7360 vdd.n7265 0.01
R48799 vdd.n7360 vdd.n7269 0.01
R48800 vdd.n7361 vdd.n7257 0.01
R48801 vdd.n7361 vdd.n7263 0.01
R48802 vdd.n7362 vdd.n7249 0.01
R48803 vdd.n7362 vdd.n7255 0.01
R48804 vdd.n7363 vdd.n7241 0.01
R48805 vdd.n7363 vdd.n7247 0.01
R48806 vdd.n7364 vdd.n7233 0.01
R48807 vdd.n7364 vdd.n7239 0.01
R48808 vdd.n7365 vdd.n7225 0.01
R48809 vdd.n7365 vdd.n7231 0.01
R48810 vdd.n7366 vdd.n7217 0.01
R48811 vdd.n7366 vdd.n7223 0.01
R48812 vdd.n7367 vdd.n7209 0.01
R48813 vdd.n7367 vdd.n7215 0.01
R48814 vdd.n7368 vdd.n7201 0.01
R48815 vdd.n7368 vdd.n7207 0.01
R48816 vdd.n7379 vdd.n7374 0.01
R48817 vdd.n7379 vdd.n7375 0.01
R48818 vdd.n7530 vdd.n7528 0.01
R48819 vdd.n7530 vdd.n7524 0.01
R48820 vdd.n7531 vdd.n7517 0.01
R48821 vdd.n7531 vdd.n7523 0.01
R48822 vdd.n7532 vdd.n7509 0.01
R48823 vdd.n7532 vdd.n7515 0.01
R48824 vdd.n7533 vdd.n7501 0.01
R48825 vdd.n7533 vdd.n7507 0.01
R48826 vdd.n7534 vdd.n7493 0.01
R48827 vdd.n7534 vdd.n7499 0.01
R48828 vdd.n7535 vdd.n7485 0.01
R48829 vdd.n7535 vdd.n7491 0.01
R48830 vdd.n7536 vdd.n7477 0.01
R48831 vdd.n7536 vdd.n7483 0.01
R48832 vdd.n7537 vdd.n7469 0.01
R48833 vdd.n7537 vdd.n7475 0.01
R48834 vdd.n7538 vdd.n7461 0.01
R48835 vdd.n7538 vdd.n7467 0.01
R48836 vdd.n7539 vdd.n7453 0.01
R48837 vdd.n7539 vdd.n7459 0.01
R48838 vdd.n7540 vdd.n7445 0.01
R48839 vdd.n7540 vdd.n7449 0.01
R48840 vdd.n7541 vdd.n7437 0.01
R48841 vdd.n7541 vdd.n7443 0.01
R48842 vdd.n7542 vdd.n7429 0.01
R48843 vdd.n7542 vdd.n7435 0.01
R48844 vdd.n7543 vdd.n7421 0.01
R48845 vdd.n7543 vdd.n7427 0.01
R48846 vdd.n7544 vdd.n7413 0.01
R48847 vdd.n7544 vdd.n7419 0.01
R48848 vdd.n7545 vdd.n7405 0.01
R48849 vdd.n7545 vdd.n7411 0.01
R48850 vdd.n7546 vdd.n7397 0.01
R48851 vdd.n7546 vdd.n7403 0.01
R48852 vdd.n7547 vdd.n7389 0.01
R48853 vdd.n7547 vdd.n7395 0.01
R48854 vdd.n7548 vdd.n7381 0.01
R48855 vdd.n7548 vdd.n7387 0.01
R48856 vdd.n7559 vdd.n7554 0.01
R48857 vdd.n7559 vdd.n7555 0.01
R48858 vdd.n7710 vdd.n7708 0.01
R48859 vdd.n7710 vdd.n7704 0.01
R48860 vdd.n7711 vdd.n7697 0.01
R48861 vdd.n7711 vdd.n7703 0.01
R48862 vdd.n7712 vdd.n7689 0.01
R48863 vdd.n7712 vdd.n7695 0.01
R48864 vdd.n7713 vdd.n7681 0.01
R48865 vdd.n7713 vdd.n7687 0.01
R48866 vdd.n7714 vdd.n7673 0.01
R48867 vdd.n7714 vdd.n7679 0.01
R48868 vdd.n7715 vdd.n7665 0.01
R48869 vdd.n7715 vdd.n7671 0.01
R48870 vdd.n7716 vdd.n7657 0.01
R48871 vdd.n7716 vdd.n7663 0.01
R48872 vdd.n7717 vdd.n7649 0.01
R48873 vdd.n7717 vdd.n7655 0.01
R48874 vdd.n7718 vdd.n7641 0.01
R48875 vdd.n7718 vdd.n7647 0.01
R48876 vdd.n7719 vdd.n7633 0.01
R48877 vdd.n7719 vdd.n7639 0.01
R48878 vdd.n7720 vdd.n7625 0.01
R48879 vdd.n7720 vdd.n7629 0.01
R48880 vdd.n7721 vdd.n7617 0.01
R48881 vdd.n7721 vdd.n7623 0.01
R48882 vdd.n7722 vdd.n7609 0.01
R48883 vdd.n7722 vdd.n7615 0.01
R48884 vdd.n7723 vdd.n7601 0.01
R48885 vdd.n7723 vdd.n7607 0.01
R48886 vdd.n7724 vdd.n7593 0.01
R48887 vdd.n7724 vdd.n7599 0.01
R48888 vdd.n7725 vdd.n7585 0.01
R48889 vdd.n7725 vdd.n7591 0.01
R48890 vdd.n7726 vdd.n7577 0.01
R48891 vdd.n7726 vdd.n7583 0.01
R48892 vdd.n7727 vdd.n7569 0.01
R48893 vdd.n7727 vdd.n7575 0.01
R48894 vdd.n7728 vdd.n7561 0.01
R48895 vdd.n7728 vdd.n7567 0.01
R48896 vdd.n7739 vdd.n7734 0.01
R48897 vdd.n7739 vdd.n7735 0.01
R48898 vdd.n7890 vdd.n7888 0.01
R48899 vdd.n7890 vdd.n7884 0.01
R48900 vdd.n7891 vdd.n7877 0.01
R48901 vdd.n7891 vdd.n7883 0.01
R48902 vdd.n7892 vdd.n7869 0.01
R48903 vdd.n7892 vdd.n7875 0.01
R48904 vdd.n7893 vdd.n7861 0.01
R48905 vdd.n7893 vdd.n7867 0.01
R48906 vdd.n7894 vdd.n7853 0.01
R48907 vdd.n7894 vdd.n7859 0.01
R48908 vdd.n7895 vdd.n7845 0.01
R48909 vdd.n7895 vdd.n7851 0.01
R48910 vdd.n7896 vdd.n7837 0.01
R48911 vdd.n7896 vdd.n7843 0.01
R48912 vdd.n7897 vdd.n7829 0.01
R48913 vdd.n7897 vdd.n7835 0.01
R48914 vdd.n7898 vdd.n7821 0.01
R48915 vdd.n7898 vdd.n7827 0.01
R48916 vdd.n7899 vdd.n7813 0.01
R48917 vdd.n7899 vdd.n7819 0.01
R48918 vdd.n7900 vdd.n7805 0.01
R48919 vdd.n7900 vdd.n7809 0.01
R48920 vdd.n7901 vdd.n7797 0.01
R48921 vdd.n7901 vdd.n7803 0.01
R48922 vdd.n7902 vdd.n7789 0.01
R48923 vdd.n7902 vdd.n7795 0.01
R48924 vdd.n7903 vdd.n7781 0.01
R48925 vdd.n7903 vdd.n7787 0.01
R48926 vdd.n7904 vdd.n7773 0.01
R48927 vdd.n7904 vdd.n7779 0.01
R48928 vdd.n7905 vdd.n7765 0.01
R48929 vdd.n7905 vdd.n7771 0.01
R48930 vdd.n7906 vdd.n7757 0.01
R48931 vdd.n7906 vdd.n7763 0.01
R48932 vdd.n7907 vdd.n7749 0.01
R48933 vdd.n7907 vdd.n7755 0.01
R48934 vdd.n7908 vdd.n7741 0.01
R48935 vdd.n7908 vdd.n7747 0.01
R48936 vdd.n7919 vdd.n7914 0.01
R48937 vdd.n7919 vdd.n7915 0.01
R48938 vdd.n8070 vdd.n8068 0.01
R48939 vdd.n8070 vdd.n8064 0.01
R48940 vdd.n8071 vdd.n8057 0.01
R48941 vdd.n8071 vdd.n8063 0.01
R48942 vdd.n8072 vdd.n8049 0.01
R48943 vdd.n8072 vdd.n8055 0.01
R48944 vdd.n8073 vdd.n8041 0.01
R48945 vdd.n8073 vdd.n8047 0.01
R48946 vdd.n8074 vdd.n8033 0.01
R48947 vdd.n8074 vdd.n8039 0.01
R48948 vdd.n8075 vdd.n8025 0.01
R48949 vdd.n8075 vdd.n8031 0.01
R48950 vdd.n8076 vdd.n8017 0.01
R48951 vdd.n8076 vdd.n8023 0.01
R48952 vdd.n8077 vdd.n8009 0.01
R48953 vdd.n8077 vdd.n8015 0.01
R48954 vdd.n8078 vdd.n8001 0.01
R48955 vdd.n8078 vdd.n8007 0.01
R48956 vdd.n8079 vdd.n7993 0.01
R48957 vdd.n8079 vdd.n7999 0.01
R48958 vdd.n8080 vdd.n7985 0.01
R48959 vdd.n8080 vdd.n7989 0.01
R48960 vdd.n8081 vdd.n7977 0.01
R48961 vdd.n8081 vdd.n7983 0.01
R48962 vdd.n8082 vdd.n7969 0.01
R48963 vdd.n8082 vdd.n7975 0.01
R48964 vdd.n8083 vdd.n7961 0.01
R48965 vdd.n8083 vdd.n7967 0.01
R48966 vdd.n8084 vdd.n7953 0.01
R48967 vdd.n8084 vdd.n7959 0.01
R48968 vdd.n8085 vdd.n7945 0.01
R48969 vdd.n8085 vdd.n7951 0.01
R48970 vdd.n8086 vdd.n7937 0.01
R48971 vdd.n8086 vdd.n7943 0.01
R48972 vdd.n8087 vdd.n7929 0.01
R48973 vdd.n8087 vdd.n7935 0.01
R48974 vdd.n8088 vdd.n7921 0.01
R48975 vdd.n8088 vdd.n7927 0.01
R48976 vdd.n8099 vdd.n8094 0.01
R48977 vdd.n8099 vdd.n8095 0.01
R48978 vdd.n8250 vdd.n8248 0.01
R48979 vdd.n8250 vdd.n8244 0.01
R48980 vdd.n8251 vdd.n8237 0.01
R48981 vdd.n8251 vdd.n8243 0.01
R48982 vdd.n8252 vdd.n8229 0.01
R48983 vdd.n8252 vdd.n8235 0.01
R48984 vdd.n8253 vdd.n8221 0.01
R48985 vdd.n8253 vdd.n8227 0.01
R48986 vdd.n8254 vdd.n8213 0.01
R48987 vdd.n8254 vdd.n8219 0.01
R48988 vdd.n8255 vdd.n8205 0.01
R48989 vdd.n8255 vdd.n8211 0.01
R48990 vdd.n8256 vdd.n8197 0.01
R48991 vdd.n8256 vdd.n8203 0.01
R48992 vdd.n8257 vdd.n8189 0.01
R48993 vdd.n8257 vdd.n8195 0.01
R48994 vdd.n8258 vdd.n8181 0.01
R48995 vdd.n8258 vdd.n8187 0.01
R48996 vdd.n8259 vdd.n8173 0.01
R48997 vdd.n8259 vdd.n8179 0.01
R48998 vdd.n8260 vdd.n8165 0.01
R48999 vdd.n8260 vdd.n8169 0.01
R49000 vdd.n8261 vdd.n8157 0.01
R49001 vdd.n8261 vdd.n8163 0.01
R49002 vdd.n8262 vdd.n8149 0.01
R49003 vdd.n8262 vdd.n8155 0.01
R49004 vdd.n8263 vdd.n8141 0.01
R49005 vdd.n8263 vdd.n8147 0.01
R49006 vdd.n8264 vdd.n8133 0.01
R49007 vdd.n8264 vdd.n8139 0.01
R49008 vdd.n8265 vdd.n8125 0.01
R49009 vdd.n8265 vdd.n8131 0.01
R49010 vdd.n8266 vdd.n8117 0.01
R49011 vdd.n8266 vdd.n8123 0.01
R49012 vdd.n8267 vdd.n8109 0.01
R49013 vdd.n8267 vdd.n8115 0.01
R49014 vdd.n8268 vdd.n8101 0.01
R49015 vdd.n8268 vdd.n8107 0.01
R49016 vdd.n8279 vdd.n8274 0.01
R49017 vdd.n8279 vdd.n8275 0.01
R49018 vdd.n8430 vdd.n8428 0.01
R49019 vdd.n8430 vdd.n8424 0.01
R49020 vdd.n8431 vdd.n8417 0.01
R49021 vdd.n8431 vdd.n8423 0.01
R49022 vdd.n8432 vdd.n8409 0.01
R49023 vdd.n8432 vdd.n8415 0.01
R49024 vdd.n8433 vdd.n8401 0.01
R49025 vdd.n8433 vdd.n8407 0.01
R49026 vdd.n8434 vdd.n8393 0.01
R49027 vdd.n8434 vdd.n8399 0.01
R49028 vdd.n8435 vdd.n8385 0.01
R49029 vdd.n8435 vdd.n8391 0.01
R49030 vdd.n8436 vdd.n8377 0.01
R49031 vdd.n8436 vdd.n8383 0.01
R49032 vdd.n8437 vdd.n8369 0.01
R49033 vdd.n8437 vdd.n8375 0.01
R49034 vdd.n8438 vdd.n8361 0.01
R49035 vdd.n8438 vdd.n8367 0.01
R49036 vdd.n8439 vdd.n8353 0.01
R49037 vdd.n8439 vdd.n8359 0.01
R49038 vdd.n8440 vdd.n8345 0.01
R49039 vdd.n8440 vdd.n8349 0.01
R49040 vdd.n8441 vdd.n8337 0.01
R49041 vdd.n8441 vdd.n8343 0.01
R49042 vdd.n8442 vdd.n8329 0.01
R49043 vdd.n8442 vdd.n8335 0.01
R49044 vdd.n8443 vdd.n8321 0.01
R49045 vdd.n8443 vdd.n8327 0.01
R49046 vdd.n8444 vdd.n8313 0.01
R49047 vdd.n8444 vdd.n8319 0.01
R49048 vdd.n8445 vdd.n8305 0.01
R49049 vdd.n8445 vdd.n8311 0.01
R49050 vdd.n8446 vdd.n8297 0.01
R49051 vdd.n8446 vdd.n8303 0.01
R49052 vdd.n8447 vdd.n8289 0.01
R49053 vdd.n8447 vdd.n8295 0.01
R49054 vdd.n8448 vdd.n8281 0.01
R49055 vdd.n8448 vdd.n8287 0.01
R49056 vdd.n8459 vdd.n8454 0.01
R49057 vdd.n8459 vdd.n8455 0.01
R49058 vdd.n8610 vdd.n8608 0.01
R49059 vdd.n8610 vdd.n8604 0.01
R49060 vdd.n8611 vdd.n8597 0.01
R49061 vdd.n8611 vdd.n8603 0.01
R49062 vdd.n8612 vdd.n8589 0.01
R49063 vdd.n8612 vdd.n8595 0.01
R49064 vdd.n8613 vdd.n8581 0.01
R49065 vdd.n8613 vdd.n8587 0.01
R49066 vdd.n8614 vdd.n8573 0.01
R49067 vdd.n8614 vdd.n8579 0.01
R49068 vdd.n8615 vdd.n8565 0.01
R49069 vdd.n8615 vdd.n8571 0.01
R49070 vdd.n8616 vdd.n8557 0.01
R49071 vdd.n8616 vdd.n8563 0.01
R49072 vdd.n8617 vdd.n8549 0.01
R49073 vdd.n8617 vdd.n8555 0.01
R49074 vdd.n8618 vdd.n8541 0.01
R49075 vdd.n8618 vdd.n8547 0.01
R49076 vdd.n8619 vdd.n8533 0.01
R49077 vdd.n8619 vdd.n8539 0.01
R49078 vdd.n8620 vdd.n8525 0.01
R49079 vdd.n8620 vdd.n8529 0.01
R49080 vdd.n8621 vdd.n8517 0.01
R49081 vdd.n8621 vdd.n8523 0.01
R49082 vdd.n8622 vdd.n8509 0.01
R49083 vdd.n8622 vdd.n8515 0.01
R49084 vdd.n8623 vdd.n8501 0.01
R49085 vdd.n8623 vdd.n8507 0.01
R49086 vdd.n8624 vdd.n8493 0.01
R49087 vdd.n8624 vdd.n8499 0.01
R49088 vdd.n8625 vdd.n8485 0.01
R49089 vdd.n8625 vdd.n8491 0.01
R49090 vdd.n8626 vdd.n8477 0.01
R49091 vdd.n8626 vdd.n8483 0.01
R49092 vdd.n8627 vdd.n8469 0.01
R49093 vdd.n8627 vdd.n8475 0.01
R49094 vdd.n8628 vdd.n8461 0.01
R49095 vdd.n8628 vdd.n8467 0.01
R49096 vdd.n8639 vdd.n8634 0.01
R49097 vdd.n8639 vdd.n8635 0.01
R49098 vdd.n8790 vdd.n8788 0.01
R49099 vdd.n8790 vdd.n8784 0.01
R49100 vdd.n8791 vdd.n8777 0.01
R49101 vdd.n8791 vdd.n8783 0.01
R49102 vdd.n8792 vdd.n8769 0.01
R49103 vdd.n8792 vdd.n8775 0.01
R49104 vdd.n8793 vdd.n8761 0.01
R49105 vdd.n8793 vdd.n8767 0.01
R49106 vdd.n8794 vdd.n8753 0.01
R49107 vdd.n8794 vdd.n8759 0.01
R49108 vdd.n8795 vdd.n8745 0.01
R49109 vdd.n8795 vdd.n8751 0.01
R49110 vdd.n8796 vdd.n8737 0.01
R49111 vdd.n8796 vdd.n8743 0.01
R49112 vdd.n8797 vdd.n8729 0.01
R49113 vdd.n8797 vdd.n8735 0.01
R49114 vdd.n8798 vdd.n8721 0.01
R49115 vdd.n8798 vdd.n8727 0.01
R49116 vdd.n8799 vdd.n8713 0.01
R49117 vdd.n8799 vdd.n8719 0.01
R49118 vdd.n8800 vdd.n8705 0.01
R49119 vdd.n8800 vdd.n8709 0.01
R49120 vdd.n8801 vdd.n8697 0.01
R49121 vdd.n8801 vdd.n8703 0.01
R49122 vdd.n8802 vdd.n8689 0.01
R49123 vdd.n8802 vdd.n8695 0.01
R49124 vdd.n8803 vdd.n8681 0.01
R49125 vdd.n8803 vdd.n8687 0.01
R49126 vdd.n8804 vdd.n8673 0.01
R49127 vdd.n8804 vdd.n8679 0.01
R49128 vdd.n8805 vdd.n8665 0.01
R49129 vdd.n8805 vdd.n8671 0.01
R49130 vdd.n8806 vdd.n8657 0.01
R49131 vdd.n8806 vdd.n8663 0.01
R49132 vdd.n8807 vdd.n8649 0.01
R49133 vdd.n8807 vdd.n8655 0.01
R49134 vdd.n8808 vdd.n8641 0.01
R49135 vdd.n8808 vdd.n8647 0.01
R49136 vdd.n8819 vdd.n8814 0.01
R49137 vdd.n8819 vdd.n8815 0.01
R49138 vdd.n8970 vdd.n8968 0.01
R49139 vdd.n8970 vdd.n8964 0.01
R49140 vdd.n8971 vdd.n8957 0.01
R49141 vdd.n8971 vdd.n8963 0.01
R49142 vdd.n8972 vdd.n8949 0.01
R49143 vdd.n8972 vdd.n8955 0.01
R49144 vdd.n8973 vdd.n8941 0.01
R49145 vdd.n8973 vdd.n8947 0.01
R49146 vdd.n8974 vdd.n8933 0.01
R49147 vdd.n8974 vdd.n8939 0.01
R49148 vdd.n8975 vdd.n8925 0.01
R49149 vdd.n8975 vdd.n8931 0.01
R49150 vdd.n8976 vdd.n8917 0.01
R49151 vdd.n8976 vdd.n8923 0.01
R49152 vdd.n8977 vdd.n8909 0.01
R49153 vdd.n8977 vdd.n8915 0.01
R49154 vdd.n8978 vdd.n8901 0.01
R49155 vdd.n8978 vdd.n8907 0.01
R49156 vdd.n8979 vdd.n8893 0.01
R49157 vdd.n8979 vdd.n8899 0.01
R49158 vdd.n8980 vdd.n8885 0.01
R49159 vdd.n8980 vdd.n8889 0.01
R49160 vdd.n8981 vdd.n8877 0.01
R49161 vdd.n8981 vdd.n8883 0.01
R49162 vdd.n8982 vdd.n8869 0.01
R49163 vdd.n8982 vdd.n8875 0.01
R49164 vdd.n8983 vdd.n8861 0.01
R49165 vdd.n8983 vdd.n8867 0.01
R49166 vdd.n8984 vdd.n8853 0.01
R49167 vdd.n8984 vdd.n8859 0.01
R49168 vdd.n8985 vdd.n8845 0.01
R49169 vdd.n8985 vdd.n8851 0.01
R49170 vdd.n8986 vdd.n8837 0.01
R49171 vdd.n8986 vdd.n8843 0.01
R49172 vdd.n8987 vdd.n8829 0.01
R49173 vdd.n8987 vdd.n8835 0.01
R49174 vdd.n8988 vdd.n8821 0.01
R49175 vdd.n8988 vdd.n8827 0.01
R49176 vdd.n8999 vdd.n8994 0.01
R49177 vdd.n8999 vdd.n8995 0.01
R49178 vdd.n9150 vdd.n9148 0.01
R49179 vdd.n9150 vdd.n9144 0.01
R49180 vdd.n9151 vdd.n9137 0.01
R49181 vdd.n9151 vdd.n9143 0.01
R49182 vdd.n9152 vdd.n9129 0.01
R49183 vdd.n9152 vdd.n9135 0.01
R49184 vdd.n9153 vdd.n9121 0.01
R49185 vdd.n9153 vdd.n9127 0.01
R49186 vdd.n9154 vdd.n9113 0.01
R49187 vdd.n9154 vdd.n9119 0.01
R49188 vdd.n9155 vdd.n9105 0.01
R49189 vdd.n9155 vdd.n9111 0.01
R49190 vdd.n9156 vdd.n9097 0.01
R49191 vdd.n9156 vdd.n9103 0.01
R49192 vdd.n9157 vdd.n9089 0.01
R49193 vdd.n9157 vdd.n9095 0.01
R49194 vdd.n9158 vdd.n9081 0.01
R49195 vdd.n9158 vdd.n9087 0.01
R49196 vdd.n9159 vdd.n9073 0.01
R49197 vdd.n9159 vdd.n9079 0.01
R49198 vdd.n9160 vdd.n9065 0.01
R49199 vdd.n9160 vdd.n9069 0.01
R49200 vdd.n9161 vdd.n9057 0.01
R49201 vdd.n9161 vdd.n9063 0.01
R49202 vdd.n9162 vdd.n9049 0.01
R49203 vdd.n9162 vdd.n9055 0.01
R49204 vdd.n9163 vdd.n9041 0.01
R49205 vdd.n9163 vdd.n9047 0.01
R49206 vdd.n9164 vdd.n9033 0.01
R49207 vdd.n9164 vdd.n9039 0.01
R49208 vdd.n9165 vdd.n9025 0.01
R49209 vdd.n9165 vdd.n9031 0.01
R49210 vdd.n9166 vdd.n9017 0.01
R49211 vdd.n9166 vdd.n9023 0.01
R49212 vdd.n9167 vdd.n9009 0.01
R49213 vdd.n9167 vdd.n9015 0.01
R49214 vdd.n9168 vdd.n9001 0.01
R49215 vdd.n9168 vdd.n9007 0.01
R49216 vdd.n9179 vdd.n9174 0.01
R49217 vdd.n9179 vdd.n9175 0.01
R49218 vdd.n9330 vdd.n9328 0.01
R49219 vdd.n9330 vdd.n9324 0.01
R49220 vdd.n9331 vdd.n9317 0.01
R49221 vdd.n9331 vdd.n9323 0.01
R49222 vdd.n9332 vdd.n9309 0.01
R49223 vdd.n9332 vdd.n9315 0.01
R49224 vdd.n9333 vdd.n9301 0.01
R49225 vdd.n9333 vdd.n9307 0.01
R49226 vdd.n9334 vdd.n9293 0.01
R49227 vdd.n9334 vdd.n9299 0.01
R49228 vdd.n9335 vdd.n9285 0.01
R49229 vdd.n9335 vdd.n9291 0.01
R49230 vdd.n9336 vdd.n9277 0.01
R49231 vdd.n9336 vdd.n9283 0.01
R49232 vdd.n9337 vdd.n9269 0.01
R49233 vdd.n9337 vdd.n9275 0.01
R49234 vdd.n9338 vdd.n9261 0.01
R49235 vdd.n9338 vdd.n9267 0.01
R49236 vdd.n9339 vdd.n9253 0.01
R49237 vdd.n9339 vdd.n9259 0.01
R49238 vdd.n9340 vdd.n9245 0.01
R49239 vdd.n9340 vdd.n9249 0.01
R49240 vdd.n9341 vdd.n9237 0.01
R49241 vdd.n9341 vdd.n9243 0.01
R49242 vdd.n9342 vdd.n9229 0.01
R49243 vdd.n9342 vdd.n9235 0.01
R49244 vdd.n9343 vdd.n9221 0.01
R49245 vdd.n9343 vdd.n9227 0.01
R49246 vdd.n9344 vdd.n9213 0.01
R49247 vdd.n9344 vdd.n9219 0.01
R49248 vdd.n9345 vdd.n9205 0.01
R49249 vdd.n9345 vdd.n9211 0.01
R49250 vdd.n9346 vdd.n9197 0.01
R49251 vdd.n9346 vdd.n9203 0.01
R49252 vdd.n9347 vdd.n9189 0.01
R49253 vdd.n9347 vdd.n9195 0.01
R49254 vdd.n9348 vdd.n9181 0.01
R49255 vdd.n9348 vdd.n9187 0.01
R49256 vdd.n9359 vdd.n9354 0.01
R49257 vdd.n9359 vdd.n9355 0.01
R49258 vdd.n9510 vdd.n9508 0.01
R49259 vdd.n9510 vdd.n9504 0.01
R49260 vdd.n9511 vdd.n9497 0.01
R49261 vdd.n9511 vdd.n9503 0.01
R49262 vdd.n9512 vdd.n9489 0.01
R49263 vdd.n9512 vdd.n9495 0.01
R49264 vdd.n9513 vdd.n9481 0.01
R49265 vdd.n9513 vdd.n9487 0.01
R49266 vdd.n9514 vdd.n9473 0.01
R49267 vdd.n9514 vdd.n9479 0.01
R49268 vdd.n9515 vdd.n9465 0.01
R49269 vdd.n9515 vdd.n9471 0.01
R49270 vdd.n9516 vdd.n9457 0.01
R49271 vdd.n9516 vdd.n9463 0.01
R49272 vdd.n9517 vdd.n9449 0.01
R49273 vdd.n9517 vdd.n9455 0.01
R49274 vdd.n9518 vdd.n9441 0.01
R49275 vdd.n9518 vdd.n9447 0.01
R49276 vdd.n9519 vdd.n9433 0.01
R49277 vdd.n9519 vdd.n9439 0.01
R49278 vdd.n9520 vdd.n9425 0.01
R49279 vdd.n9520 vdd.n9429 0.01
R49280 vdd.n9521 vdd.n9417 0.01
R49281 vdd.n9521 vdd.n9423 0.01
R49282 vdd.n9522 vdd.n9409 0.01
R49283 vdd.n9522 vdd.n9415 0.01
R49284 vdd.n9523 vdd.n9401 0.01
R49285 vdd.n9523 vdd.n9407 0.01
R49286 vdd.n9524 vdd.n9393 0.01
R49287 vdd.n9524 vdd.n9399 0.01
R49288 vdd.n9525 vdd.n9385 0.01
R49289 vdd.n9525 vdd.n9391 0.01
R49290 vdd.n9526 vdd.n9377 0.01
R49291 vdd.n9526 vdd.n9383 0.01
R49292 vdd.n9527 vdd.n9369 0.01
R49293 vdd.n9527 vdd.n9375 0.01
R49294 vdd.n9528 vdd.n9361 0.01
R49295 vdd.n9528 vdd.n9367 0.01
R49296 vdd.n9539 vdd.n9534 0.01
R49297 vdd.n9539 vdd.n9535 0.01
R49298 vdd.n9690 vdd.n9688 0.01
R49299 vdd.n9690 vdd.n9684 0.01
R49300 vdd.n9691 vdd.n9677 0.01
R49301 vdd.n9691 vdd.n9683 0.01
R49302 vdd.n9692 vdd.n9669 0.01
R49303 vdd.n9692 vdd.n9675 0.01
R49304 vdd.n9693 vdd.n9661 0.01
R49305 vdd.n9693 vdd.n9667 0.01
R49306 vdd.n9694 vdd.n9653 0.01
R49307 vdd.n9694 vdd.n9659 0.01
R49308 vdd.n9695 vdd.n9645 0.01
R49309 vdd.n9695 vdd.n9651 0.01
R49310 vdd.n9696 vdd.n9637 0.01
R49311 vdd.n9696 vdd.n9643 0.01
R49312 vdd.n9697 vdd.n9629 0.01
R49313 vdd.n9697 vdd.n9635 0.01
R49314 vdd.n9698 vdd.n9621 0.01
R49315 vdd.n9698 vdd.n9627 0.01
R49316 vdd.n9699 vdd.n9613 0.01
R49317 vdd.n9699 vdd.n9619 0.01
R49318 vdd.n9700 vdd.n9605 0.01
R49319 vdd.n9700 vdd.n9609 0.01
R49320 vdd.n9701 vdd.n9597 0.01
R49321 vdd.n9701 vdd.n9603 0.01
R49322 vdd.n9702 vdd.n9589 0.01
R49323 vdd.n9702 vdd.n9595 0.01
R49324 vdd.n9703 vdd.n9581 0.01
R49325 vdd.n9703 vdd.n9587 0.01
R49326 vdd.n9704 vdd.n9573 0.01
R49327 vdd.n9704 vdd.n9579 0.01
R49328 vdd.n9705 vdd.n9565 0.01
R49329 vdd.n9705 vdd.n9571 0.01
R49330 vdd.n9706 vdd.n9557 0.01
R49331 vdd.n9706 vdd.n9563 0.01
R49332 vdd.n9707 vdd.n9549 0.01
R49333 vdd.n9707 vdd.n9555 0.01
R49334 vdd.n9708 vdd.n9541 0.01
R49335 vdd.n9708 vdd.n9547 0.01
R49336 vdd.n9719 vdd.n9714 0.01
R49337 vdd.n9719 vdd.n9715 0.01
R49338 vdd.n9870 vdd.n9868 0.01
R49339 vdd.n9870 vdd.n9864 0.01
R49340 vdd.n9871 vdd.n9857 0.01
R49341 vdd.n9871 vdd.n9863 0.01
R49342 vdd.n9872 vdd.n9849 0.01
R49343 vdd.n9872 vdd.n9855 0.01
R49344 vdd.n9873 vdd.n9841 0.01
R49345 vdd.n9873 vdd.n9847 0.01
R49346 vdd.n9874 vdd.n9833 0.01
R49347 vdd.n9874 vdd.n9839 0.01
R49348 vdd.n9875 vdd.n9825 0.01
R49349 vdd.n9875 vdd.n9831 0.01
R49350 vdd.n9876 vdd.n9817 0.01
R49351 vdd.n9876 vdd.n9823 0.01
R49352 vdd.n9877 vdd.n9809 0.01
R49353 vdd.n9877 vdd.n9815 0.01
R49354 vdd.n9878 vdd.n9801 0.01
R49355 vdd.n9878 vdd.n9807 0.01
R49356 vdd.n9879 vdd.n9793 0.01
R49357 vdd.n9879 vdd.n9799 0.01
R49358 vdd.n9880 vdd.n9785 0.01
R49359 vdd.n9880 vdd.n9789 0.01
R49360 vdd.n9881 vdd.n9777 0.01
R49361 vdd.n9881 vdd.n9783 0.01
R49362 vdd.n9882 vdd.n9769 0.01
R49363 vdd.n9882 vdd.n9775 0.01
R49364 vdd.n9883 vdd.n9761 0.01
R49365 vdd.n9883 vdd.n9767 0.01
R49366 vdd.n9884 vdd.n9753 0.01
R49367 vdd.n9884 vdd.n9759 0.01
R49368 vdd.n9885 vdd.n9745 0.01
R49369 vdd.n9885 vdd.n9751 0.01
R49370 vdd.n9886 vdd.n9737 0.01
R49371 vdd.n9886 vdd.n9743 0.01
R49372 vdd.n9887 vdd.n9729 0.01
R49373 vdd.n9887 vdd.n9735 0.01
R49374 vdd.n9888 vdd.n9721 0.01
R49375 vdd.n9888 vdd.n9727 0.01
R49376 vdd.n9899 vdd.n9894 0.01
R49377 vdd.n9899 vdd.n9895 0.01
R49378 vdd.n10050 vdd.n10048 0.01
R49379 vdd.n10050 vdd.n10044 0.01
R49380 vdd.n10051 vdd.n10037 0.01
R49381 vdd.n10051 vdd.n10043 0.01
R49382 vdd.n10052 vdd.n10029 0.01
R49383 vdd.n10052 vdd.n10035 0.01
R49384 vdd.n10053 vdd.n10021 0.01
R49385 vdd.n10053 vdd.n10027 0.01
R49386 vdd.n10054 vdd.n10013 0.01
R49387 vdd.n10054 vdd.n10019 0.01
R49388 vdd.n10055 vdd.n10005 0.01
R49389 vdd.n10055 vdd.n10011 0.01
R49390 vdd.n10056 vdd.n9997 0.01
R49391 vdd.n10056 vdd.n10003 0.01
R49392 vdd.n10057 vdd.n9989 0.01
R49393 vdd.n10057 vdd.n9995 0.01
R49394 vdd.n10058 vdd.n9981 0.01
R49395 vdd.n10058 vdd.n9987 0.01
R49396 vdd.n10059 vdd.n9973 0.01
R49397 vdd.n10059 vdd.n9979 0.01
R49398 vdd.n10060 vdd.n9965 0.01
R49399 vdd.n10060 vdd.n9969 0.01
R49400 vdd.n10061 vdd.n9957 0.01
R49401 vdd.n10061 vdd.n9963 0.01
R49402 vdd.n10062 vdd.n9949 0.01
R49403 vdd.n10062 vdd.n9955 0.01
R49404 vdd.n10063 vdd.n9941 0.01
R49405 vdd.n10063 vdd.n9947 0.01
R49406 vdd.n10064 vdd.n9933 0.01
R49407 vdd.n10064 vdd.n9939 0.01
R49408 vdd.n10065 vdd.n9925 0.01
R49409 vdd.n10065 vdd.n9931 0.01
R49410 vdd.n10066 vdd.n9917 0.01
R49411 vdd.n10066 vdd.n9923 0.01
R49412 vdd.n10067 vdd.n9909 0.01
R49413 vdd.n10067 vdd.n9915 0.01
R49414 vdd.n10068 vdd.n9901 0.01
R49415 vdd.n10068 vdd.n9907 0.01
R49416 vdd.n10079 vdd.n10074 0.01
R49417 vdd.n10079 vdd.n10075 0.01
R49418 vdd.n10230 vdd.n10228 0.01
R49419 vdd.n10230 vdd.n10224 0.01
R49420 vdd.n10231 vdd.n10217 0.01
R49421 vdd.n10231 vdd.n10223 0.01
R49422 vdd.n10232 vdd.n10209 0.01
R49423 vdd.n10232 vdd.n10215 0.01
R49424 vdd.n10233 vdd.n10201 0.01
R49425 vdd.n10233 vdd.n10207 0.01
R49426 vdd.n10234 vdd.n10193 0.01
R49427 vdd.n10234 vdd.n10199 0.01
R49428 vdd.n10235 vdd.n10185 0.01
R49429 vdd.n10235 vdd.n10191 0.01
R49430 vdd.n10236 vdd.n10177 0.01
R49431 vdd.n10236 vdd.n10183 0.01
R49432 vdd.n10237 vdd.n10169 0.01
R49433 vdd.n10237 vdd.n10175 0.01
R49434 vdd.n10238 vdd.n10161 0.01
R49435 vdd.n10238 vdd.n10167 0.01
R49436 vdd.n10239 vdd.n10153 0.01
R49437 vdd.n10239 vdd.n10159 0.01
R49438 vdd.n10240 vdd.n10145 0.01
R49439 vdd.n10240 vdd.n10149 0.01
R49440 vdd.n10241 vdd.n10137 0.01
R49441 vdd.n10241 vdd.n10143 0.01
R49442 vdd.n10242 vdd.n10129 0.01
R49443 vdd.n10242 vdd.n10135 0.01
R49444 vdd.n10243 vdd.n10121 0.01
R49445 vdd.n10243 vdd.n10127 0.01
R49446 vdd.n10244 vdd.n10113 0.01
R49447 vdd.n10244 vdd.n10119 0.01
R49448 vdd.n10245 vdd.n10105 0.01
R49449 vdd.n10245 vdd.n10111 0.01
R49450 vdd.n10246 vdd.n10097 0.01
R49451 vdd.n10246 vdd.n10103 0.01
R49452 vdd.n10247 vdd.n10089 0.01
R49453 vdd.n10247 vdd.n10095 0.01
R49454 vdd.n10248 vdd.n10081 0.01
R49455 vdd.n10248 vdd.n10087 0.01
R49456 vdd.n10259 vdd.n10254 0.01
R49457 vdd.n10259 vdd.n10255 0.01
R49458 vdd.n10410 vdd.n10408 0.01
R49459 vdd.n10410 vdd.n10404 0.01
R49460 vdd.n10411 vdd.n10397 0.01
R49461 vdd.n10411 vdd.n10403 0.01
R49462 vdd.n10412 vdd.n10389 0.01
R49463 vdd.n10412 vdd.n10395 0.01
R49464 vdd.n10413 vdd.n10381 0.01
R49465 vdd.n10413 vdd.n10387 0.01
R49466 vdd.n10414 vdd.n10373 0.01
R49467 vdd.n10414 vdd.n10379 0.01
R49468 vdd.n10415 vdd.n10365 0.01
R49469 vdd.n10415 vdd.n10371 0.01
R49470 vdd.n10416 vdd.n10357 0.01
R49471 vdd.n10416 vdd.n10363 0.01
R49472 vdd.n10417 vdd.n10349 0.01
R49473 vdd.n10417 vdd.n10355 0.01
R49474 vdd.n10418 vdd.n10341 0.01
R49475 vdd.n10418 vdd.n10347 0.01
R49476 vdd.n10419 vdd.n10333 0.01
R49477 vdd.n10419 vdd.n10339 0.01
R49478 vdd.n10420 vdd.n10325 0.01
R49479 vdd.n10420 vdd.n10329 0.01
R49480 vdd.n10421 vdd.n10317 0.01
R49481 vdd.n10421 vdd.n10323 0.01
R49482 vdd.n10422 vdd.n10309 0.01
R49483 vdd.n10422 vdd.n10315 0.01
R49484 vdd.n10423 vdd.n10301 0.01
R49485 vdd.n10423 vdd.n10307 0.01
R49486 vdd.n10424 vdd.n10293 0.01
R49487 vdd.n10424 vdd.n10299 0.01
R49488 vdd.n10425 vdd.n10285 0.01
R49489 vdd.n10425 vdd.n10291 0.01
R49490 vdd.n10426 vdd.n10277 0.01
R49491 vdd.n10426 vdd.n10283 0.01
R49492 vdd.n10427 vdd.n10269 0.01
R49493 vdd.n10427 vdd.n10275 0.01
R49494 vdd.n10428 vdd.n10261 0.01
R49495 vdd.n10428 vdd.n10267 0.01
R49496 vdd.n10439 vdd.n10434 0.01
R49497 vdd.n10439 vdd.n10435 0.01
R49498 vdd.n10590 vdd.n10588 0.01
R49499 vdd.n10590 vdd.n10584 0.01
R49500 vdd.n10591 vdd.n10577 0.01
R49501 vdd.n10591 vdd.n10583 0.01
R49502 vdd.n10592 vdd.n10569 0.01
R49503 vdd.n10592 vdd.n10575 0.01
R49504 vdd.n10593 vdd.n10561 0.01
R49505 vdd.n10593 vdd.n10567 0.01
R49506 vdd.n10594 vdd.n10553 0.01
R49507 vdd.n10594 vdd.n10559 0.01
R49508 vdd.n10595 vdd.n10545 0.01
R49509 vdd.n10595 vdd.n10551 0.01
R49510 vdd.n10596 vdd.n10537 0.01
R49511 vdd.n10596 vdd.n10543 0.01
R49512 vdd.n10597 vdd.n10529 0.01
R49513 vdd.n10597 vdd.n10535 0.01
R49514 vdd.n10598 vdd.n10521 0.01
R49515 vdd.n10598 vdd.n10527 0.01
R49516 vdd.n10599 vdd.n10513 0.01
R49517 vdd.n10599 vdd.n10519 0.01
R49518 vdd.n10600 vdd.n10505 0.01
R49519 vdd.n10600 vdd.n10509 0.01
R49520 vdd.n10601 vdd.n10497 0.01
R49521 vdd.n10601 vdd.n10503 0.01
R49522 vdd.n10602 vdd.n10489 0.01
R49523 vdd.n10602 vdd.n10495 0.01
R49524 vdd.n10603 vdd.n10481 0.01
R49525 vdd.n10603 vdd.n10487 0.01
R49526 vdd.n10604 vdd.n10473 0.01
R49527 vdd.n10604 vdd.n10479 0.01
R49528 vdd.n10605 vdd.n10465 0.01
R49529 vdd.n10605 vdd.n10471 0.01
R49530 vdd.n10606 vdd.n10457 0.01
R49531 vdd.n10606 vdd.n10463 0.01
R49532 vdd.n10607 vdd.n10449 0.01
R49533 vdd.n10607 vdd.n10455 0.01
R49534 vdd.n10608 vdd.n10441 0.01
R49535 vdd.n10608 vdd.n10447 0.01
R49536 vdd.n10619 vdd.n10614 0.01
R49537 vdd.n10619 vdd.n10615 0.01
R49538 vdd.n10770 vdd.n10768 0.01
R49539 vdd.n10770 vdd.n10764 0.01
R49540 vdd.n10771 vdd.n10757 0.01
R49541 vdd.n10771 vdd.n10763 0.01
R49542 vdd.n10772 vdd.n10749 0.01
R49543 vdd.n10772 vdd.n10755 0.01
R49544 vdd.n10773 vdd.n10741 0.01
R49545 vdd.n10773 vdd.n10747 0.01
R49546 vdd.n10774 vdd.n10733 0.01
R49547 vdd.n10774 vdd.n10739 0.01
R49548 vdd.n10775 vdd.n10725 0.01
R49549 vdd.n10775 vdd.n10731 0.01
R49550 vdd.n10776 vdd.n10717 0.01
R49551 vdd.n10776 vdd.n10723 0.01
R49552 vdd.n10777 vdd.n10709 0.01
R49553 vdd.n10777 vdd.n10715 0.01
R49554 vdd.n10778 vdd.n10701 0.01
R49555 vdd.n10778 vdd.n10707 0.01
R49556 vdd.n10779 vdd.n10693 0.01
R49557 vdd.n10779 vdd.n10699 0.01
R49558 vdd.n10780 vdd.n10685 0.01
R49559 vdd.n10780 vdd.n10689 0.01
R49560 vdd.n10781 vdd.n10677 0.01
R49561 vdd.n10781 vdd.n10683 0.01
R49562 vdd.n10782 vdd.n10669 0.01
R49563 vdd.n10782 vdd.n10675 0.01
R49564 vdd.n10783 vdd.n10661 0.01
R49565 vdd.n10783 vdd.n10667 0.01
R49566 vdd.n10784 vdd.n10653 0.01
R49567 vdd.n10784 vdd.n10659 0.01
R49568 vdd.n10785 vdd.n10645 0.01
R49569 vdd.n10785 vdd.n10651 0.01
R49570 vdd.n10786 vdd.n10637 0.01
R49571 vdd.n10786 vdd.n10643 0.01
R49572 vdd.n10787 vdd.n10629 0.01
R49573 vdd.n10787 vdd.n10635 0.01
R49574 vdd.n10788 vdd.n10621 0.01
R49575 vdd.n10788 vdd.n10627 0.01
R49576 vdd.n10799 vdd.n10794 0.01
R49577 vdd.n10799 vdd.n10795 0.01
R49578 vdd.n10950 vdd.n10948 0.01
R49579 vdd.n10950 vdd.n10944 0.01
R49580 vdd.n10951 vdd.n10937 0.01
R49581 vdd.n10951 vdd.n10943 0.01
R49582 vdd.n10952 vdd.n10929 0.01
R49583 vdd.n10952 vdd.n10935 0.01
R49584 vdd.n10953 vdd.n10921 0.01
R49585 vdd.n10953 vdd.n10927 0.01
R49586 vdd.n10954 vdd.n10913 0.01
R49587 vdd.n10954 vdd.n10919 0.01
R49588 vdd.n10955 vdd.n10905 0.01
R49589 vdd.n10955 vdd.n10911 0.01
R49590 vdd.n10956 vdd.n10897 0.01
R49591 vdd.n10956 vdd.n10903 0.01
R49592 vdd.n10957 vdd.n10889 0.01
R49593 vdd.n10957 vdd.n10895 0.01
R49594 vdd.n10958 vdd.n10881 0.01
R49595 vdd.n10958 vdd.n10887 0.01
R49596 vdd.n10959 vdd.n10873 0.01
R49597 vdd.n10959 vdd.n10879 0.01
R49598 vdd.n10960 vdd.n10865 0.01
R49599 vdd.n10960 vdd.n10869 0.01
R49600 vdd.n10961 vdd.n10857 0.01
R49601 vdd.n10961 vdd.n10863 0.01
R49602 vdd.n10962 vdd.n10849 0.01
R49603 vdd.n10962 vdd.n10855 0.01
R49604 vdd.n10963 vdd.n10841 0.01
R49605 vdd.n10963 vdd.n10847 0.01
R49606 vdd.n10964 vdd.n10833 0.01
R49607 vdd.n10964 vdd.n10839 0.01
R49608 vdd.n10965 vdd.n10825 0.01
R49609 vdd.n10965 vdd.n10831 0.01
R49610 vdd.n10966 vdd.n10817 0.01
R49611 vdd.n10966 vdd.n10823 0.01
R49612 vdd.n10967 vdd.n10809 0.01
R49613 vdd.n10967 vdd.n10815 0.01
R49614 vdd.n10968 vdd.n10801 0.01
R49615 vdd.n10968 vdd.n10807 0.01
R49616 vdd.n10979 vdd.n10974 0.01
R49617 vdd.n10979 vdd.n10975 0.01
R49618 vdd.n11130 vdd.n11128 0.01
R49619 vdd.n11130 vdd.n11124 0.01
R49620 vdd.n11131 vdd.n11117 0.01
R49621 vdd.n11131 vdd.n11123 0.01
R49622 vdd.n11132 vdd.n11109 0.01
R49623 vdd.n11132 vdd.n11115 0.01
R49624 vdd.n11133 vdd.n11101 0.01
R49625 vdd.n11133 vdd.n11107 0.01
R49626 vdd.n11134 vdd.n11093 0.01
R49627 vdd.n11134 vdd.n11099 0.01
R49628 vdd.n11135 vdd.n11085 0.01
R49629 vdd.n11135 vdd.n11091 0.01
R49630 vdd.n11136 vdd.n11077 0.01
R49631 vdd.n11136 vdd.n11083 0.01
R49632 vdd.n11137 vdd.n11069 0.01
R49633 vdd.n11137 vdd.n11075 0.01
R49634 vdd.n11138 vdd.n11061 0.01
R49635 vdd.n11138 vdd.n11067 0.01
R49636 vdd.n11139 vdd.n11053 0.01
R49637 vdd.n11139 vdd.n11059 0.01
R49638 vdd.n11140 vdd.n11045 0.01
R49639 vdd.n11140 vdd.n11049 0.01
R49640 vdd.n11141 vdd.n11037 0.01
R49641 vdd.n11141 vdd.n11043 0.01
R49642 vdd.n11142 vdd.n11029 0.01
R49643 vdd.n11142 vdd.n11035 0.01
R49644 vdd.n11143 vdd.n11021 0.01
R49645 vdd.n11143 vdd.n11027 0.01
R49646 vdd.n11144 vdd.n11013 0.01
R49647 vdd.n11144 vdd.n11019 0.01
R49648 vdd.n11145 vdd.n11005 0.01
R49649 vdd.n11145 vdd.n11011 0.01
R49650 vdd.n11146 vdd.n10997 0.01
R49651 vdd.n11146 vdd.n11003 0.01
R49652 vdd.n11147 vdd.n10989 0.01
R49653 vdd.n11147 vdd.n10995 0.01
R49654 vdd.n11148 vdd.n10981 0.01
R49655 vdd.n11148 vdd.n10987 0.01
R49656 vdd.n11159 vdd.n11154 0.01
R49657 vdd.n11159 vdd.n11155 0.01
R49658 vdd.n11310 vdd.n11308 0.01
R49659 vdd.n11310 vdd.n11304 0.01
R49660 vdd.n11311 vdd.n11297 0.01
R49661 vdd.n11311 vdd.n11303 0.01
R49662 vdd.n11312 vdd.n11289 0.01
R49663 vdd.n11312 vdd.n11295 0.01
R49664 vdd.n11313 vdd.n11281 0.01
R49665 vdd.n11313 vdd.n11287 0.01
R49666 vdd.n11314 vdd.n11273 0.01
R49667 vdd.n11314 vdd.n11279 0.01
R49668 vdd.n11315 vdd.n11265 0.01
R49669 vdd.n11315 vdd.n11271 0.01
R49670 vdd.n11316 vdd.n11257 0.01
R49671 vdd.n11316 vdd.n11263 0.01
R49672 vdd.n11317 vdd.n11249 0.01
R49673 vdd.n11317 vdd.n11255 0.01
R49674 vdd.n11318 vdd.n11241 0.01
R49675 vdd.n11318 vdd.n11247 0.01
R49676 vdd.n11319 vdd.n11233 0.01
R49677 vdd.n11319 vdd.n11239 0.01
R49678 vdd.n11320 vdd.n11225 0.01
R49679 vdd.n11320 vdd.n11229 0.01
R49680 vdd.n11321 vdd.n11217 0.01
R49681 vdd.n11321 vdd.n11223 0.01
R49682 vdd.n11322 vdd.n11209 0.01
R49683 vdd.n11322 vdd.n11215 0.01
R49684 vdd.n11323 vdd.n11201 0.01
R49685 vdd.n11323 vdd.n11207 0.01
R49686 vdd.n11324 vdd.n11193 0.01
R49687 vdd.n11324 vdd.n11199 0.01
R49688 vdd.n11325 vdd.n11185 0.01
R49689 vdd.n11325 vdd.n11191 0.01
R49690 vdd.n11326 vdd.n11177 0.01
R49691 vdd.n11326 vdd.n11183 0.01
R49692 vdd.n11327 vdd.n11169 0.01
R49693 vdd.n11327 vdd.n11175 0.01
R49694 vdd.n11328 vdd.n11161 0.01
R49695 vdd.n11328 vdd.n11167 0.01
R49696 vdd.n11339 vdd.n11334 0.01
R49697 vdd.n11339 vdd.n11335 0.01
R49698 vdd.n11362 vdd.n11361 0.01
R49699 vdd.n11365 vdd.n11364 0.01
R49700 vdd.n11368 vdd.n11367 0.01
R49701 vdd.n11371 vdd.n11370 0.01
R49702 vdd.n11374 vdd.n11373 0.01
R49703 vdd.n11377 vdd.n11376 0.01
R49704 vdd.n11380 vdd.n11379 0.01
R49705 vdd.n11383 vdd.n11382 0.01
R49706 vdd.n11390 vdd.n11389 0.01
R49707 vdd.n11393 vdd.n11392 0.01
R49708 vdd.n11396 vdd.n11395 0.01
R49709 vdd.n11399 vdd.n11398 0.01
R49710 vdd.n11402 vdd.n11401 0.01
R49711 vdd.n11405 vdd.n11404 0.01
R49712 vdd.n11408 vdd.n11407 0.01
R49713 vdd.n11411 vdd.n11410 0.01
R49714 vdd.n11417 vdd.n11416 0.003
R49715 vdd.n11418 vdd.n11417 0.003
R49716 vdd.n11419 vdd.n11418 0.003
R49717 vdd.n11420 vdd.n11419 0.003
R49718 vdd.n11421 vdd.n11420 0.003
R49719 vdd.n11422 vdd.n11421 0.003
R49720 vdd.n11423 vdd.n11422 0.003
R49721 vdd.n11424 vdd.n11423 0.003
R49722 vdd.n11425 vdd.n11424 0.003
R49723 vdd.n11426 vdd.n11425 0.003
R49724 vdd.n11427 vdd.n11426 0.003
R49725 vdd.n11428 vdd.n11427 0.003
R49726 vdd.n11429 vdd.n11428 0.003
R49727 vdd.n11430 vdd.n11429 0.003
R49728 vdd.n11431 vdd.n11430 0.003
R49729 vdd.n11432 vdd.n11431 0.003
R49730 vdd.n11433 vdd.n11432 0.003
R49731 vdd.n11434 vdd.n11433 0.003
R49732 vdd.n11435 vdd.n11434 0.003
R49733 vdd.n11436 vdd.n11435 0.003
R49734 vdd.n11437 vdd.n11436 0.003
R49735 vdd.n11438 vdd.n11437 0.003
R49736 vdd.n11439 vdd.n11438 0.003
R49737 vdd.n11440 vdd.n11439 0.003
R49738 vdd.n11441 vdd.n11440 0.003
R49739 vdd.n11442 vdd.n11441 0.003
R49740 vdd.n11443 vdd.n11442 0.003
R49741 vdd.n11444 vdd.n11443 0.003
R49742 vdd.n11445 vdd.n11444 0.003
R49743 vdd.n11446 vdd.n11445 0.003
R49744 vdd.n11447 vdd.n11446 0.003
R49745 vdd.n11448 vdd.n11447 0.003
R49746 vdd.n11449 vdd.n11448 0.003
R49747 vdd.n11450 vdd.n11449 0.003
R49748 vdd.n11451 vdd.n11450 0.003
R49749 vdd.n11452 vdd.n11451 0.003
R49750 vdd.n11453 vdd.n11452 0.003
R49751 vdd.n11454 vdd.n11453 0.003
R49752 vdd.n11455 vdd.n11454 0.003
R49753 vdd.n11456 vdd.n11455 0.003
R49754 vdd.n11457 vdd.n11456 0.003
R49755 vdd.n11458 vdd.n11457 0.003
R49756 vdd.n11459 vdd.n11458 0.003
R49757 vdd.n11460 vdd.n11459 0.003
R49758 vdd.n11461 vdd.n11460 0.003
R49759 vdd.n11462 vdd.n11461 0.003
R49760 vdd.n11463 vdd.n11462 0.003
R49761 vdd.n11464 vdd.n11463 0.003
R49762 vdd.n11465 vdd.n11464 0.003
R49763 vdd.n11466 vdd.n11465 0.003
R49764 vdd.n11467 vdd.n11466 0.003
R49765 vdd.n11468 vdd.n11467 0.003
R49766 vdd.n11469 vdd.n11468 0.003
R49767 vdd.n11470 vdd.n11469 0.003
R49768 vdd.n11471 vdd.n11470 0.003
R49769 vdd.n11472 vdd.n11471 0.003
R49770 vdd.n11473 vdd.n11472 0.003
R49771 vdd.n11474 vdd.n11473 0.003
R49772 vdd.n11475 vdd.n11474 0.003
R49773 vdd.n11476 vdd.n11475 0.003
R49774 vdd.n11477 vdd.n11476 0.003
R49775 vdd.n11478 vdd.n11477 0.003
R49776 vdd.n13545 vdd.n13544 0.003
R49777 vdd.n13544 vdd.n13543 0.003
R49778 vdd.n13543 vdd.n13542 0.003
R49779 vdd.n13542 vdd.n13541 0.003
R49780 vdd.n13541 vdd.n13540 0.003
R49781 vdd.n13540 vdd.n13539 0.003
R49782 vdd.n13539 vdd.n13538 0.003
R49783 vdd.n13538 vdd.n13537 0.003
R49784 vdd.n13537 vdd.n13536 0.003
R49785 vdd.n13536 vdd.n13535 0.003
R49786 vdd.n13418 vdd.n13417 0.002
R49787 vdd.n13420 vdd.n13419 0.002
R49788 vdd.n13410 vdd.n13409 0.002
R49789 vdd.n13412 vdd.n13411 0.002
R49790 vdd.n13402 vdd.n13401 0.002
R49791 vdd.n13404 vdd.n13403 0.002
R49792 vdd.n13394 vdd.n13393 0.002
R49793 vdd.n13396 vdd.n13395 0.002
R49794 vdd.n13386 vdd.n13385 0.002
R49795 vdd.n13388 vdd.n13387 0.002
R49796 vdd.n13378 vdd.n13377 0.002
R49797 vdd.n13380 vdd.n13379 0.002
R49798 vdd.n13370 vdd.n13369 0.002
R49799 vdd.n13372 vdd.n13371 0.002
R49800 vdd.n13362 vdd.n13361 0.002
R49801 vdd.n13364 vdd.n13363 0.002
R49802 vdd.n13354 vdd.n13353 0.002
R49803 vdd.n13356 vdd.n13355 0.002
R49804 vdd.n13338 vdd.n13337 0.002
R49805 vdd.n13340 vdd.n13339 0.002
R49806 vdd.n13330 vdd.n13329 0.002
R49807 vdd.n13332 vdd.n13331 0.002
R49808 vdd.n13322 vdd.n13321 0.002
R49809 vdd.n13324 vdd.n13323 0.002
R49810 vdd.n13314 vdd.n13313 0.002
R49811 vdd.n13316 vdd.n13315 0.002
R49812 vdd.n13306 vdd.n13305 0.002
R49813 vdd.n13308 vdd.n13307 0.002
R49814 vdd.n13298 vdd.n13297 0.002
R49815 vdd.n13300 vdd.n13299 0.002
R49816 vdd.n13290 vdd.n13289 0.002
R49817 vdd.n13292 vdd.n13291 0.002
R49818 vdd.n13282 vdd.n13281 0.002
R49819 vdd.n13284 vdd.n13283 0.002
R49820 vdd.n13449 vdd.n13448 0.002
R49821 vdd.n13451 vdd.n13450 0.002
R49822 vdd.n13238 vdd.n13237 0.002
R49823 vdd.n13240 vdd.n13239 0.002
R49824 vdd.n13230 vdd.n13229 0.002
R49825 vdd.n13232 vdd.n13231 0.002
R49826 vdd.n13222 vdd.n13221 0.002
R49827 vdd.n13224 vdd.n13223 0.002
R49828 vdd.n13214 vdd.n13213 0.002
R49829 vdd.n13216 vdd.n13215 0.002
R49830 vdd.n13206 vdd.n13205 0.002
R49831 vdd.n13208 vdd.n13207 0.002
R49832 vdd.n13198 vdd.n13197 0.002
R49833 vdd.n13200 vdd.n13199 0.002
R49834 vdd.n13190 vdd.n13189 0.002
R49835 vdd.n13192 vdd.n13191 0.002
R49836 vdd.n13182 vdd.n13181 0.002
R49837 vdd.n13184 vdd.n13183 0.002
R49838 vdd.n13174 vdd.n13173 0.002
R49839 vdd.n13176 vdd.n13175 0.002
R49840 vdd.n13158 vdd.n13157 0.002
R49841 vdd.n13160 vdd.n13159 0.002
R49842 vdd.n13150 vdd.n13149 0.002
R49843 vdd.n13152 vdd.n13151 0.002
R49844 vdd.n13142 vdd.n13141 0.002
R49845 vdd.n13144 vdd.n13143 0.002
R49846 vdd.n13134 vdd.n13133 0.002
R49847 vdd.n13136 vdd.n13135 0.002
R49848 vdd.n13126 vdd.n13125 0.002
R49849 vdd.n13128 vdd.n13127 0.002
R49850 vdd.n13118 vdd.n13117 0.002
R49851 vdd.n13120 vdd.n13119 0.002
R49852 vdd.n13110 vdd.n13109 0.002
R49853 vdd.n13112 vdd.n13111 0.002
R49854 vdd.n13102 vdd.n13101 0.002
R49855 vdd.n13104 vdd.n13103 0.002
R49856 vdd.n13269 vdd.n13268 0.002
R49857 vdd.n13271 vdd.n13270 0.002
R49858 vdd.n13058 vdd.n13057 0.002
R49859 vdd.n13060 vdd.n13059 0.002
R49860 vdd.n13050 vdd.n13049 0.002
R49861 vdd.n13052 vdd.n13051 0.002
R49862 vdd.n13042 vdd.n13041 0.002
R49863 vdd.n13044 vdd.n13043 0.002
R49864 vdd.n13034 vdd.n13033 0.002
R49865 vdd.n13036 vdd.n13035 0.002
R49866 vdd.n13026 vdd.n13025 0.002
R49867 vdd.n13028 vdd.n13027 0.002
R49868 vdd.n13018 vdd.n13017 0.002
R49869 vdd.n13020 vdd.n13019 0.002
R49870 vdd.n13010 vdd.n13009 0.002
R49871 vdd.n13012 vdd.n13011 0.002
R49872 vdd.n13002 vdd.n13001 0.002
R49873 vdd.n13004 vdd.n13003 0.002
R49874 vdd.n12994 vdd.n12993 0.002
R49875 vdd.n12996 vdd.n12995 0.002
R49876 vdd.n12978 vdd.n12977 0.002
R49877 vdd.n12980 vdd.n12979 0.002
R49878 vdd.n12970 vdd.n12969 0.002
R49879 vdd.n12972 vdd.n12971 0.002
R49880 vdd.n12962 vdd.n12961 0.002
R49881 vdd.n12964 vdd.n12963 0.002
R49882 vdd.n12954 vdd.n12953 0.002
R49883 vdd.n12956 vdd.n12955 0.002
R49884 vdd.n12946 vdd.n12945 0.002
R49885 vdd.n12948 vdd.n12947 0.002
R49886 vdd.n12938 vdd.n12937 0.002
R49887 vdd.n12940 vdd.n12939 0.002
R49888 vdd.n12930 vdd.n12929 0.002
R49889 vdd.n12932 vdd.n12931 0.002
R49890 vdd.n12922 vdd.n12921 0.002
R49891 vdd.n12924 vdd.n12923 0.002
R49892 vdd.n13089 vdd.n13088 0.002
R49893 vdd.n13091 vdd.n13090 0.002
R49894 vdd.n12878 vdd.n12877 0.002
R49895 vdd.n12880 vdd.n12879 0.002
R49896 vdd.n12870 vdd.n12869 0.002
R49897 vdd.n12872 vdd.n12871 0.002
R49898 vdd.n12862 vdd.n12861 0.002
R49899 vdd.n12864 vdd.n12863 0.002
R49900 vdd.n12854 vdd.n12853 0.002
R49901 vdd.n12856 vdd.n12855 0.002
R49902 vdd.n12846 vdd.n12845 0.002
R49903 vdd.n12848 vdd.n12847 0.002
R49904 vdd.n12838 vdd.n12837 0.002
R49905 vdd.n12840 vdd.n12839 0.002
R49906 vdd.n12830 vdd.n12829 0.002
R49907 vdd.n12832 vdd.n12831 0.002
R49908 vdd.n12822 vdd.n12821 0.002
R49909 vdd.n12824 vdd.n12823 0.002
R49910 vdd.n12814 vdd.n12813 0.002
R49911 vdd.n12816 vdd.n12815 0.002
R49912 vdd.n12798 vdd.n12797 0.002
R49913 vdd.n12800 vdd.n12799 0.002
R49914 vdd.n12790 vdd.n12789 0.002
R49915 vdd.n12792 vdd.n12791 0.002
R49916 vdd.n12782 vdd.n12781 0.002
R49917 vdd.n12784 vdd.n12783 0.002
R49918 vdd.n12774 vdd.n12773 0.002
R49919 vdd.n12776 vdd.n12775 0.002
R49920 vdd.n12766 vdd.n12765 0.002
R49921 vdd.n12768 vdd.n12767 0.002
R49922 vdd.n12758 vdd.n12757 0.002
R49923 vdd.n12760 vdd.n12759 0.002
R49924 vdd.n12750 vdd.n12749 0.002
R49925 vdd.n12752 vdd.n12751 0.002
R49926 vdd.n12742 vdd.n12741 0.002
R49927 vdd.n12744 vdd.n12743 0.002
R49928 vdd.n12909 vdd.n12908 0.002
R49929 vdd.n12911 vdd.n12910 0.002
R49930 vdd.n12698 vdd.n12697 0.002
R49931 vdd.n12700 vdd.n12699 0.002
R49932 vdd.n12690 vdd.n12689 0.002
R49933 vdd.n12692 vdd.n12691 0.002
R49934 vdd.n12682 vdd.n12681 0.002
R49935 vdd.n12684 vdd.n12683 0.002
R49936 vdd.n12674 vdd.n12673 0.002
R49937 vdd.n12676 vdd.n12675 0.002
R49938 vdd.n12666 vdd.n12665 0.002
R49939 vdd.n12668 vdd.n12667 0.002
R49940 vdd.n12658 vdd.n12657 0.002
R49941 vdd.n12660 vdd.n12659 0.002
R49942 vdd.n12650 vdd.n12649 0.002
R49943 vdd.n12652 vdd.n12651 0.002
R49944 vdd.n12642 vdd.n12641 0.002
R49945 vdd.n12644 vdd.n12643 0.002
R49946 vdd.n12634 vdd.n12633 0.002
R49947 vdd.n12636 vdd.n12635 0.002
R49948 vdd.n12618 vdd.n12617 0.002
R49949 vdd.n12620 vdd.n12619 0.002
R49950 vdd.n12610 vdd.n12609 0.002
R49951 vdd.n12612 vdd.n12611 0.002
R49952 vdd.n12602 vdd.n12601 0.002
R49953 vdd.n12604 vdd.n12603 0.002
R49954 vdd.n12594 vdd.n12593 0.002
R49955 vdd.n12596 vdd.n12595 0.002
R49956 vdd.n12586 vdd.n12585 0.002
R49957 vdd.n12588 vdd.n12587 0.002
R49958 vdd.n12578 vdd.n12577 0.002
R49959 vdd.n12580 vdd.n12579 0.002
R49960 vdd.n12570 vdd.n12569 0.002
R49961 vdd.n12572 vdd.n12571 0.002
R49962 vdd.n12562 vdd.n12561 0.002
R49963 vdd.n12564 vdd.n12563 0.002
R49964 vdd.n12729 vdd.n12728 0.002
R49965 vdd.n12731 vdd.n12730 0.002
R49966 vdd.n12518 vdd.n12517 0.002
R49967 vdd.n12520 vdd.n12519 0.002
R49968 vdd.n12510 vdd.n12509 0.002
R49969 vdd.n12512 vdd.n12511 0.002
R49970 vdd.n12502 vdd.n12501 0.002
R49971 vdd.n12504 vdd.n12503 0.002
R49972 vdd.n12494 vdd.n12493 0.002
R49973 vdd.n12496 vdd.n12495 0.002
R49974 vdd.n12486 vdd.n12485 0.002
R49975 vdd.n12488 vdd.n12487 0.002
R49976 vdd.n12478 vdd.n12477 0.002
R49977 vdd.n12480 vdd.n12479 0.002
R49978 vdd.n12470 vdd.n12469 0.002
R49979 vdd.n12472 vdd.n12471 0.002
R49980 vdd.n12462 vdd.n12461 0.002
R49981 vdd.n12464 vdd.n12463 0.002
R49982 vdd.n12454 vdd.n12453 0.002
R49983 vdd.n12456 vdd.n12455 0.002
R49984 vdd.n12438 vdd.n12437 0.002
R49985 vdd.n12440 vdd.n12439 0.002
R49986 vdd.n12430 vdd.n12429 0.002
R49987 vdd.n12432 vdd.n12431 0.002
R49988 vdd.n12422 vdd.n12421 0.002
R49989 vdd.n12424 vdd.n12423 0.002
R49990 vdd.n12414 vdd.n12413 0.002
R49991 vdd.n12416 vdd.n12415 0.002
R49992 vdd.n12406 vdd.n12405 0.002
R49993 vdd.n12408 vdd.n12407 0.002
R49994 vdd.n12398 vdd.n12397 0.002
R49995 vdd.n12400 vdd.n12399 0.002
R49996 vdd.n12390 vdd.n12389 0.002
R49997 vdd.n12392 vdd.n12391 0.002
R49998 vdd.n12382 vdd.n12381 0.002
R49999 vdd.n12384 vdd.n12383 0.002
R50000 vdd.n12549 vdd.n12548 0.002
R50001 vdd.n12551 vdd.n12550 0.002
R50002 vdd.n12338 vdd.n12337 0.002
R50003 vdd.n12340 vdd.n12339 0.002
R50004 vdd.n12330 vdd.n12329 0.002
R50005 vdd.n12332 vdd.n12331 0.002
R50006 vdd.n12322 vdd.n12321 0.002
R50007 vdd.n12324 vdd.n12323 0.002
R50008 vdd.n12314 vdd.n12313 0.002
R50009 vdd.n12316 vdd.n12315 0.002
R50010 vdd.n12306 vdd.n12305 0.002
R50011 vdd.n12308 vdd.n12307 0.002
R50012 vdd.n12298 vdd.n12297 0.002
R50013 vdd.n12300 vdd.n12299 0.002
R50014 vdd.n12290 vdd.n12289 0.002
R50015 vdd.n12292 vdd.n12291 0.002
R50016 vdd.n12282 vdd.n12281 0.002
R50017 vdd.n12284 vdd.n12283 0.002
R50018 vdd.n12274 vdd.n12273 0.002
R50019 vdd.n12276 vdd.n12275 0.002
R50020 vdd.n12258 vdd.n12257 0.002
R50021 vdd.n12260 vdd.n12259 0.002
R50022 vdd.n12250 vdd.n12249 0.002
R50023 vdd.n12252 vdd.n12251 0.002
R50024 vdd.n12242 vdd.n12241 0.002
R50025 vdd.n12244 vdd.n12243 0.002
R50026 vdd.n12234 vdd.n12233 0.002
R50027 vdd.n12236 vdd.n12235 0.002
R50028 vdd.n12226 vdd.n12225 0.002
R50029 vdd.n12228 vdd.n12227 0.002
R50030 vdd.n12218 vdd.n12217 0.002
R50031 vdd.n12220 vdd.n12219 0.002
R50032 vdd.n12210 vdd.n12209 0.002
R50033 vdd.n12212 vdd.n12211 0.002
R50034 vdd.n12202 vdd.n12201 0.002
R50035 vdd.n12204 vdd.n12203 0.002
R50036 vdd.n12369 vdd.n12368 0.002
R50037 vdd.n12371 vdd.n12370 0.002
R50038 vdd.n12158 vdd.n12157 0.002
R50039 vdd.n12160 vdd.n12159 0.002
R50040 vdd.n12150 vdd.n12149 0.002
R50041 vdd.n12152 vdd.n12151 0.002
R50042 vdd.n12142 vdd.n12141 0.002
R50043 vdd.n12144 vdd.n12143 0.002
R50044 vdd.n12134 vdd.n12133 0.002
R50045 vdd.n12136 vdd.n12135 0.002
R50046 vdd.n12126 vdd.n12125 0.002
R50047 vdd.n12128 vdd.n12127 0.002
R50048 vdd.n12118 vdd.n12117 0.002
R50049 vdd.n12120 vdd.n12119 0.002
R50050 vdd.n12110 vdd.n12109 0.002
R50051 vdd.n12112 vdd.n12111 0.002
R50052 vdd.n12102 vdd.n12101 0.002
R50053 vdd.n12104 vdd.n12103 0.002
R50054 vdd.n12094 vdd.n12093 0.002
R50055 vdd.n12096 vdd.n12095 0.002
R50056 vdd.n12078 vdd.n12077 0.002
R50057 vdd.n12080 vdd.n12079 0.002
R50058 vdd.n12070 vdd.n12069 0.002
R50059 vdd.n12072 vdd.n12071 0.002
R50060 vdd.n12062 vdd.n12061 0.002
R50061 vdd.n12064 vdd.n12063 0.002
R50062 vdd.n12054 vdd.n12053 0.002
R50063 vdd.n12056 vdd.n12055 0.002
R50064 vdd.n12046 vdd.n12045 0.002
R50065 vdd.n12048 vdd.n12047 0.002
R50066 vdd.n12038 vdd.n12037 0.002
R50067 vdd.n12040 vdd.n12039 0.002
R50068 vdd.n12030 vdd.n12029 0.002
R50069 vdd.n12032 vdd.n12031 0.002
R50070 vdd.n12022 vdd.n12021 0.002
R50071 vdd.n12024 vdd.n12023 0.002
R50072 vdd.n12189 vdd.n12188 0.002
R50073 vdd.n12191 vdd.n12190 0.002
R50074 vdd.n11978 vdd.n11977 0.002
R50075 vdd.n11980 vdd.n11979 0.002
R50076 vdd.n11970 vdd.n11969 0.002
R50077 vdd.n11972 vdd.n11971 0.002
R50078 vdd.n11962 vdd.n11961 0.002
R50079 vdd.n11964 vdd.n11963 0.002
R50080 vdd.n11954 vdd.n11953 0.002
R50081 vdd.n11956 vdd.n11955 0.002
R50082 vdd.n11946 vdd.n11945 0.002
R50083 vdd.n11948 vdd.n11947 0.002
R50084 vdd.n11938 vdd.n11937 0.002
R50085 vdd.n11940 vdd.n11939 0.002
R50086 vdd.n11930 vdd.n11929 0.002
R50087 vdd.n11932 vdd.n11931 0.002
R50088 vdd.n11922 vdd.n11921 0.002
R50089 vdd.n11924 vdd.n11923 0.002
R50090 vdd.n11914 vdd.n11913 0.002
R50091 vdd.n11916 vdd.n11915 0.002
R50092 vdd.n11898 vdd.n11897 0.002
R50093 vdd.n11900 vdd.n11899 0.002
R50094 vdd.n11890 vdd.n11889 0.002
R50095 vdd.n11892 vdd.n11891 0.002
R50096 vdd.n11882 vdd.n11881 0.002
R50097 vdd.n11884 vdd.n11883 0.002
R50098 vdd.n11874 vdd.n11873 0.002
R50099 vdd.n11876 vdd.n11875 0.002
R50100 vdd.n11866 vdd.n11865 0.002
R50101 vdd.n11868 vdd.n11867 0.002
R50102 vdd.n11858 vdd.n11857 0.002
R50103 vdd.n11860 vdd.n11859 0.002
R50104 vdd.n11850 vdd.n11849 0.002
R50105 vdd.n11852 vdd.n11851 0.002
R50106 vdd.n11842 vdd.n11841 0.002
R50107 vdd.n11844 vdd.n11843 0.002
R50108 vdd.n12009 vdd.n12008 0.002
R50109 vdd.n12011 vdd.n12010 0.002
R50110 vdd.n11798 vdd.n11797 0.002
R50111 vdd.n11800 vdd.n11799 0.002
R50112 vdd.n11790 vdd.n11789 0.002
R50113 vdd.n11792 vdd.n11791 0.002
R50114 vdd.n11782 vdd.n11781 0.002
R50115 vdd.n11784 vdd.n11783 0.002
R50116 vdd.n11774 vdd.n11773 0.002
R50117 vdd.n11776 vdd.n11775 0.002
R50118 vdd.n11766 vdd.n11765 0.002
R50119 vdd.n11768 vdd.n11767 0.002
R50120 vdd.n11758 vdd.n11757 0.002
R50121 vdd.n11760 vdd.n11759 0.002
R50122 vdd.n11750 vdd.n11749 0.002
R50123 vdd.n11752 vdd.n11751 0.002
R50124 vdd.n11742 vdd.n11741 0.002
R50125 vdd.n11744 vdd.n11743 0.002
R50126 vdd.n11734 vdd.n11733 0.002
R50127 vdd.n11736 vdd.n11735 0.002
R50128 vdd.n11718 vdd.n11717 0.002
R50129 vdd.n11720 vdd.n11719 0.002
R50130 vdd.n11710 vdd.n11709 0.002
R50131 vdd.n11712 vdd.n11711 0.002
R50132 vdd.n11702 vdd.n11701 0.002
R50133 vdd.n11704 vdd.n11703 0.002
R50134 vdd.n11694 vdd.n11693 0.002
R50135 vdd.n11696 vdd.n11695 0.002
R50136 vdd.n11686 vdd.n11685 0.002
R50137 vdd.n11688 vdd.n11687 0.002
R50138 vdd.n11678 vdd.n11677 0.002
R50139 vdd.n11680 vdd.n11679 0.002
R50140 vdd.n11670 vdd.n11669 0.002
R50141 vdd.n11672 vdd.n11671 0.002
R50142 vdd.n11662 vdd.n11661 0.002
R50143 vdd.n11664 vdd.n11663 0.002
R50144 vdd.n11829 vdd.n11828 0.002
R50145 vdd.n11831 vdd.n11830 0.002
R50146 vdd.n11618 vdd.n11617 0.002
R50147 vdd.n11620 vdd.n11619 0.002
R50148 vdd.n11610 vdd.n11609 0.002
R50149 vdd.n11612 vdd.n11611 0.002
R50150 vdd.n11602 vdd.n11601 0.002
R50151 vdd.n11604 vdd.n11603 0.002
R50152 vdd.n11594 vdd.n11593 0.002
R50153 vdd.n11596 vdd.n11595 0.002
R50154 vdd.n11586 vdd.n11585 0.002
R50155 vdd.n11588 vdd.n11587 0.002
R50156 vdd.n11578 vdd.n11577 0.002
R50157 vdd.n11580 vdd.n11579 0.002
R50158 vdd.n11570 vdd.n11569 0.002
R50159 vdd.n11572 vdd.n11571 0.002
R50160 vdd.n11562 vdd.n11561 0.002
R50161 vdd.n11564 vdd.n11563 0.002
R50162 vdd.n11554 vdd.n11553 0.002
R50163 vdd.n11556 vdd.n11555 0.002
R50164 vdd.n11538 vdd.n11537 0.002
R50165 vdd.n11540 vdd.n11539 0.002
R50166 vdd.n11530 vdd.n11529 0.002
R50167 vdd.n11532 vdd.n11531 0.002
R50168 vdd.n11522 vdd.n11521 0.002
R50169 vdd.n11524 vdd.n11523 0.002
R50170 vdd.n11514 vdd.n11513 0.002
R50171 vdd.n11516 vdd.n11515 0.002
R50172 vdd.n11506 vdd.n11505 0.002
R50173 vdd.n11508 vdd.n11507 0.002
R50174 vdd.n11498 vdd.n11497 0.002
R50175 vdd.n11500 vdd.n11499 0.002
R50176 vdd.n11490 vdd.n11489 0.002
R50177 vdd.n11492 vdd.n11491 0.002
R50178 vdd.n11482 vdd.n11481 0.002
R50179 vdd.n11484 vdd.n11483 0.002
R50180 vdd.n11649 vdd.n11648 0.002
R50181 vdd.n11651 vdd.n11650 0.002
R50182 vdd.n139 vdd.n138 0.002
R50183 vdd.n141 vdd.n140 0.002
R50184 vdd.n131 vdd.n130 0.002
R50185 vdd.n133 vdd.n132 0.002
R50186 vdd.n123 vdd.n122 0.002
R50187 vdd.n125 vdd.n124 0.002
R50188 vdd.n115 vdd.n114 0.002
R50189 vdd.n117 vdd.n116 0.002
R50190 vdd.n107 vdd.n106 0.002
R50191 vdd.n109 vdd.n108 0.002
R50192 vdd.n99 vdd.n98 0.002
R50193 vdd.n101 vdd.n100 0.002
R50194 vdd.n91 vdd.n90 0.002
R50195 vdd.n93 vdd.n92 0.002
R50196 vdd.n83 vdd.n82 0.002
R50197 vdd.n85 vdd.n84 0.002
R50198 vdd.n75 vdd.n74 0.002
R50199 vdd.n77 vdd.n76 0.002
R50200 vdd.n59 vdd.n58 0.002
R50201 vdd.n61 vdd.n60 0.002
R50202 vdd.n51 vdd.n50 0.002
R50203 vdd.n53 vdd.n52 0.002
R50204 vdd.n43 vdd.n42 0.002
R50205 vdd.n45 vdd.n44 0.002
R50206 vdd.n35 vdd.n34 0.002
R50207 vdd.n37 vdd.n36 0.002
R50208 vdd.n27 vdd.n26 0.002
R50209 vdd.n29 vdd.n28 0.002
R50210 vdd.n19 vdd.n18 0.002
R50211 vdd.n21 vdd.n20 0.002
R50212 vdd.n11 vdd.n10 0.002
R50213 vdd.n13 vdd.n12 0.002
R50214 vdd.n3 vdd.n2 0.002
R50215 vdd.n5 vdd.n4 0.002
R50216 vdd.n170 vdd.n169 0.002
R50217 vdd.n172 vdd.n171 0.002
R50218 vdd.n319 vdd.n318 0.002
R50219 vdd.n321 vdd.n320 0.002
R50220 vdd.n311 vdd.n310 0.002
R50221 vdd.n313 vdd.n312 0.002
R50222 vdd.n303 vdd.n302 0.002
R50223 vdd.n305 vdd.n304 0.002
R50224 vdd.n295 vdd.n294 0.002
R50225 vdd.n297 vdd.n296 0.002
R50226 vdd.n287 vdd.n286 0.002
R50227 vdd.n289 vdd.n288 0.002
R50228 vdd.n279 vdd.n278 0.002
R50229 vdd.n281 vdd.n280 0.002
R50230 vdd.n271 vdd.n270 0.002
R50231 vdd.n273 vdd.n272 0.002
R50232 vdd.n263 vdd.n262 0.002
R50233 vdd.n265 vdd.n264 0.002
R50234 vdd.n255 vdd.n254 0.002
R50235 vdd.n257 vdd.n256 0.002
R50236 vdd.n239 vdd.n238 0.002
R50237 vdd.n241 vdd.n240 0.002
R50238 vdd.n231 vdd.n230 0.002
R50239 vdd.n233 vdd.n232 0.002
R50240 vdd.n223 vdd.n222 0.002
R50241 vdd.n225 vdd.n224 0.002
R50242 vdd.n215 vdd.n214 0.002
R50243 vdd.n217 vdd.n216 0.002
R50244 vdd.n207 vdd.n206 0.002
R50245 vdd.n209 vdd.n208 0.002
R50246 vdd.n199 vdd.n198 0.002
R50247 vdd.n201 vdd.n200 0.002
R50248 vdd.n191 vdd.n190 0.002
R50249 vdd.n193 vdd.n192 0.002
R50250 vdd.n183 vdd.n182 0.002
R50251 vdd.n185 vdd.n184 0.002
R50252 vdd.n350 vdd.n349 0.002
R50253 vdd.n352 vdd.n351 0.002
R50254 vdd.n499 vdd.n498 0.002
R50255 vdd.n501 vdd.n500 0.002
R50256 vdd.n491 vdd.n490 0.002
R50257 vdd.n493 vdd.n492 0.002
R50258 vdd.n483 vdd.n482 0.002
R50259 vdd.n485 vdd.n484 0.002
R50260 vdd.n475 vdd.n474 0.002
R50261 vdd.n477 vdd.n476 0.002
R50262 vdd.n467 vdd.n466 0.002
R50263 vdd.n469 vdd.n468 0.002
R50264 vdd.n459 vdd.n458 0.002
R50265 vdd.n461 vdd.n460 0.002
R50266 vdd.n451 vdd.n450 0.002
R50267 vdd.n453 vdd.n452 0.002
R50268 vdd.n443 vdd.n442 0.002
R50269 vdd.n445 vdd.n444 0.002
R50270 vdd.n435 vdd.n434 0.002
R50271 vdd.n437 vdd.n436 0.002
R50272 vdd.n419 vdd.n418 0.002
R50273 vdd.n421 vdd.n420 0.002
R50274 vdd.n411 vdd.n410 0.002
R50275 vdd.n413 vdd.n412 0.002
R50276 vdd.n403 vdd.n402 0.002
R50277 vdd.n405 vdd.n404 0.002
R50278 vdd.n395 vdd.n394 0.002
R50279 vdd.n397 vdd.n396 0.002
R50280 vdd.n387 vdd.n386 0.002
R50281 vdd.n389 vdd.n388 0.002
R50282 vdd.n379 vdd.n378 0.002
R50283 vdd.n381 vdd.n380 0.002
R50284 vdd.n371 vdd.n370 0.002
R50285 vdd.n373 vdd.n372 0.002
R50286 vdd.n363 vdd.n362 0.002
R50287 vdd.n365 vdd.n364 0.002
R50288 vdd.n530 vdd.n529 0.002
R50289 vdd.n532 vdd.n531 0.002
R50290 vdd.n679 vdd.n678 0.002
R50291 vdd.n681 vdd.n680 0.002
R50292 vdd.n671 vdd.n670 0.002
R50293 vdd.n673 vdd.n672 0.002
R50294 vdd.n663 vdd.n662 0.002
R50295 vdd.n665 vdd.n664 0.002
R50296 vdd.n655 vdd.n654 0.002
R50297 vdd.n657 vdd.n656 0.002
R50298 vdd.n647 vdd.n646 0.002
R50299 vdd.n649 vdd.n648 0.002
R50300 vdd.n639 vdd.n638 0.002
R50301 vdd.n641 vdd.n640 0.002
R50302 vdd.n631 vdd.n630 0.002
R50303 vdd.n633 vdd.n632 0.002
R50304 vdd.n623 vdd.n622 0.002
R50305 vdd.n625 vdd.n624 0.002
R50306 vdd.n615 vdd.n614 0.002
R50307 vdd.n617 vdd.n616 0.002
R50308 vdd.n599 vdd.n598 0.002
R50309 vdd.n601 vdd.n600 0.002
R50310 vdd.n591 vdd.n590 0.002
R50311 vdd.n593 vdd.n592 0.002
R50312 vdd.n583 vdd.n582 0.002
R50313 vdd.n585 vdd.n584 0.002
R50314 vdd.n575 vdd.n574 0.002
R50315 vdd.n577 vdd.n576 0.002
R50316 vdd.n567 vdd.n566 0.002
R50317 vdd.n569 vdd.n568 0.002
R50318 vdd.n559 vdd.n558 0.002
R50319 vdd.n561 vdd.n560 0.002
R50320 vdd.n551 vdd.n550 0.002
R50321 vdd.n553 vdd.n552 0.002
R50322 vdd.n543 vdd.n542 0.002
R50323 vdd.n545 vdd.n544 0.002
R50324 vdd.n710 vdd.n709 0.002
R50325 vdd.n712 vdd.n711 0.002
R50326 vdd.n859 vdd.n858 0.002
R50327 vdd.n861 vdd.n860 0.002
R50328 vdd.n851 vdd.n850 0.002
R50329 vdd.n853 vdd.n852 0.002
R50330 vdd.n843 vdd.n842 0.002
R50331 vdd.n845 vdd.n844 0.002
R50332 vdd.n835 vdd.n834 0.002
R50333 vdd.n837 vdd.n836 0.002
R50334 vdd.n827 vdd.n826 0.002
R50335 vdd.n829 vdd.n828 0.002
R50336 vdd.n819 vdd.n818 0.002
R50337 vdd.n821 vdd.n820 0.002
R50338 vdd.n811 vdd.n810 0.002
R50339 vdd.n813 vdd.n812 0.002
R50340 vdd.n803 vdd.n802 0.002
R50341 vdd.n805 vdd.n804 0.002
R50342 vdd.n795 vdd.n794 0.002
R50343 vdd.n797 vdd.n796 0.002
R50344 vdd.n779 vdd.n778 0.002
R50345 vdd.n781 vdd.n780 0.002
R50346 vdd.n771 vdd.n770 0.002
R50347 vdd.n773 vdd.n772 0.002
R50348 vdd.n763 vdd.n762 0.002
R50349 vdd.n765 vdd.n764 0.002
R50350 vdd.n755 vdd.n754 0.002
R50351 vdd.n757 vdd.n756 0.002
R50352 vdd.n747 vdd.n746 0.002
R50353 vdd.n749 vdd.n748 0.002
R50354 vdd.n739 vdd.n738 0.002
R50355 vdd.n741 vdd.n740 0.002
R50356 vdd.n731 vdd.n730 0.002
R50357 vdd.n733 vdd.n732 0.002
R50358 vdd.n723 vdd.n722 0.002
R50359 vdd.n725 vdd.n724 0.002
R50360 vdd.n890 vdd.n889 0.002
R50361 vdd.n892 vdd.n891 0.002
R50362 vdd.n1039 vdd.n1038 0.002
R50363 vdd.n1041 vdd.n1040 0.002
R50364 vdd.n1031 vdd.n1030 0.002
R50365 vdd.n1033 vdd.n1032 0.002
R50366 vdd.n1023 vdd.n1022 0.002
R50367 vdd.n1025 vdd.n1024 0.002
R50368 vdd.n1015 vdd.n1014 0.002
R50369 vdd.n1017 vdd.n1016 0.002
R50370 vdd.n1007 vdd.n1006 0.002
R50371 vdd.n1009 vdd.n1008 0.002
R50372 vdd.n999 vdd.n998 0.002
R50373 vdd.n1001 vdd.n1000 0.002
R50374 vdd.n991 vdd.n990 0.002
R50375 vdd.n993 vdd.n992 0.002
R50376 vdd.n983 vdd.n982 0.002
R50377 vdd.n985 vdd.n984 0.002
R50378 vdd.n975 vdd.n974 0.002
R50379 vdd.n977 vdd.n976 0.002
R50380 vdd.n959 vdd.n958 0.002
R50381 vdd.n961 vdd.n960 0.002
R50382 vdd.n951 vdd.n950 0.002
R50383 vdd.n953 vdd.n952 0.002
R50384 vdd.n943 vdd.n942 0.002
R50385 vdd.n945 vdd.n944 0.002
R50386 vdd.n935 vdd.n934 0.002
R50387 vdd.n937 vdd.n936 0.002
R50388 vdd.n927 vdd.n926 0.002
R50389 vdd.n929 vdd.n928 0.002
R50390 vdd.n919 vdd.n918 0.002
R50391 vdd.n921 vdd.n920 0.002
R50392 vdd.n911 vdd.n910 0.002
R50393 vdd.n913 vdd.n912 0.002
R50394 vdd.n903 vdd.n902 0.002
R50395 vdd.n905 vdd.n904 0.002
R50396 vdd.n1070 vdd.n1069 0.002
R50397 vdd.n1072 vdd.n1071 0.002
R50398 vdd.n1219 vdd.n1218 0.002
R50399 vdd.n1221 vdd.n1220 0.002
R50400 vdd.n1211 vdd.n1210 0.002
R50401 vdd.n1213 vdd.n1212 0.002
R50402 vdd.n1203 vdd.n1202 0.002
R50403 vdd.n1205 vdd.n1204 0.002
R50404 vdd.n1195 vdd.n1194 0.002
R50405 vdd.n1197 vdd.n1196 0.002
R50406 vdd.n1187 vdd.n1186 0.002
R50407 vdd.n1189 vdd.n1188 0.002
R50408 vdd.n1179 vdd.n1178 0.002
R50409 vdd.n1181 vdd.n1180 0.002
R50410 vdd.n1171 vdd.n1170 0.002
R50411 vdd.n1173 vdd.n1172 0.002
R50412 vdd.n1163 vdd.n1162 0.002
R50413 vdd.n1165 vdd.n1164 0.002
R50414 vdd.n1155 vdd.n1154 0.002
R50415 vdd.n1157 vdd.n1156 0.002
R50416 vdd.n1139 vdd.n1138 0.002
R50417 vdd.n1141 vdd.n1140 0.002
R50418 vdd.n1131 vdd.n1130 0.002
R50419 vdd.n1133 vdd.n1132 0.002
R50420 vdd.n1123 vdd.n1122 0.002
R50421 vdd.n1125 vdd.n1124 0.002
R50422 vdd.n1115 vdd.n1114 0.002
R50423 vdd.n1117 vdd.n1116 0.002
R50424 vdd.n1107 vdd.n1106 0.002
R50425 vdd.n1109 vdd.n1108 0.002
R50426 vdd.n1099 vdd.n1098 0.002
R50427 vdd.n1101 vdd.n1100 0.002
R50428 vdd.n1091 vdd.n1090 0.002
R50429 vdd.n1093 vdd.n1092 0.002
R50430 vdd.n1083 vdd.n1082 0.002
R50431 vdd.n1085 vdd.n1084 0.002
R50432 vdd.n1250 vdd.n1249 0.002
R50433 vdd.n1252 vdd.n1251 0.002
R50434 vdd.n1399 vdd.n1398 0.002
R50435 vdd.n1401 vdd.n1400 0.002
R50436 vdd.n1391 vdd.n1390 0.002
R50437 vdd.n1393 vdd.n1392 0.002
R50438 vdd.n1383 vdd.n1382 0.002
R50439 vdd.n1385 vdd.n1384 0.002
R50440 vdd.n1375 vdd.n1374 0.002
R50441 vdd.n1377 vdd.n1376 0.002
R50442 vdd.n1367 vdd.n1366 0.002
R50443 vdd.n1369 vdd.n1368 0.002
R50444 vdd.n1359 vdd.n1358 0.002
R50445 vdd.n1361 vdd.n1360 0.002
R50446 vdd.n1351 vdd.n1350 0.002
R50447 vdd.n1353 vdd.n1352 0.002
R50448 vdd.n1343 vdd.n1342 0.002
R50449 vdd.n1345 vdd.n1344 0.002
R50450 vdd.n1335 vdd.n1334 0.002
R50451 vdd.n1337 vdd.n1336 0.002
R50452 vdd.n1319 vdd.n1318 0.002
R50453 vdd.n1321 vdd.n1320 0.002
R50454 vdd.n1311 vdd.n1310 0.002
R50455 vdd.n1313 vdd.n1312 0.002
R50456 vdd.n1303 vdd.n1302 0.002
R50457 vdd.n1305 vdd.n1304 0.002
R50458 vdd.n1295 vdd.n1294 0.002
R50459 vdd.n1297 vdd.n1296 0.002
R50460 vdd.n1287 vdd.n1286 0.002
R50461 vdd.n1289 vdd.n1288 0.002
R50462 vdd.n1279 vdd.n1278 0.002
R50463 vdd.n1281 vdd.n1280 0.002
R50464 vdd.n1271 vdd.n1270 0.002
R50465 vdd.n1273 vdd.n1272 0.002
R50466 vdd.n1263 vdd.n1262 0.002
R50467 vdd.n1265 vdd.n1264 0.002
R50468 vdd.n1430 vdd.n1429 0.002
R50469 vdd.n1432 vdd.n1431 0.002
R50470 vdd.n1579 vdd.n1578 0.002
R50471 vdd.n1581 vdd.n1580 0.002
R50472 vdd.n1571 vdd.n1570 0.002
R50473 vdd.n1573 vdd.n1572 0.002
R50474 vdd.n1563 vdd.n1562 0.002
R50475 vdd.n1565 vdd.n1564 0.002
R50476 vdd.n1555 vdd.n1554 0.002
R50477 vdd.n1557 vdd.n1556 0.002
R50478 vdd.n1547 vdd.n1546 0.002
R50479 vdd.n1549 vdd.n1548 0.002
R50480 vdd.n1539 vdd.n1538 0.002
R50481 vdd.n1541 vdd.n1540 0.002
R50482 vdd.n1531 vdd.n1530 0.002
R50483 vdd.n1533 vdd.n1532 0.002
R50484 vdd.n1523 vdd.n1522 0.002
R50485 vdd.n1525 vdd.n1524 0.002
R50486 vdd.n1515 vdd.n1514 0.002
R50487 vdd.n1517 vdd.n1516 0.002
R50488 vdd.n1499 vdd.n1498 0.002
R50489 vdd.n1501 vdd.n1500 0.002
R50490 vdd.n1491 vdd.n1490 0.002
R50491 vdd.n1493 vdd.n1492 0.002
R50492 vdd.n1483 vdd.n1482 0.002
R50493 vdd.n1485 vdd.n1484 0.002
R50494 vdd.n1475 vdd.n1474 0.002
R50495 vdd.n1477 vdd.n1476 0.002
R50496 vdd.n1467 vdd.n1466 0.002
R50497 vdd.n1469 vdd.n1468 0.002
R50498 vdd.n1459 vdd.n1458 0.002
R50499 vdd.n1461 vdd.n1460 0.002
R50500 vdd.n1451 vdd.n1450 0.002
R50501 vdd.n1453 vdd.n1452 0.002
R50502 vdd.n1443 vdd.n1442 0.002
R50503 vdd.n1445 vdd.n1444 0.002
R50504 vdd.n1610 vdd.n1609 0.002
R50505 vdd.n1612 vdd.n1611 0.002
R50506 vdd.n1759 vdd.n1758 0.002
R50507 vdd.n1761 vdd.n1760 0.002
R50508 vdd.n1751 vdd.n1750 0.002
R50509 vdd.n1753 vdd.n1752 0.002
R50510 vdd.n1743 vdd.n1742 0.002
R50511 vdd.n1745 vdd.n1744 0.002
R50512 vdd.n1735 vdd.n1734 0.002
R50513 vdd.n1737 vdd.n1736 0.002
R50514 vdd.n1727 vdd.n1726 0.002
R50515 vdd.n1729 vdd.n1728 0.002
R50516 vdd.n1719 vdd.n1718 0.002
R50517 vdd.n1721 vdd.n1720 0.002
R50518 vdd.n1711 vdd.n1710 0.002
R50519 vdd.n1713 vdd.n1712 0.002
R50520 vdd.n1703 vdd.n1702 0.002
R50521 vdd.n1705 vdd.n1704 0.002
R50522 vdd.n1695 vdd.n1694 0.002
R50523 vdd.n1697 vdd.n1696 0.002
R50524 vdd.n1679 vdd.n1678 0.002
R50525 vdd.n1681 vdd.n1680 0.002
R50526 vdd.n1671 vdd.n1670 0.002
R50527 vdd.n1673 vdd.n1672 0.002
R50528 vdd.n1663 vdd.n1662 0.002
R50529 vdd.n1665 vdd.n1664 0.002
R50530 vdd.n1655 vdd.n1654 0.002
R50531 vdd.n1657 vdd.n1656 0.002
R50532 vdd.n1647 vdd.n1646 0.002
R50533 vdd.n1649 vdd.n1648 0.002
R50534 vdd.n1639 vdd.n1638 0.002
R50535 vdd.n1641 vdd.n1640 0.002
R50536 vdd.n1631 vdd.n1630 0.002
R50537 vdd.n1633 vdd.n1632 0.002
R50538 vdd.n1623 vdd.n1622 0.002
R50539 vdd.n1625 vdd.n1624 0.002
R50540 vdd.n1790 vdd.n1789 0.002
R50541 vdd.n1792 vdd.n1791 0.002
R50542 vdd.n1939 vdd.n1938 0.002
R50543 vdd.n1941 vdd.n1940 0.002
R50544 vdd.n1931 vdd.n1930 0.002
R50545 vdd.n1933 vdd.n1932 0.002
R50546 vdd.n1923 vdd.n1922 0.002
R50547 vdd.n1925 vdd.n1924 0.002
R50548 vdd.n1915 vdd.n1914 0.002
R50549 vdd.n1917 vdd.n1916 0.002
R50550 vdd.n1907 vdd.n1906 0.002
R50551 vdd.n1909 vdd.n1908 0.002
R50552 vdd.n1899 vdd.n1898 0.002
R50553 vdd.n1901 vdd.n1900 0.002
R50554 vdd.n1891 vdd.n1890 0.002
R50555 vdd.n1893 vdd.n1892 0.002
R50556 vdd.n1883 vdd.n1882 0.002
R50557 vdd.n1885 vdd.n1884 0.002
R50558 vdd.n1875 vdd.n1874 0.002
R50559 vdd.n1877 vdd.n1876 0.002
R50560 vdd.n1859 vdd.n1858 0.002
R50561 vdd.n1861 vdd.n1860 0.002
R50562 vdd.n1851 vdd.n1850 0.002
R50563 vdd.n1853 vdd.n1852 0.002
R50564 vdd.n1843 vdd.n1842 0.002
R50565 vdd.n1845 vdd.n1844 0.002
R50566 vdd.n1835 vdd.n1834 0.002
R50567 vdd.n1837 vdd.n1836 0.002
R50568 vdd.n1827 vdd.n1826 0.002
R50569 vdd.n1829 vdd.n1828 0.002
R50570 vdd.n1819 vdd.n1818 0.002
R50571 vdd.n1821 vdd.n1820 0.002
R50572 vdd.n1811 vdd.n1810 0.002
R50573 vdd.n1813 vdd.n1812 0.002
R50574 vdd.n1803 vdd.n1802 0.002
R50575 vdd.n1805 vdd.n1804 0.002
R50576 vdd.n1970 vdd.n1969 0.002
R50577 vdd.n1972 vdd.n1971 0.002
R50578 vdd.n2119 vdd.n2118 0.002
R50579 vdd.n2121 vdd.n2120 0.002
R50580 vdd.n2111 vdd.n2110 0.002
R50581 vdd.n2113 vdd.n2112 0.002
R50582 vdd.n2103 vdd.n2102 0.002
R50583 vdd.n2105 vdd.n2104 0.002
R50584 vdd.n2095 vdd.n2094 0.002
R50585 vdd.n2097 vdd.n2096 0.002
R50586 vdd.n2087 vdd.n2086 0.002
R50587 vdd.n2089 vdd.n2088 0.002
R50588 vdd.n2079 vdd.n2078 0.002
R50589 vdd.n2081 vdd.n2080 0.002
R50590 vdd.n2071 vdd.n2070 0.002
R50591 vdd.n2073 vdd.n2072 0.002
R50592 vdd.n2063 vdd.n2062 0.002
R50593 vdd.n2065 vdd.n2064 0.002
R50594 vdd.n2055 vdd.n2054 0.002
R50595 vdd.n2057 vdd.n2056 0.002
R50596 vdd.n2039 vdd.n2038 0.002
R50597 vdd.n2041 vdd.n2040 0.002
R50598 vdd.n2031 vdd.n2030 0.002
R50599 vdd.n2033 vdd.n2032 0.002
R50600 vdd.n2023 vdd.n2022 0.002
R50601 vdd.n2025 vdd.n2024 0.002
R50602 vdd.n2015 vdd.n2014 0.002
R50603 vdd.n2017 vdd.n2016 0.002
R50604 vdd.n2007 vdd.n2006 0.002
R50605 vdd.n2009 vdd.n2008 0.002
R50606 vdd.n1999 vdd.n1998 0.002
R50607 vdd.n2001 vdd.n2000 0.002
R50608 vdd.n1991 vdd.n1990 0.002
R50609 vdd.n1993 vdd.n1992 0.002
R50610 vdd.n1983 vdd.n1982 0.002
R50611 vdd.n1985 vdd.n1984 0.002
R50612 vdd.n2150 vdd.n2149 0.002
R50613 vdd.n2152 vdd.n2151 0.002
R50614 vdd.n2299 vdd.n2298 0.002
R50615 vdd.n2301 vdd.n2300 0.002
R50616 vdd.n2291 vdd.n2290 0.002
R50617 vdd.n2293 vdd.n2292 0.002
R50618 vdd.n2283 vdd.n2282 0.002
R50619 vdd.n2285 vdd.n2284 0.002
R50620 vdd.n2275 vdd.n2274 0.002
R50621 vdd.n2277 vdd.n2276 0.002
R50622 vdd.n2267 vdd.n2266 0.002
R50623 vdd.n2269 vdd.n2268 0.002
R50624 vdd.n2259 vdd.n2258 0.002
R50625 vdd.n2261 vdd.n2260 0.002
R50626 vdd.n2251 vdd.n2250 0.002
R50627 vdd.n2253 vdd.n2252 0.002
R50628 vdd.n2243 vdd.n2242 0.002
R50629 vdd.n2245 vdd.n2244 0.002
R50630 vdd.n2235 vdd.n2234 0.002
R50631 vdd.n2237 vdd.n2236 0.002
R50632 vdd.n2219 vdd.n2218 0.002
R50633 vdd.n2221 vdd.n2220 0.002
R50634 vdd.n2211 vdd.n2210 0.002
R50635 vdd.n2213 vdd.n2212 0.002
R50636 vdd.n2203 vdd.n2202 0.002
R50637 vdd.n2205 vdd.n2204 0.002
R50638 vdd.n2195 vdd.n2194 0.002
R50639 vdd.n2197 vdd.n2196 0.002
R50640 vdd.n2187 vdd.n2186 0.002
R50641 vdd.n2189 vdd.n2188 0.002
R50642 vdd.n2179 vdd.n2178 0.002
R50643 vdd.n2181 vdd.n2180 0.002
R50644 vdd.n2171 vdd.n2170 0.002
R50645 vdd.n2173 vdd.n2172 0.002
R50646 vdd.n2163 vdd.n2162 0.002
R50647 vdd.n2165 vdd.n2164 0.002
R50648 vdd.n2330 vdd.n2329 0.002
R50649 vdd.n2332 vdd.n2331 0.002
R50650 vdd.n2479 vdd.n2478 0.002
R50651 vdd.n2481 vdd.n2480 0.002
R50652 vdd.n2471 vdd.n2470 0.002
R50653 vdd.n2473 vdd.n2472 0.002
R50654 vdd.n2463 vdd.n2462 0.002
R50655 vdd.n2465 vdd.n2464 0.002
R50656 vdd.n2455 vdd.n2454 0.002
R50657 vdd.n2457 vdd.n2456 0.002
R50658 vdd.n2447 vdd.n2446 0.002
R50659 vdd.n2449 vdd.n2448 0.002
R50660 vdd.n2439 vdd.n2438 0.002
R50661 vdd.n2441 vdd.n2440 0.002
R50662 vdd.n2431 vdd.n2430 0.002
R50663 vdd.n2433 vdd.n2432 0.002
R50664 vdd.n2423 vdd.n2422 0.002
R50665 vdd.n2425 vdd.n2424 0.002
R50666 vdd.n2415 vdd.n2414 0.002
R50667 vdd.n2417 vdd.n2416 0.002
R50668 vdd.n2399 vdd.n2398 0.002
R50669 vdd.n2401 vdd.n2400 0.002
R50670 vdd.n2391 vdd.n2390 0.002
R50671 vdd.n2393 vdd.n2392 0.002
R50672 vdd.n2383 vdd.n2382 0.002
R50673 vdd.n2385 vdd.n2384 0.002
R50674 vdd.n2375 vdd.n2374 0.002
R50675 vdd.n2377 vdd.n2376 0.002
R50676 vdd.n2367 vdd.n2366 0.002
R50677 vdd.n2369 vdd.n2368 0.002
R50678 vdd.n2359 vdd.n2358 0.002
R50679 vdd.n2361 vdd.n2360 0.002
R50680 vdd.n2351 vdd.n2350 0.002
R50681 vdd.n2353 vdd.n2352 0.002
R50682 vdd.n2343 vdd.n2342 0.002
R50683 vdd.n2345 vdd.n2344 0.002
R50684 vdd.n2510 vdd.n2509 0.002
R50685 vdd.n2512 vdd.n2511 0.002
R50686 vdd.n2659 vdd.n2658 0.002
R50687 vdd.n2661 vdd.n2660 0.002
R50688 vdd.n2651 vdd.n2650 0.002
R50689 vdd.n2653 vdd.n2652 0.002
R50690 vdd.n2643 vdd.n2642 0.002
R50691 vdd.n2645 vdd.n2644 0.002
R50692 vdd.n2635 vdd.n2634 0.002
R50693 vdd.n2637 vdd.n2636 0.002
R50694 vdd.n2627 vdd.n2626 0.002
R50695 vdd.n2629 vdd.n2628 0.002
R50696 vdd.n2619 vdd.n2618 0.002
R50697 vdd.n2621 vdd.n2620 0.002
R50698 vdd.n2611 vdd.n2610 0.002
R50699 vdd.n2613 vdd.n2612 0.002
R50700 vdd.n2603 vdd.n2602 0.002
R50701 vdd.n2605 vdd.n2604 0.002
R50702 vdd.n2595 vdd.n2594 0.002
R50703 vdd.n2597 vdd.n2596 0.002
R50704 vdd.n2579 vdd.n2578 0.002
R50705 vdd.n2581 vdd.n2580 0.002
R50706 vdd.n2571 vdd.n2570 0.002
R50707 vdd.n2573 vdd.n2572 0.002
R50708 vdd.n2563 vdd.n2562 0.002
R50709 vdd.n2565 vdd.n2564 0.002
R50710 vdd.n2555 vdd.n2554 0.002
R50711 vdd.n2557 vdd.n2556 0.002
R50712 vdd.n2547 vdd.n2546 0.002
R50713 vdd.n2549 vdd.n2548 0.002
R50714 vdd.n2539 vdd.n2538 0.002
R50715 vdd.n2541 vdd.n2540 0.002
R50716 vdd.n2531 vdd.n2530 0.002
R50717 vdd.n2533 vdd.n2532 0.002
R50718 vdd.n2523 vdd.n2522 0.002
R50719 vdd.n2525 vdd.n2524 0.002
R50720 vdd.n2690 vdd.n2689 0.002
R50721 vdd.n2692 vdd.n2691 0.002
R50722 vdd.n2839 vdd.n2838 0.002
R50723 vdd.n2841 vdd.n2840 0.002
R50724 vdd.n2831 vdd.n2830 0.002
R50725 vdd.n2833 vdd.n2832 0.002
R50726 vdd.n2823 vdd.n2822 0.002
R50727 vdd.n2825 vdd.n2824 0.002
R50728 vdd.n2815 vdd.n2814 0.002
R50729 vdd.n2817 vdd.n2816 0.002
R50730 vdd.n2807 vdd.n2806 0.002
R50731 vdd.n2809 vdd.n2808 0.002
R50732 vdd.n2799 vdd.n2798 0.002
R50733 vdd.n2801 vdd.n2800 0.002
R50734 vdd.n2791 vdd.n2790 0.002
R50735 vdd.n2793 vdd.n2792 0.002
R50736 vdd.n2783 vdd.n2782 0.002
R50737 vdd.n2785 vdd.n2784 0.002
R50738 vdd.n2775 vdd.n2774 0.002
R50739 vdd.n2777 vdd.n2776 0.002
R50740 vdd.n2759 vdd.n2758 0.002
R50741 vdd.n2761 vdd.n2760 0.002
R50742 vdd.n2751 vdd.n2750 0.002
R50743 vdd.n2753 vdd.n2752 0.002
R50744 vdd.n2743 vdd.n2742 0.002
R50745 vdd.n2745 vdd.n2744 0.002
R50746 vdd.n2735 vdd.n2734 0.002
R50747 vdd.n2737 vdd.n2736 0.002
R50748 vdd.n2727 vdd.n2726 0.002
R50749 vdd.n2729 vdd.n2728 0.002
R50750 vdd.n2719 vdd.n2718 0.002
R50751 vdd.n2721 vdd.n2720 0.002
R50752 vdd.n2711 vdd.n2710 0.002
R50753 vdd.n2713 vdd.n2712 0.002
R50754 vdd.n2703 vdd.n2702 0.002
R50755 vdd.n2705 vdd.n2704 0.002
R50756 vdd.n2870 vdd.n2869 0.002
R50757 vdd.n2872 vdd.n2871 0.002
R50758 vdd.n3019 vdd.n3018 0.002
R50759 vdd.n3021 vdd.n3020 0.002
R50760 vdd.n3011 vdd.n3010 0.002
R50761 vdd.n3013 vdd.n3012 0.002
R50762 vdd.n3003 vdd.n3002 0.002
R50763 vdd.n3005 vdd.n3004 0.002
R50764 vdd.n2995 vdd.n2994 0.002
R50765 vdd.n2997 vdd.n2996 0.002
R50766 vdd.n2987 vdd.n2986 0.002
R50767 vdd.n2989 vdd.n2988 0.002
R50768 vdd.n2979 vdd.n2978 0.002
R50769 vdd.n2981 vdd.n2980 0.002
R50770 vdd.n2971 vdd.n2970 0.002
R50771 vdd.n2973 vdd.n2972 0.002
R50772 vdd.n2963 vdd.n2962 0.002
R50773 vdd.n2965 vdd.n2964 0.002
R50774 vdd.n2955 vdd.n2954 0.002
R50775 vdd.n2957 vdd.n2956 0.002
R50776 vdd.n2939 vdd.n2938 0.002
R50777 vdd.n2941 vdd.n2940 0.002
R50778 vdd.n2931 vdd.n2930 0.002
R50779 vdd.n2933 vdd.n2932 0.002
R50780 vdd.n2923 vdd.n2922 0.002
R50781 vdd.n2925 vdd.n2924 0.002
R50782 vdd.n2915 vdd.n2914 0.002
R50783 vdd.n2917 vdd.n2916 0.002
R50784 vdd.n2907 vdd.n2906 0.002
R50785 vdd.n2909 vdd.n2908 0.002
R50786 vdd.n2899 vdd.n2898 0.002
R50787 vdd.n2901 vdd.n2900 0.002
R50788 vdd.n2891 vdd.n2890 0.002
R50789 vdd.n2893 vdd.n2892 0.002
R50790 vdd.n2883 vdd.n2882 0.002
R50791 vdd.n2885 vdd.n2884 0.002
R50792 vdd.n3050 vdd.n3049 0.002
R50793 vdd.n3052 vdd.n3051 0.002
R50794 vdd.n3199 vdd.n3198 0.002
R50795 vdd.n3201 vdd.n3200 0.002
R50796 vdd.n3191 vdd.n3190 0.002
R50797 vdd.n3193 vdd.n3192 0.002
R50798 vdd.n3183 vdd.n3182 0.002
R50799 vdd.n3185 vdd.n3184 0.002
R50800 vdd.n3175 vdd.n3174 0.002
R50801 vdd.n3177 vdd.n3176 0.002
R50802 vdd.n3167 vdd.n3166 0.002
R50803 vdd.n3169 vdd.n3168 0.002
R50804 vdd.n3159 vdd.n3158 0.002
R50805 vdd.n3161 vdd.n3160 0.002
R50806 vdd.n3151 vdd.n3150 0.002
R50807 vdd.n3153 vdd.n3152 0.002
R50808 vdd.n3143 vdd.n3142 0.002
R50809 vdd.n3145 vdd.n3144 0.002
R50810 vdd.n3135 vdd.n3134 0.002
R50811 vdd.n3137 vdd.n3136 0.002
R50812 vdd.n3119 vdd.n3118 0.002
R50813 vdd.n3121 vdd.n3120 0.002
R50814 vdd.n3111 vdd.n3110 0.002
R50815 vdd.n3113 vdd.n3112 0.002
R50816 vdd.n3103 vdd.n3102 0.002
R50817 vdd.n3105 vdd.n3104 0.002
R50818 vdd.n3095 vdd.n3094 0.002
R50819 vdd.n3097 vdd.n3096 0.002
R50820 vdd.n3087 vdd.n3086 0.002
R50821 vdd.n3089 vdd.n3088 0.002
R50822 vdd.n3079 vdd.n3078 0.002
R50823 vdd.n3081 vdd.n3080 0.002
R50824 vdd.n3071 vdd.n3070 0.002
R50825 vdd.n3073 vdd.n3072 0.002
R50826 vdd.n3063 vdd.n3062 0.002
R50827 vdd.n3065 vdd.n3064 0.002
R50828 vdd.n3230 vdd.n3229 0.002
R50829 vdd.n3232 vdd.n3231 0.002
R50830 vdd.n3379 vdd.n3378 0.002
R50831 vdd.n3381 vdd.n3380 0.002
R50832 vdd.n3371 vdd.n3370 0.002
R50833 vdd.n3373 vdd.n3372 0.002
R50834 vdd.n3363 vdd.n3362 0.002
R50835 vdd.n3365 vdd.n3364 0.002
R50836 vdd.n3355 vdd.n3354 0.002
R50837 vdd.n3357 vdd.n3356 0.002
R50838 vdd.n3347 vdd.n3346 0.002
R50839 vdd.n3349 vdd.n3348 0.002
R50840 vdd.n3339 vdd.n3338 0.002
R50841 vdd.n3341 vdd.n3340 0.002
R50842 vdd.n3331 vdd.n3330 0.002
R50843 vdd.n3333 vdd.n3332 0.002
R50844 vdd.n3323 vdd.n3322 0.002
R50845 vdd.n3325 vdd.n3324 0.002
R50846 vdd.n3315 vdd.n3314 0.002
R50847 vdd.n3317 vdd.n3316 0.002
R50848 vdd.n3299 vdd.n3298 0.002
R50849 vdd.n3301 vdd.n3300 0.002
R50850 vdd.n3291 vdd.n3290 0.002
R50851 vdd.n3293 vdd.n3292 0.002
R50852 vdd.n3283 vdd.n3282 0.002
R50853 vdd.n3285 vdd.n3284 0.002
R50854 vdd.n3275 vdd.n3274 0.002
R50855 vdd.n3277 vdd.n3276 0.002
R50856 vdd.n3267 vdd.n3266 0.002
R50857 vdd.n3269 vdd.n3268 0.002
R50858 vdd.n3259 vdd.n3258 0.002
R50859 vdd.n3261 vdd.n3260 0.002
R50860 vdd.n3251 vdd.n3250 0.002
R50861 vdd.n3253 vdd.n3252 0.002
R50862 vdd.n3243 vdd.n3242 0.002
R50863 vdd.n3245 vdd.n3244 0.002
R50864 vdd.n3410 vdd.n3409 0.002
R50865 vdd.n3412 vdd.n3411 0.002
R50866 vdd.n3559 vdd.n3558 0.002
R50867 vdd.n3561 vdd.n3560 0.002
R50868 vdd.n3551 vdd.n3550 0.002
R50869 vdd.n3553 vdd.n3552 0.002
R50870 vdd.n3543 vdd.n3542 0.002
R50871 vdd.n3545 vdd.n3544 0.002
R50872 vdd.n3535 vdd.n3534 0.002
R50873 vdd.n3537 vdd.n3536 0.002
R50874 vdd.n3527 vdd.n3526 0.002
R50875 vdd.n3529 vdd.n3528 0.002
R50876 vdd.n3519 vdd.n3518 0.002
R50877 vdd.n3521 vdd.n3520 0.002
R50878 vdd.n3511 vdd.n3510 0.002
R50879 vdd.n3513 vdd.n3512 0.002
R50880 vdd.n3503 vdd.n3502 0.002
R50881 vdd.n3505 vdd.n3504 0.002
R50882 vdd.n3495 vdd.n3494 0.002
R50883 vdd.n3497 vdd.n3496 0.002
R50884 vdd.n3479 vdd.n3478 0.002
R50885 vdd.n3481 vdd.n3480 0.002
R50886 vdd.n3471 vdd.n3470 0.002
R50887 vdd.n3473 vdd.n3472 0.002
R50888 vdd.n3463 vdd.n3462 0.002
R50889 vdd.n3465 vdd.n3464 0.002
R50890 vdd.n3455 vdd.n3454 0.002
R50891 vdd.n3457 vdd.n3456 0.002
R50892 vdd.n3447 vdd.n3446 0.002
R50893 vdd.n3449 vdd.n3448 0.002
R50894 vdd.n3439 vdd.n3438 0.002
R50895 vdd.n3441 vdd.n3440 0.002
R50896 vdd.n3431 vdd.n3430 0.002
R50897 vdd.n3433 vdd.n3432 0.002
R50898 vdd.n3423 vdd.n3422 0.002
R50899 vdd.n3425 vdd.n3424 0.002
R50900 vdd.n3590 vdd.n3589 0.002
R50901 vdd.n3592 vdd.n3591 0.002
R50902 vdd.n3739 vdd.n3738 0.002
R50903 vdd.n3741 vdd.n3740 0.002
R50904 vdd.n3731 vdd.n3730 0.002
R50905 vdd.n3733 vdd.n3732 0.002
R50906 vdd.n3723 vdd.n3722 0.002
R50907 vdd.n3725 vdd.n3724 0.002
R50908 vdd.n3715 vdd.n3714 0.002
R50909 vdd.n3717 vdd.n3716 0.002
R50910 vdd.n3707 vdd.n3706 0.002
R50911 vdd.n3709 vdd.n3708 0.002
R50912 vdd.n3699 vdd.n3698 0.002
R50913 vdd.n3701 vdd.n3700 0.002
R50914 vdd.n3691 vdd.n3690 0.002
R50915 vdd.n3693 vdd.n3692 0.002
R50916 vdd.n3683 vdd.n3682 0.002
R50917 vdd.n3685 vdd.n3684 0.002
R50918 vdd.n3675 vdd.n3674 0.002
R50919 vdd.n3677 vdd.n3676 0.002
R50920 vdd.n3659 vdd.n3658 0.002
R50921 vdd.n3661 vdd.n3660 0.002
R50922 vdd.n3651 vdd.n3650 0.002
R50923 vdd.n3653 vdd.n3652 0.002
R50924 vdd.n3643 vdd.n3642 0.002
R50925 vdd.n3645 vdd.n3644 0.002
R50926 vdd.n3635 vdd.n3634 0.002
R50927 vdd.n3637 vdd.n3636 0.002
R50928 vdd.n3627 vdd.n3626 0.002
R50929 vdd.n3629 vdd.n3628 0.002
R50930 vdd.n3619 vdd.n3618 0.002
R50931 vdd.n3621 vdd.n3620 0.002
R50932 vdd.n3611 vdd.n3610 0.002
R50933 vdd.n3613 vdd.n3612 0.002
R50934 vdd.n3603 vdd.n3602 0.002
R50935 vdd.n3605 vdd.n3604 0.002
R50936 vdd.n3770 vdd.n3769 0.002
R50937 vdd.n3772 vdd.n3771 0.002
R50938 vdd.n3919 vdd.n3918 0.002
R50939 vdd.n3921 vdd.n3920 0.002
R50940 vdd.n3911 vdd.n3910 0.002
R50941 vdd.n3913 vdd.n3912 0.002
R50942 vdd.n3903 vdd.n3902 0.002
R50943 vdd.n3905 vdd.n3904 0.002
R50944 vdd.n3895 vdd.n3894 0.002
R50945 vdd.n3897 vdd.n3896 0.002
R50946 vdd.n3887 vdd.n3886 0.002
R50947 vdd.n3889 vdd.n3888 0.002
R50948 vdd.n3879 vdd.n3878 0.002
R50949 vdd.n3881 vdd.n3880 0.002
R50950 vdd.n3871 vdd.n3870 0.002
R50951 vdd.n3873 vdd.n3872 0.002
R50952 vdd.n3863 vdd.n3862 0.002
R50953 vdd.n3865 vdd.n3864 0.002
R50954 vdd.n3855 vdd.n3854 0.002
R50955 vdd.n3857 vdd.n3856 0.002
R50956 vdd.n3839 vdd.n3838 0.002
R50957 vdd.n3841 vdd.n3840 0.002
R50958 vdd.n3831 vdd.n3830 0.002
R50959 vdd.n3833 vdd.n3832 0.002
R50960 vdd.n3823 vdd.n3822 0.002
R50961 vdd.n3825 vdd.n3824 0.002
R50962 vdd.n3815 vdd.n3814 0.002
R50963 vdd.n3817 vdd.n3816 0.002
R50964 vdd.n3807 vdd.n3806 0.002
R50965 vdd.n3809 vdd.n3808 0.002
R50966 vdd.n3799 vdd.n3798 0.002
R50967 vdd.n3801 vdd.n3800 0.002
R50968 vdd.n3791 vdd.n3790 0.002
R50969 vdd.n3793 vdd.n3792 0.002
R50970 vdd.n3783 vdd.n3782 0.002
R50971 vdd.n3785 vdd.n3784 0.002
R50972 vdd.n3950 vdd.n3949 0.002
R50973 vdd.n3952 vdd.n3951 0.002
R50974 vdd.n4099 vdd.n4098 0.002
R50975 vdd.n4101 vdd.n4100 0.002
R50976 vdd.n4091 vdd.n4090 0.002
R50977 vdd.n4093 vdd.n4092 0.002
R50978 vdd.n4083 vdd.n4082 0.002
R50979 vdd.n4085 vdd.n4084 0.002
R50980 vdd.n4075 vdd.n4074 0.002
R50981 vdd.n4077 vdd.n4076 0.002
R50982 vdd.n4067 vdd.n4066 0.002
R50983 vdd.n4069 vdd.n4068 0.002
R50984 vdd.n4059 vdd.n4058 0.002
R50985 vdd.n4061 vdd.n4060 0.002
R50986 vdd.n4051 vdd.n4050 0.002
R50987 vdd.n4053 vdd.n4052 0.002
R50988 vdd.n4043 vdd.n4042 0.002
R50989 vdd.n4045 vdd.n4044 0.002
R50990 vdd.n4035 vdd.n4034 0.002
R50991 vdd.n4037 vdd.n4036 0.002
R50992 vdd.n4019 vdd.n4018 0.002
R50993 vdd.n4021 vdd.n4020 0.002
R50994 vdd.n4011 vdd.n4010 0.002
R50995 vdd.n4013 vdd.n4012 0.002
R50996 vdd.n4003 vdd.n4002 0.002
R50997 vdd.n4005 vdd.n4004 0.002
R50998 vdd.n3995 vdd.n3994 0.002
R50999 vdd.n3997 vdd.n3996 0.002
R51000 vdd.n3987 vdd.n3986 0.002
R51001 vdd.n3989 vdd.n3988 0.002
R51002 vdd.n3979 vdd.n3978 0.002
R51003 vdd.n3981 vdd.n3980 0.002
R51004 vdd.n3971 vdd.n3970 0.002
R51005 vdd.n3973 vdd.n3972 0.002
R51006 vdd.n3963 vdd.n3962 0.002
R51007 vdd.n3965 vdd.n3964 0.002
R51008 vdd.n4130 vdd.n4129 0.002
R51009 vdd.n4132 vdd.n4131 0.002
R51010 vdd.n4279 vdd.n4278 0.002
R51011 vdd.n4281 vdd.n4280 0.002
R51012 vdd.n4271 vdd.n4270 0.002
R51013 vdd.n4273 vdd.n4272 0.002
R51014 vdd.n4263 vdd.n4262 0.002
R51015 vdd.n4265 vdd.n4264 0.002
R51016 vdd.n4255 vdd.n4254 0.002
R51017 vdd.n4257 vdd.n4256 0.002
R51018 vdd.n4247 vdd.n4246 0.002
R51019 vdd.n4249 vdd.n4248 0.002
R51020 vdd.n4239 vdd.n4238 0.002
R51021 vdd.n4241 vdd.n4240 0.002
R51022 vdd.n4231 vdd.n4230 0.002
R51023 vdd.n4233 vdd.n4232 0.002
R51024 vdd.n4223 vdd.n4222 0.002
R51025 vdd.n4225 vdd.n4224 0.002
R51026 vdd.n4215 vdd.n4214 0.002
R51027 vdd.n4217 vdd.n4216 0.002
R51028 vdd.n4199 vdd.n4198 0.002
R51029 vdd.n4201 vdd.n4200 0.002
R51030 vdd.n4191 vdd.n4190 0.002
R51031 vdd.n4193 vdd.n4192 0.002
R51032 vdd.n4183 vdd.n4182 0.002
R51033 vdd.n4185 vdd.n4184 0.002
R51034 vdd.n4175 vdd.n4174 0.002
R51035 vdd.n4177 vdd.n4176 0.002
R51036 vdd.n4167 vdd.n4166 0.002
R51037 vdd.n4169 vdd.n4168 0.002
R51038 vdd.n4159 vdd.n4158 0.002
R51039 vdd.n4161 vdd.n4160 0.002
R51040 vdd.n4151 vdd.n4150 0.002
R51041 vdd.n4153 vdd.n4152 0.002
R51042 vdd.n4143 vdd.n4142 0.002
R51043 vdd.n4145 vdd.n4144 0.002
R51044 vdd.n4310 vdd.n4309 0.002
R51045 vdd.n4312 vdd.n4311 0.002
R51046 vdd.n4459 vdd.n4458 0.002
R51047 vdd.n4461 vdd.n4460 0.002
R51048 vdd.n4451 vdd.n4450 0.002
R51049 vdd.n4453 vdd.n4452 0.002
R51050 vdd.n4443 vdd.n4442 0.002
R51051 vdd.n4445 vdd.n4444 0.002
R51052 vdd.n4435 vdd.n4434 0.002
R51053 vdd.n4437 vdd.n4436 0.002
R51054 vdd.n4427 vdd.n4426 0.002
R51055 vdd.n4429 vdd.n4428 0.002
R51056 vdd.n4419 vdd.n4418 0.002
R51057 vdd.n4421 vdd.n4420 0.002
R51058 vdd.n4411 vdd.n4410 0.002
R51059 vdd.n4413 vdd.n4412 0.002
R51060 vdd.n4403 vdd.n4402 0.002
R51061 vdd.n4405 vdd.n4404 0.002
R51062 vdd.n4395 vdd.n4394 0.002
R51063 vdd.n4397 vdd.n4396 0.002
R51064 vdd.n4379 vdd.n4378 0.002
R51065 vdd.n4381 vdd.n4380 0.002
R51066 vdd.n4371 vdd.n4370 0.002
R51067 vdd.n4373 vdd.n4372 0.002
R51068 vdd.n4363 vdd.n4362 0.002
R51069 vdd.n4365 vdd.n4364 0.002
R51070 vdd.n4355 vdd.n4354 0.002
R51071 vdd.n4357 vdd.n4356 0.002
R51072 vdd.n4347 vdd.n4346 0.002
R51073 vdd.n4349 vdd.n4348 0.002
R51074 vdd.n4339 vdd.n4338 0.002
R51075 vdd.n4341 vdd.n4340 0.002
R51076 vdd.n4331 vdd.n4330 0.002
R51077 vdd.n4333 vdd.n4332 0.002
R51078 vdd.n4323 vdd.n4322 0.002
R51079 vdd.n4325 vdd.n4324 0.002
R51080 vdd.n4490 vdd.n4489 0.002
R51081 vdd.n4492 vdd.n4491 0.002
R51082 vdd.n4639 vdd.n4638 0.002
R51083 vdd.n4641 vdd.n4640 0.002
R51084 vdd.n4631 vdd.n4630 0.002
R51085 vdd.n4633 vdd.n4632 0.002
R51086 vdd.n4623 vdd.n4622 0.002
R51087 vdd.n4625 vdd.n4624 0.002
R51088 vdd.n4615 vdd.n4614 0.002
R51089 vdd.n4617 vdd.n4616 0.002
R51090 vdd.n4607 vdd.n4606 0.002
R51091 vdd.n4609 vdd.n4608 0.002
R51092 vdd.n4599 vdd.n4598 0.002
R51093 vdd.n4601 vdd.n4600 0.002
R51094 vdd.n4591 vdd.n4590 0.002
R51095 vdd.n4593 vdd.n4592 0.002
R51096 vdd.n4583 vdd.n4582 0.002
R51097 vdd.n4585 vdd.n4584 0.002
R51098 vdd.n4575 vdd.n4574 0.002
R51099 vdd.n4577 vdd.n4576 0.002
R51100 vdd.n4559 vdd.n4558 0.002
R51101 vdd.n4561 vdd.n4560 0.002
R51102 vdd.n4551 vdd.n4550 0.002
R51103 vdd.n4553 vdd.n4552 0.002
R51104 vdd.n4543 vdd.n4542 0.002
R51105 vdd.n4545 vdd.n4544 0.002
R51106 vdd.n4535 vdd.n4534 0.002
R51107 vdd.n4537 vdd.n4536 0.002
R51108 vdd.n4527 vdd.n4526 0.002
R51109 vdd.n4529 vdd.n4528 0.002
R51110 vdd.n4519 vdd.n4518 0.002
R51111 vdd.n4521 vdd.n4520 0.002
R51112 vdd.n4511 vdd.n4510 0.002
R51113 vdd.n4513 vdd.n4512 0.002
R51114 vdd.n4503 vdd.n4502 0.002
R51115 vdd.n4505 vdd.n4504 0.002
R51116 vdd.n4670 vdd.n4669 0.002
R51117 vdd.n4672 vdd.n4671 0.002
R51118 vdd.n4819 vdd.n4818 0.002
R51119 vdd.n4821 vdd.n4820 0.002
R51120 vdd.n4811 vdd.n4810 0.002
R51121 vdd.n4813 vdd.n4812 0.002
R51122 vdd.n4803 vdd.n4802 0.002
R51123 vdd.n4805 vdd.n4804 0.002
R51124 vdd.n4795 vdd.n4794 0.002
R51125 vdd.n4797 vdd.n4796 0.002
R51126 vdd.n4787 vdd.n4786 0.002
R51127 vdd.n4789 vdd.n4788 0.002
R51128 vdd.n4779 vdd.n4778 0.002
R51129 vdd.n4781 vdd.n4780 0.002
R51130 vdd.n4771 vdd.n4770 0.002
R51131 vdd.n4773 vdd.n4772 0.002
R51132 vdd.n4763 vdd.n4762 0.002
R51133 vdd.n4765 vdd.n4764 0.002
R51134 vdd.n4755 vdd.n4754 0.002
R51135 vdd.n4757 vdd.n4756 0.002
R51136 vdd.n4739 vdd.n4738 0.002
R51137 vdd.n4741 vdd.n4740 0.002
R51138 vdd.n4731 vdd.n4730 0.002
R51139 vdd.n4733 vdd.n4732 0.002
R51140 vdd.n4723 vdd.n4722 0.002
R51141 vdd.n4725 vdd.n4724 0.002
R51142 vdd.n4715 vdd.n4714 0.002
R51143 vdd.n4717 vdd.n4716 0.002
R51144 vdd.n4707 vdd.n4706 0.002
R51145 vdd.n4709 vdd.n4708 0.002
R51146 vdd.n4699 vdd.n4698 0.002
R51147 vdd.n4701 vdd.n4700 0.002
R51148 vdd.n4691 vdd.n4690 0.002
R51149 vdd.n4693 vdd.n4692 0.002
R51150 vdd.n4683 vdd.n4682 0.002
R51151 vdd.n4685 vdd.n4684 0.002
R51152 vdd.n4850 vdd.n4849 0.002
R51153 vdd.n4852 vdd.n4851 0.002
R51154 vdd.n4999 vdd.n4998 0.002
R51155 vdd.n5001 vdd.n5000 0.002
R51156 vdd.n4991 vdd.n4990 0.002
R51157 vdd.n4993 vdd.n4992 0.002
R51158 vdd.n4983 vdd.n4982 0.002
R51159 vdd.n4985 vdd.n4984 0.002
R51160 vdd.n4975 vdd.n4974 0.002
R51161 vdd.n4977 vdd.n4976 0.002
R51162 vdd.n4967 vdd.n4966 0.002
R51163 vdd.n4969 vdd.n4968 0.002
R51164 vdd.n4959 vdd.n4958 0.002
R51165 vdd.n4961 vdd.n4960 0.002
R51166 vdd.n4951 vdd.n4950 0.002
R51167 vdd.n4953 vdd.n4952 0.002
R51168 vdd.n4943 vdd.n4942 0.002
R51169 vdd.n4945 vdd.n4944 0.002
R51170 vdd.n4935 vdd.n4934 0.002
R51171 vdd.n4937 vdd.n4936 0.002
R51172 vdd.n4919 vdd.n4918 0.002
R51173 vdd.n4921 vdd.n4920 0.002
R51174 vdd.n4911 vdd.n4910 0.002
R51175 vdd.n4913 vdd.n4912 0.002
R51176 vdd.n4903 vdd.n4902 0.002
R51177 vdd.n4905 vdd.n4904 0.002
R51178 vdd.n4895 vdd.n4894 0.002
R51179 vdd.n4897 vdd.n4896 0.002
R51180 vdd.n4887 vdd.n4886 0.002
R51181 vdd.n4889 vdd.n4888 0.002
R51182 vdd.n4879 vdd.n4878 0.002
R51183 vdd.n4881 vdd.n4880 0.002
R51184 vdd.n4871 vdd.n4870 0.002
R51185 vdd.n4873 vdd.n4872 0.002
R51186 vdd.n4863 vdd.n4862 0.002
R51187 vdd.n4865 vdd.n4864 0.002
R51188 vdd.n5030 vdd.n5029 0.002
R51189 vdd.n5032 vdd.n5031 0.002
R51190 vdd.n5179 vdd.n5178 0.002
R51191 vdd.n5181 vdd.n5180 0.002
R51192 vdd.n5171 vdd.n5170 0.002
R51193 vdd.n5173 vdd.n5172 0.002
R51194 vdd.n5163 vdd.n5162 0.002
R51195 vdd.n5165 vdd.n5164 0.002
R51196 vdd.n5155 vdd.n5154 0.002
R51197 vdd.n5157 vdd.n5156 0.002
R51198 vdd.n5147 vdd.n5146 0.002
R51199 vdd.n5149 vdd.n5148 0.002
R51200 vdd.n5139 vdd.n5138 0.002
R51201 vdd.n5141 vdd.n5140 0.002
R51202 vdd.n5131 vdd.n5130 0.002
R51203 vdd.n5133 vdd.n5132 0.002
R51204 vdd.n5123 vdd.n5122 0.002
R51205 vdd.n5125 vdd.n5124 0.002
R51206 vdd.n5115 vdd.n5114 0.002
R51207 vdd.n5117 vdd.n5116 0.002
R51208 vdd.n5099 vdd.n5098 0.002
R51209 vdd.n5101 vdd.n5100 0.002
R51210 vdd.n5091 vdd.n5090 0.002
R51211 vdd.n5093 vdd.n5092 0.002
R51212 vdd.n5083 vdd.n5082 0.002
R51213 vdd.n5085 vdd.n5084 0.002
R51214 vdd.n5075 vdd.n5074 0.002
R51215 vdd.n5077 vdd.n5076 0.002
R51216 vdd.n5067 vdd.n5066 0.002
R51217 vdd.n5069 vdd.n5068 0.002
R51218 vdd.n5059 vdd.n5058 0.002
R51219 vdd.n5061 vdd.n5060 0.002
R51220 vdd.n5051 vdd.n5050 0.002
R51221 vdd.n5053 vdd.n5052 0.002
R51222 vdd.n5043 vdd.n5042 0.002
R51223 vdd.n5045 vdd.n5044 0.002
R51224 vdd.n5210 vdd.n5209 0.002
R51225 vdd.n5212 vdd.n5211 0.002
R51226 vdd.n5359 vdd.n5358 0.002
R51227 vdd.n5361 vdd.n5360 0.002
R51228 vdd.n5351 vdd.n5350 0.002
R51229 vdd.n5353 vdd.n5352 0.002
R51230 vdd.n5343 vdd.n5342 0.002
R51231 vdd.n5345 vdd.n5344 0.002
R51232 vdd.n5335 vdd.n5334 0.002
R51233 vdd.n5337 vdd.n5336 0.002
R51234 vdd.n5327 vdd.n5326 0.002
R51235 vdd.n5329 vdd.n5328 0.002
R51236 vdd.n5319 vdd.n5318 0.002
R51237 vdd.n5321 vdd.n5320 0.002
R51238 vdd.n5311 vdd.n5310 0.002
R51239 vdd.n5313 vdd.n5312 0.002
R51240 vdd.n5303 vdd.n5302 0.002
R51241 vdd.n5305 vdd.n5304 0.002
R51242 vdd.n5295 vdd.n5294 0.002
R51243 vdd.n5297 vdd.n5296 0.002
R51244 vdd.n5279 vdd.n5278 0.002
R51245 vdd.n5281 vdd.n5280 0.002
R51246 vdd.n5271 vdd.n5270 0.002
R51247 vdd.n5273 vdd.n5272 0.002
R51248 vdd.n5263 vdd.n5262 0.002
R51249 vdd.n5265 vdd.n5264 0.002
R51250 vdd.n5255 vdd.n5254 0.002
R51251 vdd.n5257 vdd.n5256 0.002
R51252 vdd.n5247 vdd.n5246 0.002
R51253 vdd.n5249 vdd.n5248 0.002
R51254 vdd.n5239 vdd.n5238 0.002
R51255 vdd.n5241 vdd.n5240 0.002
R51256 vdd.n5231 vdd.n5230 0.002
R51257 vdd.n5233 vdd.n5232 0.002
R51258 vdd.n5223 vdd.n5222 0.002
R51259 vdd.n5225 vdd.n5224 0.002
R51260 vdd.n5390 vdd.n5389 0.002
R51261 vdd.n5392 vdd.n5391 0.002
R51262 vdd.n5539 vdd.n5538 0.002
R51263 vdd.n5541 vdd.n5540 0.002
R51264 vdd.n5531 vdd.n5530 0.002
R51265 vdd.n5533 vdd.n5532 0.002
R51266 vdd.n5523 vdd.n5522 0.002
R51267 vdd.n5525 vdd.n5524 0.002
R51268 vdd.n5515 vdd.n5514 0.002
R51269 vdd.n5517 vdd.n5516 0.002
R51270 vdd.n5507 vdd.n5506 0.002
R51271 vdd.n5509 vdd.n5508 0.002
R51272 vdd.n5499 vdd.n5498 0.002
R51273 vdd.n5501 vdd.n5500 0.002
R51274 vdd.n5491 vdd.n5490 0.002
R51275 vdd.n5493 vdd.n5492 0.002
R51276 vdd.n5483 vdd.n5482 0.002
R51277 vdd.n5485 vdd.n5484 0.002
R51278 vdd.n5475 vdd.n5474 0.002
R51279 vdd.n5477 vdd.n5476 0.002
R51280 vdd.n5459 vdd.n5458 0.002
R51281 vdd.n5461 vdd.n5460 0.002
R51282 vdd.n5451 vdd.n5450 0.002
R51283 vdd.n5453 vdd.n5452 0.002
R51284 vdd.n5443 vdd.n5442 0.002
R51285 vdd.n5445 vdd.n5444 0.002
R51286 vdd.n5435 vdd.n5434 0.002
R51287 vdd.n5437 vdd.n5436 0.002
R51288 vdd.n5427 vdd.n5426 0.002
R51289 vdd.n5429 vdd.n5428 0.002
R51290 vdd.n5419 vdd.n5418 0.002
R51291 vdd.n5421 vdd.n5420 0.002
R51292 vdd.n5411 vdd.n5410 0.002
R51293 vdd.n5413 vdd.n5412 0.002
R51294 vdd.n5403 vdd.n5402 0.002
R51295 vdd.n5405 vdd.n5404 0.002
R51296 vdd.n5570 vdd.n5569 0.002
R51297 vdd.n5572 vdd.n5571 0.002
R51298 vdd.n5719 vdd.n5718 0.002
R51299 vdd.n5721 vdd.n5720 0.002
R51300 vdd.n5711 vdd.n5710 0.002
R51301 vdd.n5713 vdd.n5712 0.002
R51302 vdd.n5703 vdd.n5702 0.002
R51303 vdd.n5705 vdd.n5704 0.002
R51304 vdd.n5695 vdd.n5694 0.002
R51305 vdd.n5697 vdd.n5696 0.002
R51306 vdd.n5687 vdd.n5686 0.002
R51307 vdd.n5689 vdd.n5688 0.002
R51308 vdd.n5679 vdd.n5678 0.002
R51309 vdd.n5681 vdd.n5680 0.002
R51310 vdd.n5671 vdd.n5670 0.002
R51311 vdd.n5673 vdd.n5672 0.002
R51312 vdd.n5663 vdd.n5662 0.002
R51313 vdd.n5665 vdd.n5664 0.002
R51314 vdd.n5655 vdd.n5654 0.002
R51315 vdd.n5657 vdd.n5656 0.002
R51316 vdd.n5639 vdd.n5638 0.002
R51317 vdd.n5641 vdd.n5640 0.002
R51318 vdd.n5631 vdd.n5630 0.002
R51319 vdd.n5633 vdd.n5632 0.002
R51320 vdd.n5623 vdd.n5622 0.002
R51321 vdd.n5625 vdd.n5624 0.002
R51322 vdd.n5615 vdd.n5614 0.002
R51323 vdd.n5617 vdd.n5616 0.002
R51324 vdd.n5607 vdd.n5606 0.002
R51325 vdd.n5609 vdd.n5608 0.002
R51326 vdd.n5599 vdd.n5598 0.002
R51327 vdd.n5601 vdd.n5600 0.002
R51328 vdd.n5591 vdd.n5590 0.002
R51329 vdd.n5593 vdd.n5592 0.002
R51330 vdd.n5583 vdd.n5582 0.002
R51331 vdd.n5585 vdd.n5584 0.002
R51332 vdd.n5750 vdd.n5749 0.002
R51333 vdd.n5752 vdd.n5751 0.002
R51334 vdd.n5899 vdd.n5898 0.002
R51335 vdd.n5901 vdd.n5900 0.002
R51336 vdd.n5891 vdd.n5890 0.002
R51337 vdd.n5893 vdd.n5892 0.002
R51338 vdd.n5883 vdd.n5882 0.002
R51339 vdd.n5885 vdd.n5884 0.002
R51340 vdd.n5875 vdd.n5874 0.002
R51341 vdd.n5877 vdd.n5876 0.002
R51342 vdd.n5867 vdd.n5866 0.002
R51343 vdd.n5869 vdd.n5868 0.002
R51344 vdd.n5859 vdd.n5858 0.002
R51345 vdd.n5861 vdd.n5860 0.002
R51346 vdd.n5851 vdd.n5850 0.002
R51347 vdd.n5853 vdd.n5852 0.002
R51348 vdd.n5843 vdd.n5842 0.002
R51349 vdd.n5845 vdd.n5844 0.002
R51350 vdd.n5835 vdd.n5834 0.002
R51351 vdd.n5837 vdd.n5836 0.002
R51352 vdd.n5819 vdd.n5818 0.002
R51353 vdd.n5821 vdd.n5820 0.002
R51354 vdd.n5811 vdd.n5810 0.002
R51355 vdd.n5813 vdd.n5812 0.002
R51356 vdd.n5803 vdd.n5802 0.002
R51357 vdd.n5805 vdd.n5804 0.002
R51358 vdd.n5795 vdd.n5794 0.002
R51359 vdd.n5797 vdd.n5796 0.002
R51360 vdd.n5787 vdd.n5786 0.002
R51361 vdd.n5789 vdd.n5788 0.002
R51362 vdd.n5779 vdd.n5778 0.002
R51363 vdd.n5781 vdd.n5780 0.002
R51364 vdd.n5771 vdd.n5770 0.002
R51365 vdd.n5773 vdd.n5772 0.002
R51366 vdd.n5763 vdd.n5762 0.002
R51367 vdd.n5765 vdd.n5764 0.002
R51368 vdd.n5930 vdd.n5929 0.002
R51369 vdd.n5932 vdd.n5931 0.002
R51370 vdd.n6079 vdd.n6078 0.002
R51371 vdd.n6081 vdd.n6080 0.002
R51372 vdd.n6071 vdd.n6070 0.002
R51373 vdd.n6073 vdd.n6072 0.002
R51374 vdd.n6063 vdd.n6062 0.002
R51375 vdd.n6065 vdd.n6064 0.002
R51376 vdd.n6055 vdd.n6054 0.002
R51377 vdd.n6057 vdd.n6056 0.002
R51378 vdd.n6047 vdd.n6046 0.002
R51379 vdd.n6049 vdd.n6048 0.002
R51380 vdd.n6039 vdd.n6038 0.002
R51381 vdd.n6041 vdd.n6040 0.002
R51382 vdd.n6031 vdd.n6030 0.002
R51383 vdd.n6033 vdd.n6032 0.002
R51384 vdd.n6023 vdd.n6022 0.002
R51385 vdd.n6025 vdd.n6024 0.002
R51386 vdd.n6015 vdd.n6014 0.002
R51387 vdd.n6017 vdd.n6016 0.002
R51388 vdd.n5999 vdd.n5998 0.002
R51389 vdd.n6001 vdd.n6000 0.002
R51390 vdd.n5991 vdd.n5990 0.002
R51391 vdd.n5993 vdd.n5992 0.002
R51392 vdd.n5983 vdd.n5982 0.002
R51393 vdd.n5985 vdd.n5984 0.002
R51394 vdd.n5975 vdd.n5974 0.002
R51395 vdd.n5977 vdd.n5976 0.002
R51396 vdd.n5967 vdd.n5966 0.002
R51397 vdd.n5969 vdd.n5968 0.002
R51398 vdd.n5959 vdd.n5958 0.002
R51399 vdd.n5961 vdd.n5960 0.002
R51400 vdd.n5951 vdd.n5950 0.002
R51401 vdd.n5953 vdd.n5952 0.002
R51402 vdd.n5943 vdd.n5942 0.002
R51403 vdd.n5945 vdd.n5944 0.002
R51404 vdd.n6110 vdd.n6109 0.002
R51405 vdd.n6112 vdd.n6111 0.002
R51406 vdd.n6259 vdd.n6258 0.002
R51407 vdd.n6261 vdd.n6260 0.002
R51408 vdd.n6251 vdd.n6250 0.002
R51409 vdd.n6253 vdd.n6252 0.002
R51410 vdd.n6243 vdd.n6242 0.002
R51411 vdd.n6245 vdd.n6244 0.002
R51412 vdd.n6235 vdd.n6234 0.002
R51413 vdd.n6237 vdd.n6236 0.002
R51414 vdd.n6227 vdd.n6226 0.002
R51415 vdd.n6229 vdd.n6228 0.002
R51416 vdd.n6219 vdd.n6218 0.002
R51417 vdd.n6221 vdd.n6220 0.002
R51418 vdd.n6211 vdd.n6210 0.002
R51419 vdd.n6213 vdd.n6212 0.002
R51420 vdd.n6203 vdd.n6202 0.002
R51421 vdd.n6205 vdd.n6204 0.002
R51422 vdd.n6195 vdd.n6194 0.002
R51423 vdd.n6197 vdd.n6196 0.002
R51424 vdd.n6179 vdd.n6178 0.002
R51425 vdd.n6181 vdd.n6180 0.002
R51426 vdd.n6171 vdd.n6170 0.002
R51427 vdd.n6173 vdd.n6172 0.002
R51428 vdd.n6163 vdd.n6162 0.002
R51429 vdd.n6165 vdd.n6164 0.002
R51430 vdd.n6155 vdd.n6154 0.002
R51431 vdd.n6157 vdd.n6156 0.002
R51432 vdd.n6147 vdd.n6146 0.002
R51433 vdd.n6149 vdd.n6148 0.002
R51434 vdd.n6139 vdd.n6138 0.002
R51435 vdd.n6141 vdd.n6140 0.002
R51436 vdd.n6131 vdd.n6130 0.002
R51437 vdd.n6133 vdd.n6132 0.002
R51438 vdd.n6123 vdd.n6122 0.002
R51439 vdd.n6125 vdd.n6124 0.002
R51440 vdd.n6290 vdd.n6289 0.002
R51441 vdd.n6292 vdd.n6291 0.002
R51442 vdd.n6439 vdd.n6438 0.002
R51443 vdd.n6441 vdd.n6440 0.002
R51444 vdd.n6431 vdd.n6430 0.002
R51445 vdd.n6433 vdd.n6432 0.002
R51446 vdd.n6423 vdd.n6422 0.002
R51447 vdd.n6425 vdd.n6424 0.002
R51448 vdd.n6415 vdd.n6414 0.002
R51449 vdd.n6417 vdd.n6416 0.002
R51450 vdd.n6407 vdd.n6406 0.002
R51451 vdd.n6409 vdd.n6408 0.002
R51452 vdd.n6399 vdd.n6398 0.002
R51453 vdd.n6401 vdd.n6400 0.002
R51454 vdd.n6391 vdd.n6390 0.002
R51455 vdd.n6393 vdd.n6392 0.002
R51456 vdd.n6383 vdd.n6382 0.002
R51457 vdd.n6385 vdd.n6384 0.002
R51458 vdd.n6375 vdd.n6374 0.002
R51459 vdd.n6377 vdd.n6376 0.002
R51460 vdd.n6359 vdd.n6358 0.002
R51461 vdd.n6361 vdd.n6360 0.002
R51462 vdd.n6351 vdd.n6350 0.002
R51463 vdd.n6353 vdd.n6352 0.002
R51464 vdd.n6343 vdd.n6342 0.002
R51465 vdd.n6345 vdd.n6344 0.002
R51466 vdd.n6335 vdd.n6334 0.002
R51467 vdd.n6337 vdd.n6336 0.002
R51468 vdd.n6327 vdd.n6326 0.002
R51469 vdd.n6329 vdd.n6328 0.002
R51470 vdd.n6319 vdd.n6318 0.002
R51471 vdd.n6321 vdd.n6320 0.002
R51472 vdd.n6311 vdd.n6310 0.002
R51473 vdd.n6313 vdd.n6312 0.002
R51474 vdd.n6303 vdd.n6302 0.002
R51475 vdd.n6305 vdd.n6304 0.002
R51476 vdd.n6470 vdd.n6469 0.002
R51477 vdd.n6472 vdd.n6471 0.002
R51478 vdd.n6619 vdd.n6618 0.002
R51479 vdd.n6621 vdd.n6620 0.002
R51480 vdd.n6611 vdd.n6610 0.002
R51481 vdd.n6613 vdd.n6612 0.002
R51482 vdd.n6603 vdd.n6602 0.002
R51483 vdd.n6605 vdd.n6604 0.002
R51484 vdd.n6595 vdd.n6594 0.002
R51485 vdd.n6597 vdd.n6596 0.002
R51486 vdd.n6587 vdd.n6586 0.002
R51487 vdd.n6589 vdd.n6588 0.002
R51488 vdd.n6579 vdd.n6578 0.002
R51489 vdd.n6581 vdd.n6580 0.002
R51490 vdd.n6571 vdd.n6570 0.002
R51491 vdd.n6573 vdd.n6572 0.002
R51492 vdd.n6563 vdd.n6562 0.002
R51493 vdd.n6565 vdd.n6564 0.002
R51494 vdd.n6555 vdd.n6554 0.002
R51495 vdd.n6557 vdd.n6556 0.002
R51496 vdd.n6539 vdd.n6538 0.002
R51497 vdd.n6541 vdd.n6540 0.002
R51498 vdd.n6531 vdd.n6530 0.002
R51499 vdd.n6533 vdd.n6532 0.002
R51500 vdd.n6523 vdd.n6522 0.002
R51501 vdd.n6525 vdd.n6524 0.002
R51502 vdd.n6515 vdd.n6514 0.002
R51503 vdd.n6517 vdd.n6516 0.002
R51504 vdd.n6507 vdd.n6506 0.002
R51505 vdd.n6509 vdd.n6508 0.002
R51506 vdd.n6499 vdd.n6498 0.002
R51507 vdd.n6501 vdd.n6500 0.002
R51508 vdd.n6491 vdd.n6490 0.002
R51509 vdd.n6493 vdd.n6492 0.002
R51510 vdd.n6483 vdd.n6482 0.002
R51511 vdd.n6485 vdd.n6484 0.002
R51512 vdd.n6650 vdd.n6649 0.002
R51513 vdd.n6652 vdd.n6651 0.002
R51514 vdd.n6799 vdd.n6798 0.002
R51515 vdd.n6801 vdd.n6800 0.002
R51516 vdd.n6791 vdd.n6790 0.002
R51517 vdd.n6793 vdd.n6792 0.002
R51518 vdd.n6783 vdd.n6782 0.002
R51519 vdd.n6785 vdd.n6784 0.002
R51520 vdd.n6775 vdd.n6774 0.002
R51521 vdd.n6777 vdd.n6776 0.002
R51522 vdd.n6767 vdd.n6766 0.002
R51523 vdd.n6769 vdd.n6768 0.002
R51524 vdd.n6759 vdd.n6758 0.002
R51525 vdd.n6761 vdd.n6760 0.002
R51526 vdd.n6751 vdd.n6750 0.002
R51527 vdd.n6753 vdd.n6752 0.002
R51528 vdd.n6743 vdd.n6742 0.002
R51529 vdd.n6745 vdd.n6744 0.002
R51530 vdd.n6735 vdd.n6734 0.002
R51531 vdd.n6737 vdd.n6736 0.002
R51532 vdd.n6719 vdd.n6718 0.002
R51533 vdd.n6721 vdd.n6720 0.002
R51534 vdd.n6711 vdd.n6710 0.002
R51535 vdd.n6713 vdd.n6712 0.002
R51536 vdd.n6703 vdd.n6702 0.002
R51537 vdd.n6705 vdd.n6704 0.002
R51538 vdd.n6695 vdd.n6694 0.002
R51539 vdd.n6697 vdd.n6696 0.002
R51540 vdd.n6687 vdd.n6686 0.002
R51541 vdd.n6689 vdd.n6688 0.002
R51542 vdd.n6679 vdd.n6678 0.002
R51543 vdd.n6681 vdd.n6680 0.002
R51544 vdd.n6671 vdd.n6670 0.002
R51545 vdd.n6673 vdd.n6672 0.002
R51546 vdd.n6663 vdd.n6662 0.002
R51547 vdd.n6665 vdd.n6664 0.002
R51548 vdd.n6830 vdd.n6829 0.002
R51549 vdd.n6832 vdd.n6831 0.002
R51550 vdd.n6979 vdd.n6978 0.002
R51551 vdd.n6981 vdd.n6980 0.002
R51552 vdd.n6971 vdd.n6970 0.002
R51553 vdd.n6973 vdd.n6972 0.002
R51554 vdd.n6963 vdd.n6962 0.002
R51555 vdd.n6965 vdd.n6964 0.002
R51556 vdd.n6955 vdd.n6954 0.002
R51557 vdd.n6957 vdd.n6956 0.002
R51558 vdd.n6947 vdd.n6946 0.002
R51559 vdd.n6949 vdd.n6948 0.002
R51560 vdd.n6939 vdd.n6938 0.002
R51561 vdd.n6941 vdd.n6940 0.002
R51562 vdd.n6931 vdd.n6930 0.002
R51563 vdd.n6933 vdd.n6932 0.002
R51564 vdd.n6923 vdd.n6922 0.002
R51565 vdd.n6925 vdd.n6924 0.002
R51566 vdd.n6915 vdd.n6914 0.002
R51567 vdd.n6917 vdd.n6916 0.002
R51568 vdd.n6899 vdd.n6898 0.002
R51569 vdd.n6901 vdd.n6900 0.002
R51570 vdd.n6891 vdd.n6890 0.002
R51571 vdd.n6893 vdd.n6892 0.002
R51572 vdd.n6883 vdd.n6882 0.002
R51573 vdd.n6885 vdd.n6884 0.002
R51574 vdd.n6875 vdd.n6874 0.002
R51575 vdd.n6877 vdd.n6876 0.002
R51576 vdd.n6867 vdd.n6866 0.002
R51577 vdd.n6869 vdd.n6868 0.002
R51578 vdd.n6859 vdd.n6858 0.002
R51579 vdd.n6861 vdd.n6860 0.002
R51580 vdd.n6851 vdd.n6850 0.002
R51581 vdd.n6853 vdd.n6852 0.002
R51582 vdd.n6843 vdd.n6842 0.002
R51583 vdd.n6845 vdd.n6844 0.002
R51584 vdd.n7010 vdd.n7009 0.002
R51585 vdd.n7012 vdd.n7011 0.002
R51586 vdd.n7159 vdd.n7158 0.002
R51587 vdd.n7161 vdd.n7160 0.002
R51588 vdd.n7151 vdd.n7150 0.002
R51589 vdd.n7153 vdd.n7152 0.002
R51590 vdd.n7143 vdd.n7142 0.002
R51591 vdd.n7145 vdd.n7144 0.002
R51592 vdd.n7135 vdd.n7134 0.002
R51593 vdd.n7137 vdd.n7136 0.002
R51594 vdd.n7127 vdd.n7126 0.002
R51595 vdd.n7129 vdd.n7128 0.002
R51596 vdd.n7119 vdd.n7118 0.002
R51597 vdd.n7121 vdd.n7120 0.002
R51598 vdd.n7111 vdd.n7110 0.002
R51599 vdd.n7113 vdd.n7112 0.002
R51600 vdd.n7103 vdd.n7102 0.002
R51601 vdd.n7105 vdd.n7104 0.002
R51602 vdd.n7095 vdd.n7094 0.002
R51603 vdd.n7097 vdd.n7096 0.002
R51604 vdd.n7079 vdd.n7078 0.002
R51605 vdd.n7081 vdd.n7080 0.002
R51606 vdd.n7071 vdd.n7070 0.002
R51607 vdd.n7073 vdd.n7072 0.002
R51608 vdd.n7063 vdd.n7062 0.002
R51609 vdd.n7065 vdd.n7064 0.002
R51610 vdd.n7055 vdd.n7054 0.002
R51611 vdd.n7057 vdd.n7056 0.002
R51612 vdd.n7047 vdd.n7046 0.002
R51613 vdd.n7049 vdd.n7048 0.002
R51614 vdd.n7039 vdd.n7038 0.002
R51615 vdd.n7041 vdd.n7040 0.002
R51616 vdd.n7031 vdd.n7030 0.002
R51617 vdd.n7033 vdd.n7032 0.002
R51618 vdd.n7023 vdd.n7022 0.002
R51619 vdd.n7025 vdd.n7024 0.002
R51620 vdd.n7190 vdd.n7189 0.002
R51621 vdd.n7192 vdd.n7191 0.002
R51622 vdd.n7339 vdd.n7338 0.002
R51623 vdd.n7341 vdd.n7340 0.002
R51624 vdd.n7331 vdd.n7330 0.002
R51625 vdd.n7333 vdd.n7332 0.002
R51626 vdd.n7323 vdd.n7322 0.002
R51627 vdd.n7325 vdd.n7324 0.002
R51628 vdd.n7315 vdd.n7314 0.002
R51629 vdd.n7317 vdd.n7316 0.002
R51630 vdd.n7307 vdd.n7306 0.002
R51631 vdd.n7309 vdd.n7308 0.002
R51632 vdd.n7299 vdd.n7298 0.002
R51633 vdd.n7301 vdd.n7300 0.002
R51634 vdd.n7291 vdd.n7290 0.002
R51635 vdd.n7293 vdd.n7292 0.002
R51636 vdd.n7283 vdd.n7282 0.002
R51637 vdd.n7285 vdd.n7284 0.002
R51638 vdd.n7275 vdd.n7274 0.002
R51639 vdd.n7277 vdd.n7276 0.002
R51640 vdd.n7259 vdd.n7258 0.002
R51641 vdd.n7261 vdd.n7260 0.002
R51642 vdd.n7251 vdd.n7250 0.002
R51643 vdd.n7253 vdd.n7252 0.002
R51644 vdd.n7243 vdd.n7242 0.002
R51645 vdd.n7245 vdd.n7244 0.002
R51646 vdd.n7235 vdd.n7234 0.002
R51647 vdd.n7237 vdd.n7236 0.002
R51648 vdd.n7227 vdd.n7226 0.002
R51649 vdd.n7229 vdd.n7228 0.002
R51650 vdd.n7219 vdd.n7218 0.002
R51651 vdd.n7221 vdd.n7220 0.002
R51652 vdd.n7211 vdd.n7210 0.002
R51653 vdd.n7213 vdd.n7212 0.002
R51654 vdd.n7203 vdd.n7202 0.002
R51655 vdd.n7205 vdd.n7204 0.002
R51656 vdd.n7370 vdd.n7369 0.002
R51657 vdd.n7372 vdd.n7371 0.002
R51658 vdd.n7519 vdd.n7518 0.002
R51659 vdd.n7521 vdd.n7520 0.002
R51660 vdd.n7511 vdd.n7510 0.002
R51661 vdd.n7513 vdd.n7512 0.002
R51662 vdd.n7503 vdd.n7502 0.002
R51663 vdd.n7505 vdd.n7504 0.002
R51664 vdd.n7495 vdd.n7494 0.002
R51665 vdd.n7497 vdd.n7496 0.002
R51666 vdd.n7487 vdd.n7486 0.002
R51667 vdd.n7489 vdd.n7488 0.002
R51668 vdd.n7479 vdd.n7478 0.002
R51669 vdd.n7481 vdd.n7480 0.002
R51670 vdd.n7471 vdd.n7470 0.002
R51671 vdd.n7473 vdd.n7472 0.002
R51672 vdd.n7463 vdd.n7462 0.002
R51673 vdd.n7465 vdd.n7464 0.002
R51674 vdd.n7455 vdd.n7454 0.002
R51675 vdd.n7457 vdd.n7456 0.002
R51676 vdd.n7439 vdd.n7438 0.002
R51677 vdd.n7441 vdd.n7440 0.002
R51678 vdd.n7431 vdd.n7430 0.002
R51679 vdd.n7433 vdd.n7432 0.002
R51680 vdd.n7423 vdd.n7422 0.002
R51681 vdd.n7425 vdd.n7424 0.002
R51682 vdd.n7415 vdd.n7414 0.002
R51683 vdd.n7417 vdd.n7416 0.002
R51684 vdd.n7407 vdd.n7406 0.002
R51685 vdd.n7409 vdd.n7408 0.002
R51686 vdd.n7399 vdd.n7398 0.002
R51687 vdd.n7401 vdd.n7400 0.002
R51688 vdd.n7391 vdd.n7390 0.002
R51689 vdd.n7393 vdd.n7392 0.002
R51690 vdd.n7383 vdd.n7382 0.002
R51691 vdd.n7385 vdd.n7384 0.002
R51692 vdd.n7550 vdd.n7549 0.002
R51693 vdd.n7552 vdd.n7551 0.002
R51694 vdd.n7699 vdd.n7698 0.002
R51695 vdd.n7701 vdd.n7700 0.002
R51696 vdd.n7691 vdd.n7690 0.002
R51697 vdd.n7693 vdd.n7692 0.002
R51698 vdd.n7683 vdd.n7682 0.002
R51699 vdd.n7685 vdd.n7684 0.002
R51700 vdd.n7675 vdd.n7674 0.002
R51701 vdd.n7677 vdd.n7676 0.002
R51702 vdd.n7667 vdd.n7666 0.002
R51703 vdd.n7669 vdd.n7668 0.002
R51704 vdd.n7659 vdd.n7658 0.002
R51705 vdd.n7661 vdd.n7660 0.002
R51706 vdd.n7651 vdd.n7650 0.002
R51707 vdd.n7653 vdd.n7652 0.002
R51708 vdd.n7643 vdd.n7642 0.002
R51709 vdd.n7645 vdd.n7644 0.002
R51710 vdd.n7635 vdd.n7634 0.002
R51711 vdd.n7637 vdd.n7636 0.002
R51712 vdd.n7619 vdd.n7618 0.002
R51713 vdd.n7621 vdd.n7620 0.002
R51714 vdd.n7611 vdd.n7610 0.002
R51715 vdd.n7613 vdd.n7612 0.002
R51716 vdd.n7603 vdd.n7602 0.002
R51717 vdd.n7605 vdd.n7604 0.002
R51718 vdd.n7595 vdd.n7594 0.002
R51719 vdd.n7597 vdd.n7596 0.002
R51720 vdd.n7587 vdd.n7586 0.002
R51721 vdd.n7589 vdd.n7588 0.002
R51722 vdd.n7579 vdd.n7578 0.002
R51723 vdd.n7581 vdd.n7580 0.002
R51724 vdd.n7571 vdd.n7570 0.002
R51725 vdd.n7573 vdd.n7572 0.002
R51726 vdd.n7563 vdd.n7562 0.002
R51727 vdd.n7565 vdd.n7564 0.002
R51728 vdd.n7730 vdd.n7729 0.002
R51729 vdd.n7732 vdd.n7731 0.002
R51730 vdd.n7879 vdd.n7878 0.002
R51731 vdd.n7881 vdd.n7880 0.002
R51732 vdd.n7871 vdd.n7870 0.002
R51733 vdd.n7873 vdd.n7872 0.002
R51734 vdd.n7863 vdd.n7862 0.002
R51735 vdd.n7865 vdd.n7864 0.002
R51736 vdd.n7855 vdd.n7854 0.002
R51737 vdd.n7857 vdd.n7856 0.002
R51738 vdd.n7847 vdd.n7846 0.002
R51739 vdd.n7849 vdd.n7848 0.002
R51740 vdd.n7839 vdd.n7838 0.002
R51741 vdd.n7841 vdd.n7840 0.002
R51742 vdd.n7831 vdd.n7830 0.002
R51743 vdd.n7833 vdd.n7832 0.002
R51744 vdd.n7823 vdd.n7822 0.002
R51745 vdd.n7825 vdd.n7824 0.002
R51746 vdd.n7815 vdd.n7814 0.002
R51747 vdd.n7817 vdd.n7816 0.002
R51748 vdd.n7799 vdd.n7798 0.002
R51749 vdd.n7801 vdd.n7800 0.002
R51750 vdd.n7791 vdd.n7790 0.002
R51751 vdd.n7793 vdd.n7792 0.002
R51752 vdd.n7783 vdd.n7782 0.002
R51753 vdd.n7785 vdd.n7784 0.002
R51754 vdd.n7775 vdd.n7774 0.002
R51755 vdd.n7777 vdd.n7776 0.002
R51756 vdd.n7767 vdd.n7766 0.002
R51757 vdd.n7769 vdd.n7768 0.002
R51758 vdd.n7759 vdd.n7758 0.002
R51759 vdd.n7761 vdd.n7760 0.002
R51760 vdd.n7751 vdd.n7750 0.002
R51761 vdd.n7753 vdd.n7752 0.002
R51762 vdd.n7743 vdd.n7742 0.002
R51763 vdd.n7745 vdd.n7744 0.002
R51764 vdd.n7910 vdd.n7909 0.002
R51765 vdd.n7912 vdd.n7911 0.002
R51766 vdd.n8059 vdd.n8058 0.002
R51767 vdd.n8061 vdd.n8060 0.002
R51768 vdd.n8051 vdd.n8050 0.002
R51769 vdd.n8053 vdd.n8052 0.002
R51770 vdd.n8043 vdd.n8042 0.002
R51771 vdd.n8045 vdd.n8044 0.002
R51772 vdd.n8035 vdd.n8034 0.002
R51773 vdd.n8037 vdd.n8036 0.002
R51774 vdd.n8027 vdd.n8026 0.002
R51775 vdd.n8029 vdd.n8028 0.002
R51776 vdd.n8019 vdd.n8018 0.002
R51777 vdd.n8021 vdd.n8020 0.002
R51778 vdd.n8011 vdd.n8010 0.002
R51779 vdd.n8013 vdd.n8012 0.002
R51780 vdd.n8003 vdd.n8002 0.002
R51781 vdd.n8005 vdd.n8004 0.002
R51782 vdd.n7995 vdd.n7994 0.002
R51783 vdd.n7997 vdd.n7996 0.002
R51784 vdd.n7979 vdd.n7978 0.002
R51785 vdd.n7981 vdd.n7980 0.002
R51786 vdd.n7971 vdd.n7970 0.002
R51787 vdd.n7973 vdd.n7972 0.002
R51788 vdd.n7963 vdd.n7962 0.002
R51789 vdd.n7965 vdd.n7964 0.002
R51790 vdd.n7955 vdd.n7954 0.002
R51791 vdd.n7957 vdd.n7956 0.002
R51792 vdd.n7947 vdd.n7946 0.002
R51793 vdd.n7949 vdd.n7948 0.002
R51794 vdd.n7939 vdd.n7938 0.002
R51795 vdd.n7941 vdd.n7940 0.002
R51796 vdd.n7931 vdd.n7930 0.002
R51797 vdd.n7933 vdd.n7932 0.002
R51798 vdd.n7923 vdd.n7922 0.002
R51799 vdd.n7925 vdd.n7924 0.002
R51800 vdd.n8090 vdd.n8089 0.002
R51801 vdd.n8092 vdd.n8091 0.002
R51802 vdd.n8239 vdd.n8238 0.002
R51803 vdd.n8241 vdd.n8240 0.002
R51804 vdd.n8231 vdd.n8230 0.002
R51805 vdd.n8233 vdd.n8232 0.002
R51806 vdd.n8223 vdd.n8222 0.002
R51807 vdd.n8225 vdd.n8224 0.002
R51808 vdd.n8215 vdd.n8214 0.002
R51809 vdd.n8217 vdd.n8216 0.002
R51810 vdd.n8207 vdd.n8206 0.002
R51811 vdd.n8209 vdd.n8208 0.002
R51812 vdd.n8199 vdd.n8198 0.002
R51813 vdd.n8201 vdd.n8200 0.002
R51814 vdd.n8191 vdd.n8190 0.002
R51815 vdd.n8193 vdd.n8192 0.002
R51816 vdd.n8183 vdd.n8182 0.002
R51817 vdd.n8185 vdd.n8184 0.002
R51818 vdd.n8175 vdd.n8174 0.002
R51819 vdd.n8177 vdd.n8176 0.002
R51820 vdd.n8159 vdd.n8158 0.002
R51821 vdd.n8161 vdd.n8160 0.002
R51822 vdd.n8151 vdd.n8150 0.002
R51823 vdd.n8153 vdd.n8152 0.002
R51824 vdd.n8143 vdd.n8142 0.002
R51825 vdd.n8145 vdd.n8144 0.002
R51826 vdd.n8135 vdd.n8134 0.002
R51827 vdd.n8137 vdd.n8136 0.002
R51828 vdd.n8127 vdd.n8126 0.002
R51829 vdd.n8129 vdd.n8128 0.002
R51830 vdd.n8119 vdd.n8118 0.002
R51831 vdd.n8121 vdd.n8120 0.002
R51832 vdd.n8111 vdd.n8110 0.002
R51833 vdd.n8113 vdd.n8112 0.002
R51834 vdd.n8103 vdd.n8102 0.002
R51835 vdd.n8105 vdd.n8104 0.002
R51836 vdd.n8270 vdd.n8269 0.002
R51837 vdd.n8272 vdd.n8271 0.002
R51838 vdd.n8419 vdd.n8418 0.002
R51839 vdd.n8421 vdd.n8420 0.002
R51840 vdd.n8411 vdd.n8410 0.002
R51841 vdd.n8413 vdd.n8412 0.002
R51842 vdd.n8403 vdd.n8402 0.002
R51843 vdd.n8405 vdd.n8404 0.002
R51844 vdd.n8395 vdd.n8394 0.002
R51845 vdd.n8397 vdd.n8396 0.002
R51846 vdd.n8387 vdd.n8386 0.002
R51847 vdd.n8389 vdd.n8388 0.002
R51848 vdd.n8379 vdd.n8378 0.002
R51849 vdd.n8381 vdd.n8380 0.002
R51850 vdd.n8371 vdd.n8370 0.002
R51851 vdd.n8373 vdd.n8372 0.002
R51852 vdd.n8363 vdd.n8362 0.002
R51853 vdd.n8365 vdd.n8364 0.002
R51854 vdd.n8355 vdd.n8354 0.002
R51855 vdd.n8357 vdd.n8356 0.002
R51856 vdd.n8339 vdd.n8338 0.002
R51857 vdd.n8341 vdd.n8340 0.002
R51858 vdd.n8331 vdd.n8330 0.002
R51859 vdd.n8333 vdd.n8332 0.002
R51860 vdd.n8323 vdd.n8322 0.002
R51861 vdd.n8325 vdd.n8324 0.002
R51862 vdd.n8315 vdd.n8314 0.002
R51863 vdd.n8317 vdd.n8316 0.002
R51864 vdd.n8307 vdd.n8306 0.002
R51865 vdd.n8309 vdd.n8308 0.002
R51866 vdd.n8299 vdd.n8298 0.002
R51867 vdd.n8301 vdd.n8300 0.002
R51868 vdd.n8291 vdd.n8290 0.002
R51869 vdd.n8293 vdd.n8292 0.002
R51870 vdd.n8283 vdd.n8282 0.002
R51871 vdd.n8285 vdd.n8284 0.002
R51872 vdd.n8450 vdd.n8449 0.002
R51873 vdd.n8452 vdd.n8451 0.002
R51874 vdd.n8599 vdd.n8598 0.002
R51875 vdd.n8601 vdd.n8600 0.002
R51876 vdd.n8591 vdd.n8590 0.002
R51877 vdd.n8593 vdd.n8592 0.002
R51878 vdd.n8583 vdd.n8582 0.002
R51879 vdd.n8585 vdd.n8584 0.002
R51880 vdd.n8575 vdd.n8574 0.002
R51881 vdd.n8577 vdd.n8576 0.002
R51882 vdd.n8567 vdd.n8566 0.002
R51883 vdd.n8569 vdd.n8568 0.002
R51884 vdd.n8559 vdd.n8558 0.002
R51885 vdd.n8561 vdd.n8560 0.002
R51886 vdd.n8551 vdd.n8550 0.002
R51887 vdd.n8553 vdd.n8552 0.002
R51888 vdd.n8543 vdd.n8542 0.002
R51889 vdd.n8545 vdd.n8544 0.002
R51890 vdd.n8535 vdd.n8534 0.002
R51891 vdd.n8537 vdd.n8536 0.002
R51892 vdd.n8519 vdd.n8518 0.002
R51893 vdd.n8521 vdd.n8520 0.002
R51894 vdd.n8511 vdd.n8510 0.002
R51895 vdd.n8513 vdd.n8512 0.002
R51896 vdd.n8503 vdd.n8502 0.002
R51897 vdd.n8505 vdd.n8504 0.002
R51898 vdd.n8495 vdd.n8494 0.002
R51899 vdd.n8497 vdd.n8496 0.002
R51900 vdd.n8487 vdd.n8486 0.002
R51901 vdd.n8489 vdd.n8488 0.002
R51902 vdd.n8479 vdd.n8478 0.002
R51903 vdd.n8481 vdd.n8480 0.002
R51904 vdd.n8471 vdd.n8470 0.002
R51905 vdd.n8473 vdd.n8472 0.002
R51906 vdd.n8463 vdd.n8462 0.002
R51907 vdd.n8465 vdd.n8464 0.002
R51908 vdd.n8630 vdd.n8629 0.002
R51909 vdd.n8632 vdd.n8631 0.002
R51910 vdd.n8779 vdd.n8778 0.002
R51911 vdd.n8781 vdd.n8780 0.002
R51912 vdd.n8771 vdd.n8770 0.002
R51913 vdd.n8773 vdd.n8772 0.002
R51914 vdd.n8763 vdd.n8762 0.002
R51915 vdd.n8765 vdd.n8764 0.002
R51916 vdd.n8755 vdd.n8754 0.002
R51917 vdd.n8757 vdd.n8756 0.002
R51918 vdd.n8747 vdd.n8746 0.002
R51919 vdd.n8749 vdd.n8748 0.002
R51920 vdd.n8739 vdd.n8738 0.002
R51921 vdd.n8741 vdd.n8740 0.002
R51922 vdd.n8731 vdd.n8730 0.002
R51923 vdd.n8733 vdd.n8732 0.002
R51924 vdd.n8723 vdd.n8722 0.002
R51925 vdd.n8725 vdd.n8724 0.002
R51926 vdd.n8715 vdd.n8714 0.002
R51927 vdd.n8717 vdd.n8716 0.002
R51928 vdd.n8699 vdd.n8698 0.002
R51929 vdd.n8701 vdd.n8700 0.002
R51930 vdd.n8691 vdd.n8690 0.002
R51931 vdd.n8693 vdd.n8692 0.002
R51932 vdd.n8683 vdd.n8682 0.002
R51933 vdd.n8685 vdd.n8684 0.002
R51934 vdd.n8675 vdd.n8674 0.002
R51935 vdd.n8677 vdd.n8676 0.002
R51936 vdd.n8667 vdd.n8666 0.002
R51937 vdd.n8669 vdd.n8668 0.002
R51938 vdd.n8659 vdd.n8658 0.002
R51939 vdd.n8661 vdd.n8660 0.002
R51940 vdd.n8651 vdd.n8650 0.002
R51941 vdd.n8653 vdd.n8652 0.002
R51942 vdd.n8643 vdd.n8642 0.002
R51943 vdd.n8645 vdd.n8644 0.002
R51944 vdd.n8810 vdd.n8809 0.002
R51945 vdd.n8812 vdd.n8811 0.002
R51946 vdd.n8959 vdd.n8958 0.002
R51947 vdd.n8961 vdd.n8960 0.002
R51948 vdd.n8951 vdd.n8950 0.002
R51949 vdd.n8953 vdd.n8952 0.002
R51950 vdd.n8943 vdd.n8942 0.002
R51951 vdd.n8945 vdd.n8944 0.002
R51952 vdd.n8935 vdd.n8934 0.002
R51953 vdd.n8937 vdd.n8936 0.002
R51954 vdd.n8927 vdd.n8926 0.002
R51955 vdd.n8929 vdd.n8928 0.002
R51956 vdd.n8919 vdd.n8918 0.002
R51957 vdd.n8921 vdd.n8920 0.002
R51958 vdd.n8911 vdd.n8910 0.002
R51959 vdd.n8913 vdd.n8912 0.002
R51960 vdd.n8903 vdd.n8902 0.002
R51961 vdd.n8905 vdd.n8904 0.002
R51962 vdd.n8895 vdd.n8894 0.002
R51963 vdd.n8897 vdd.n8896 0.002
R51964 vdd.n8879 vdd.n8878 0.002
R51965 vdd.n8881 vdd.n8880 0.002
R51966 vdd.n8871 vdd.n8870 0.002
R51967 vdd.n8873 vdd.n8872 0.002
R51968 vdd.n8863 vdd.n8862 0.002
R51969 vdd.n8865 vdd.n8864 0.002
R51970 vdd.n8855 vdd.n8854 0.002
R51971 vdd.n8857 vdd.n8856 0.002
R51972 vdd.n8847 vdd.n8846 0.002
R51973 vdd.n8849 vdd.n8848 0.002
R51974 vdd.n8839 vdd.n8838 0.002
R51975 vdd.n8841 vdd.n8840 0.002
R51976 vdd.n8831 vdd.n8830 0.002
R51977 vdd.n8833 vdd.n8832 0.002
R51978 vdd.n8823 vdd.n8822 0.002
R51979 vdd.n8825 vdd.n8824 0.002
R51980 vdd.n8990 vdd.n8989 0.002
R51981 vdd.n8992 vdd.n8991 0.002
R51982 vdd.n9139 vdd.n9138 0.002
R51983 vdd.n9141 vdd.n9140 0.002
R51984 vdd.n9131 vdd.n9130 0.002
R51985 vdd.n9133 vdd.n9132 0.002
R51986 vdd.n9123 vdd.n9122 0.002
R51987 vdd.n9125 vdd.n9124 0.002
R51988 vdd.n9115 vdd.n9114 0.002
R51989 vdd.n9117 vdd.n9116 0.002
R51990 vdd.n9107 vdd.n9106 0.002
R51991 vdd.n9109 vdd.n9108 0.002
R51992 vdd.n9099 vdd.n9098 0.002
R51993 vdd.n9101 vdd.n9100 0.002
R51994 vdd.n9091 vdd.n9090 0.002
R51995 vdd.n9093 vdd.n9092 0.002
R51996 vdd.n9083 vdd.n9082 0.002
R51997 vdd.n9085 vdd.n9084 0.002
R51998 vdd.n9075 vdd.n9074 0.002
R51999 vdd.n9077 vdd.n9076 0.002
R52000 vdd.n9059 vdd.n9058 0.002
R52001 vdd.n9061 vdd.n9060 0.002
R52002 vdd.n9051 vdd.n9050 0.002
R52003 vdd.n9053 vdd.n9052 0.002
R52004 vdd.n9043 vdd.n9042 0.002
R52005 vdd.n9045 vdd.n9044 0.002
R52006 vdd.n9035 vdd.n9034 0.002
R52007 vdd.n9037 vdd.n9036 0.002
R52008 vdd.n9027 vdd.n9026 0.002
R52009 vdd.n9029 vdd.n9028 0.002
R52010 vdd.n9019 vdd.n9018 0.002
R52011 vdd.n9021 vdd.n9020 0.002
R52012 vdd.n9011 vdd.n9010 0.002
R52013 vdd.n9013 vdd.n9012 0.002
R52014 vdd.n9003 vdd.n9002 0.002
R52015 vdd.n9005 vdd.n9004 0.002
R52016 vdd.n9170 vdd.n9169 0.002
R52017 vdd.n9172 vdd.n9171 0.002
R52018 vdd.n9319 vdd.n9318 0.002
R52019 vdd.n9321 vdd.n9320 0.002
R52020 vdd.n9311 vdd.n9310 0.002
R52021 vdd.n9313 vdd.n9312 0.002
R52022 vdd.n9303 vdd.n9302 0.002
R52023 vdd.n9305 vdd.n9304 0.002
R52024 vdd.n9295 vdd.n9294 0.002
R52025 vdd.n9297 vdd.n9296 0.002
R52026 vdd.n9287 vdd.n9286 0.002
R52027 vdd.n9289 vdd.n9288 0.002
R52028 vdd.n9279 vdd.n9278 0.002
R52029 vdd.n9281 vdd.n9280 0.002
R52030 vdd.n9271 vdd.n9270 0.002
R52031 vdd.n9273 vdd.n9272 0.002
R52032 vdd.n9263 vdd.n9262 0.002
R52033 vdd.n9265 vdd.n9264 0.002
R52034 vdd.n9255 vdd.n9254 0.002
R52035 vdd.n9257 vdd.n9256 0.002
R52036 vdd.n9239 vdd.n9238 0.002
R52037 vdd.n9241 vdd.n9240 0.002
R52038 vdd.n9231 vdd.n9230 0.002
R52039 vdd.n9233 vdd.n9232 0.002
R52040 vdd.n9223 vdd.n9222 0.002
R52041 vdd.n9225 vdd.n9224 0.002
R52042 vdd.n9215 vdd.n9214 0.002
R52043 vdd.n9217 vdd.n9216 0.002
R52044 vdd.n9207 vdd.n9206 0.002
R52045 vdd.n9209 vdd.n9208 0.002
R52046 vdd.n9199 vdd.n9198 0.002
R52047 vdd.n9201 vdd.n9200 0.002
R52048 vdd.n9191 vdd.n9190 0.002
R52049 vdd.n9193 vdd.n9192 0.002
R52050 vdd.n9183 vdd.n9182 0.002
R52051 vdd.n9185 vdd.n9184 0.002
R52052 vdd.n9350 vdd.n9349 0.002
R52053 vdd.n9352 vdd.n9351 0.002
R52054 vdd.n9499 vdd.n9498 0.002
R52055 vdd.n9501 vdd.n9500 0.002
R52056 vdd.n9491 vdd.n9490 0.002
R52057 vdd.n9493 vdd.n9492 0.002
R52058 vdd.n9483 vdd.n9482 0.002
R52059 vdd.n9485 vdd.n9484 0.002
R52060 vdd.n9475 vdd.n9474 0.002
R52061 vdd.n9477 vdd.n9476 0.002
R52062 vdd.n9467 vdd.n9466 0.002
R52063 vdd.n9469 vdd.n9468 0.002
R52064 vdd.n9459 vdd.n9458 0.002
R52065 vdd.n9461 vdd.n9460 0.002
R52066 vdd.n9451 vdd.n9450 0.002
R52067 vdd.n9453 vdd.n9452 0.002
R52068 vdd.n9443 vdd.n9442 0.002
R52069 vdd.n9445 vdd.n9444 0.002
R52070 vdd.n9435 vdd.n9434 0.002
R52071 vdd.n9437 vdd.n9436 0.002
R52072 vdd.n9419 vdd.n9418 0.002
R52073 vdd.n9421 vdd.n9420 0.002
R52074 vdd.n9411 vdd.n9410 0.002
R52075 vdd.n9413 vdd.n9412 0.002
R52076 vdd.n9403 vdd.n9402 0.002
R52077 vdd.n9405 vdd.n9404 0.002
R52078 vdd.n9395 vdd.n9394 0.002
R52079 vdd.n9397 vdd.n9396 0.002
R52080 vdd.n9387 vdd.n9386 0.002
R52081 vdd.n9389 vdd.n9388 0.002
R52082 vdd.n9379 vdd.n9378 0.002
R52083 vdd.n9381 vdd.n9380 0.002
R52084 vdd.n9371 vdd.n9370 0.002
R52085 vdd.n9373 vdd.n9372 0.002
R52086 vdd.n9363 vdd.n9362 0.002
R52087 vdd.n9365 vdd.n9364 0.002
R52088 vdd.n9530 vdd.n9529 0.002
R52089 vdd.n9532 vdd.n9531 0.002
R52090 vdd.n9679 vdd.n9678 0.002
R52091 vdd.n9681 vdd.n9680 0.002
R52092 vdd.n9671 vdd.n9670 0.002
R52093 vdd.n9673 vdd.n9672 0.002
R52094 vdd.n9663 vdd.n9662 0.002
R52095 vdd.n9665 vdd.n9664 0.002
R52096 vdd.n9655 vdd.n9654 0.002
R52097 vdd.n9657 vdd.n9656 0.002
R52098 vdd.n9647 vdd.n9646 0.002
R52099 vdd.n9649 vdd.n9648 0.002
R52100 vdd.n9639 vdd.n9638 0.002
R52101 vdd.n9641 vdd.n9640 0.002
R52102 vdd.n9631 vdd.n9630 0.002
R52103 vdd.n9633 vdd.n9632 0.002
R52104 vdd.n9623 vdd.n9622 0.002
R52105 vdd.n9625 vdd.n9624 0.002
R52106 vdd.n9615 vdd.n9614 0.002
R52107 vdd.n9617 vdd.n9616 0.002
R52108 vdd.n9599 vdd.n9598 0.002
R52109 vdd.n9601 vdd.n9600 0.002
R52110 vdd.n9591 vdd.n9590 0.002
R52111 vdd.n9593 vdd.n9592 0.002
R52112 vdd.n9583 vdd.n9582 0.002
R52113 vdd.n9585 vdd.n9584 0.002
R52114 vdd.n9575 vdd.n9574 0.002
R52115 vdd.n9577 vdd.n9576 0.002
R52116 vdd.n9567 vdd.n9566 0.002
R52117 vdd.n9569 vdd.n9568 0.002
R52118 vdd.n9559 vdd.n9558 0.002
R52119 vdd.n9561 vdd.n9560 0.002
R52120 vdd.n9551 vdd.n9550 0.002
R52121 vdd.n9553 vdd.n9552 0.002
R52122 vdd.n9543 vdd.n9542 0.002
R52123 vdd.n9545 vdd.n9544 0.002
R52124 vdd.n9710 vdd.n9709 0.002
R52125 vdd.n9712 vdd.n9711 0.002
R52126 vdd.n9859 vdd.n9858 0.002
R52127 vdd.n9861 vdd.n9860 0.002
R52128 vdd.n9851 vdd.n9850 0.002
R52129 vdd.n9853 vdd.n9852 0.002
R52130 vdd.n9843 vdd.n9842 0.002
R52131 vdd.n9845 vdd.n9844 0.002
R52132 vdd.n9835 vdd.n9834 0.002
R52133 vdd.n9837 vdd.n9836 0.002
R52134 vdd.n9827 vdd.n9826 0.002
R52135 vdd.n9829 vdd.n9828 0.002
R52136 vdd.n9819 vdd.n9818 0.002
R52137 vdd.n9821 vdd.n9820 0.002
R52138 vdd.n9811 vdd.n9810 0.002
R52139 vdd.n9813 vdd.n9812 0.002
R52140 vdd.n9803 vdd.n9802 0.002
R52141 vdd.n9805 vdd.n9804 0.002
R52142 vdd.n9795 vdd.n9794 0.002
R52143 vdd.n9797 vdd.n9796 0.002
R52144 vdd.n9779 vdd.n9778 0.002
R52145 vdd.n9781 vdd.n9780 0.002
R52146 vdd.n9771 vdd.n9770 0.002
R52147 vdd.n9773 vdd.n9772 0.002
R52148 vdd.n9763 vdd.n9762 0.002
R52149 vdd.n9765 vdd.n9764 0.002
R52150 vdd.n9755 vdd.n9754 0.002
R52151 vdd.n9757 vdd.n9756 0.002
R52152 vdd.n9747 vdd.n9746 0.002
R52153 vdd.n9749 vdd.n9748 0.002
R52154 vdd.n9739 vdd.n9738 0.002
R52155 vdd.n9741 vdd.n9740 0.002
R52156 vdd.n9731 vdd.n9730 0.002
R52157 vdd.n9733 vdd.n9732 0.002
R52158 vdd.n9723 vdd.n9722 0.002
R52159 vdd.n9725 vdd.n9724 0.002
R52160 vdd.n9890 vdd.n9889 0.002
R52161 vdd.n9892 vdd.n9891 0.002
R52162 vdd.n10039 vdd.n10038 0.002
R52163 vdd.n10041 vdd.n10040 0.002
R52164 vdd.n10031 vdd.n10030 0.002
R52165 vdd.n10033 vdd.n10032 0.002
R52166 vdd.n10023 vdd.n10022 0.002
R52167 vdd.n10025 vdd.n10024 0.002
R52168 vdd.n10015 vdd.n10014 0.002
R52169 vdd.n10017 vdd.n10016 0.002
R52170 vdd.n10007 vdd.n10006 0.002
R52171 vdd.n10009 vdd.n10008 0.002
R52172 vdd.n9999 vdd.n9998 0.002
R52173 vdd.n10001 vdd.n10000 0.002
R52174 vdd.n9991 vdd.n9990 0.002
R52175 vdd.n9993 vdd.n9992 0.002
R52176 vdd.n9983 vdd.n9982 0.002
R52177 vdd.n9985 vdd.n9984 0.002
R52178 vdd.n9975 vdd.n9974 0.002
R52179 vdd.n9977 vdd.n9976 0.002
R52180 vdd.n9959 vdd.n9958 0.002
R52181 vdd.n9961 vdd.n9960 0.002
R52182 vdd.n9951 vdd.n9950 0.002
R52183 vdd.n9953 vdd.n9952 0.002
R52184 vdd.n9943 vdd.n9942 0.002
R52185 vdd.n9945 vdd.n9944 0.002
R52186 vdd.n9935 vdd.n9934 0.002
R52187 vdd.n9937 vdd.n9936 0.002
R52188 vdd.n9927 vdd.n9926 0.002
R52189 vdd.n9929 vdd.n9928 0.002
R52190 vdd.n9919 vdd.n9918 0.002
R52191 vdd.n9921 vdd.n9920 0.002
R52192 vdd.n9911 vdd.n9910 0.002
R52193 vdd.n9913 vdd.n9912 0.002
R52194 vdd.n9903 vdd.n9902 0.002
R52195 vdd.n9905 vdd.n9904 0.002
R52196 vdd.n10070 vdd.n10069 0.002
R52197 vdd.n10072 vdd.n10071 0.002
R52198 vdd.n10219 vdd.n10218 0.002
R52199 vdd.n10221 vdd.n10220 0.002
R52200 vdd.n10211 vdd.n10210 0.002
R52201 vdd.n10213 vdd.n10212 0.002
R52202 vdd.n10203 vdd.n10202 0.002
R52203 vdd.n10205 vdd.n10204 0.002
R52204 vdd.n10195 vdd.n10194 0.002
R52205 vdd.n10197 vdd.n10196 0.002
R52206 vdd.n10187 vdd.n10186 0.002
R52207 vdd.n10189 vdd.n10188 0.002
R52208 vdd.n10179 vdd.n10178 0.002
R52209 vdd.n10181 vdd.n10180 0.002
R52210 vdd.n10171 vdd.n10170 0.002
R52211 vdd.n10173 vdd.n10172 0.002
R52212 vdd.n10163 vdd.n10162 0.002
R52213 vdd.n10165 vdd.n10164 0.002
R52214 vdd.n10155 vdd.n10154 0.002
R52215 vdd.n10157 vdd.n10156 0.002
R52216 vdd.n10139 vdd.n10138 0.002
R52217 vdd.n10141 vdd.n10140 0.002
R52218 vdd.n10131 vdd.n10130 0.002
R52219 vdd.n10133 vdd.n10132 0.002
R52220 vdd.n10123 vdd.n10122 0.002
R52221 vdd.n10125 vdd.n10124 0.002
R52222 vdd.n10115 vdd.n10114 0.002
R52223 vdd.n10117 vdd.n10116 0.002
R52224 vdd.n10107 vdd.n10106 0.002
R52225 vdd.n10109 vdd.n10108 0.002
R52226 vdd.n10099 vdd.n10098 0.002
R52227 vdd.n10101 vdd.n10100 0.002
R52228 vdd.n10091 vdd.n10090 0.002
R52229 vdd.n10093 vdd.n10092 0.002
R52230 vdd.n10083 vdd.n10082 0.002
R52231 vdd.n10085 vdd.n10084 0.002
R52232 vdd.n10250 vdd.n10249 0.002
R52233 vdd.n10252 vdd.n10251 0.002
R52234 vdd.n10399 vdd.n10398 0.002
R52235 vdd.n10401 vdd.n10400 0.002
R52236 vdd.n10391 vdd.n10390 0.002
R52237 vdd.n10393 vdd.n10392 0.002
R52238 vdd.n10383 vdd.n10382 0.002
R52239 vdd.n10385 vdd.n10384 0.002
R52240 vdd.n10375 vdd.n10374 0.002
R52241 vdd.n10377 vdd.n10376 0.002
R52242 vdd.n10367 vdd.n10366 0.002
R52243 vdd.n10369 vdd.n10368 0.002
R52244 vdd.n10359 vdd.n10358 0.002
R52245 vdd.n10361 vdd.n10360 0.002
R52246 vdd.n10351 vdd.n10350 0.002
R52247 vdd.n10353 vdd.n10352 0.002
R52248 vdd.n10343 vdd.n10342 0.002
R52249 vdd.n10345 vdd.n10344 0.002
R52250 vdd.n10335 vdd.n10334 0.002
R52251 vdd.n10337 vdd.n10336 0.002
R52252 vdd.n10319 vdd.n10318 0.002
R52253 vdd.n10321 vdd.n10320 0.002
R52254 vdd.n10311 vdd.n10310 0.002
R52255 vdd.n10313 vdd.n10312 0.002
R52256 vdd.n10303 vdd.n10302 0.002
R52257 vdd.n10305 vdd.n10304 0.002
R52258 vdd.n10295 vdd.n10294 0.002
R52259 vdd.n10297 vdd.n10296 0.002
R52260 vdd.n10287 vdd.n10286 0.002
R52261 vdd.n10289 vdd.n10288 0.002
R52262 vdd.n10279 vdd.n10278 0.002
R52263 vdd.n10281 vdd.n10280 0.002
R52264 vdd.n10271 vdd.n10270 0.002
R52265 vdd.n10273 vdd.n10272 0.002
R52266 vdd.n10263 vdd.n10262 0.002
R52267 vdd.n10265 vdd.n10264 0.002
R52268 vdd.n10430 vdd.n10429 0.002
R52269 vdd.n10432 vdd.n10431 0.002
R52270 vdd.n10579 vdd.n10578 0.002
R52271 vdd.n10581 vdd.n10580 0.002
R52272 vdd.n10571 vdd.n10570 0.002
R52273 vdd.n10573 vdd.n10572 0.002
R52274 vdd.n10563 vdd.n10562 0.002
R52275 vdd.n10565 vdd.n10564 0.002
R52276 vdd.n10555 vdd.n10554 0.002
R52277 vdd.n10557 vdd.n10556 0.002
R52278 vdd.n10547 vdd.n10546 0.002
R52279 vdd.n10549 vdd.n10548 0.002
R52280 vdd.n10539 vdd.n10538 0.002
R52281 vdd.n10541 vdd.n10540 0.002
R52282 vdd.n10531 vdd.n10530 0.002
R52283 vdd.n10533 vdd.n10532 0.002
R52284 vdd.n10523 vdd.n10522 0.002
R52285 vdd.n10525 vdd.n10524 0.002
R52286 vdd.n10515 vdd.n10514 0.002
R52287 vdd.n10517 vdd.n10516 0.002
R52288 vdd.n10499 vdd.n10498 0.002
R52289 vdd.n10501 vdd.n10500 0.002
R52290 vdd.n10491 vdd.n10490 0.002
R52291 vdd.n10493 vdd.n10492 0.002
R52292 vdd.n10483 vdd.n10482 0.002
R52293 vdd.n10485 vdd.n10484 0.002
R52294 vdd.n10475 vdd.n10474 0.002
R52295 vdd.n10477 vdd.n10476 0.002
R52296 vdd.n10467 vdd.n10466 0.002
R52297 vdd.n10469 vdd.n10468 0.002
R52298 vdd.n10459 vdd.n10458 0.002
R52299 vdd.n10461 vdd.n10460 0.002
R52300 vdd.n10451 vdd.n10450 0.002
R52301 vdd.n10453 vdd.n10452 0.002
R52302 vdd.n10443 vdd.n10442 0.002
R52303 vdd.n10445 vdd.n10444 0.002
R52304 vdd.n10610 vdd.n10609 0.002
R52305 vdd.n10612 vdd.n10611 0.002
R52306 vdd.n10759 vdd.n10758 0.002
R52307 vdd.n10761 vdd.n10760 0.002
R52308 vdd.n10751 vdd.n10750 0.002
R52309 vdd.n10753 vdd.n10752 0.002
R52310 vdd.n10743 vdd.n10742 0.002
R52311 vdd.n10745 vdd.n10744 0.002
R52312 vdd.n10735 vdd.n10734 0.002
R52313 vdd.n10737 vdd.n10736 0.002
R52314 vdd.n10727 vdd.n10726 0.002
R52315 vdd.n10729 vdd.n10728 0.002
R52316 vdd.n10719 vdd.n10718 0.002
R52317 vdd.n10721 vdd.n10720 0.002
R52318 vdd.n10711 vdd.n10710 0.002
R52319 vdd.n10713 vdd.n10712 0.002
R52320 vdd.n10703 vdd.n10702 0.002
R52321 vdd.n10705 vdd.n10704 0.002
R52322 vdd.n10695 vdd.n10694 0.002
R52323 vdd.n10697 vdd.n10696 0.002
R52324 vdd.n10679 vdd.n10678 0.002
R52325 vdd.n10681 vdd.n10680 0.002
R52326 vdd.n10671 vdd.n10670 0.002
R52327 vdd.n10673 vdd.n10672 0.002
R52328 vdd.n10663 vdd.n10662 0.002
R52329 vdd.n10665 vdd.n10664 0.002
R52330 vdd.n10655 vdd.n10654 0.002
R52331 vdd.n10657 vdd.n10656 0.002
R52332 vdd.n10647 vdd.n10646 0.002
R52333 vdd.n10649 vdd.n10648 0.002
R52334 vdd.n10639 vdd.n10638 0.002
R52335 vdd.n10641 vdd.n10640 0.002
R52336 vdd.n10631 vdd.n10630 0.002
R52337 vdd.n10633 vdd.n10632 0.002
R52338 vdd.n10623 vdd.n10622 0.002
R52339 vdd.n10625 vdd.n10624 0.002
R52340 vdd.n10790 vdd.n10789 0.002
R52341 vdd.n10792 vdd.n10791 0.002
R52342 vdd.n10939 vdd.n10938 0.002
R52343 vdd.n10941 vdd.n10940 0.002
R52344 vdd.n10931 vdd.n10930 0.002
R52345 vdd.n10933 vdd.n10932 0.002
R52346 vdd.n10923 vdd.n10922 0.002
R52347 vdd.n10925 vdd.n10924 0.002
R52348 vdd.n10915 vdd.n10914 0.002
R52349 vdd.n10917 vdd.n10916 0.002
R52350 vdd.n10907 vdd.n10906 0.002
R52351 vdd.n10909 vdd.n10908 0.002
R52352 vdd.n10899 vdd.n10898 0.002
R52353 vdd.n10901 vdd.n10900 0.002
R52354 vdd.n10891 vdd.n10890 0.002
R52355 vdd.n10893 vdd.n10892 0.002
R52356 vdd.n10883 vdd.n10882 0.002
R52357 vdd.n10885 vdd.n10884 0.002
R52358 vdd.n10875 vdd.n10874 0.002
R52359 vdd.n10877 vdd.n10876 0.002
R52360 vdd.n10859 vdd.n10858 0.002
R52361 vdd.n10861 vdd.n10860 0.002
R52362 vdd.n10851 vdd.n10850 0.002
R52363 vdd.n10853 vdd.n10852 0.002
R52364 vdd.n10843 vdd.n10842 0.002
R52365 vdd.n10845 vdd.n10844 0.002
R52366 vdd.n10835 vdd.n10834 0.002
R52367 vdd.n10837 vdd.n10836 0.002
R52368 vdd.n10827 vdd.n10826 0.002
R52369 vdd.n10829 vdd.n10828 0.002
R52370 vdd.n10819 vdd.n10818 0.002
R52371 vdd.n10821 vdd.n10820 0.002
R52372 vdd.n10811 vdd.n10810 0.002
R52373 vdd.n10813 vdd.n10812 0.002
R52374 vdd.n10803 vdd.n10802 0.002
R52375 vdd.n10805 vdd.n10804 0.002
R52376 vdd.n10970 vdd.n10969 0.002
R52377 vdd.n10972 vdd.n10971 0.002
R52378 vdd.n11119 vdd.n11118 0.002
R52379 vdd.n11121 vdd.n11120 0.002
R52380 vdd.n11111 vdd.n11110 0.002
R52381 vdd.n11113 vdd.n11112 0.002
R52382 vdd.n11103 vdd.n11102 0.002
R52383 vdd.n11105 vdd.n11104 0.002
R52384 vdd.n11095 vdd.n11094 0.002
R52385 vdd.n11097 vdd.n11096 0.002
R52386 vdd.n11087 vdd.n11086 0.002
R52387 vdd.n11089 vdd.n11088 0.002
R52388 vdd.n11079 vdd.n11078 0.002
R52389 vdd.n11081 vdd.n11080 0.002
R52390 vdd.n11071 vdd.n11070 0.002
R52391 vdd.n11073 vdd.n11072 0.002
R52392 vdd.n11063 vdd.n11062 0.002
R52393 vdd.n11065 vdd.n11064 0.002
R52394 vdd.n11055 vdd.n11054 0.002
R52395 vdd.n11057 vdd.n11056 0.002
R52396 vdd.n11039 vdd.n11038 0.002
R52397 vdd.n11041 vdd.n11040 0.002
R52398 vdd.n11031 vdd.n11030 0.002
R52399 vdd.n11033 vdd.n11032 0.002
R52400 vdd.n11023 vdd.n11022 0.002
R52401 vdd.n11025 vdd.n11024 0.002
R52402 vdd.n11015 vdd.n11014 0.002
R52403 vdd.n11017 vdd.n11016 0.002
R52404 vdd.n11007 vdd.n11006 0.002
R52405 vdd.n11009 vdd.n11008 0.002
R52406 vdd.n10999 vdd.n10998 0.002
R52407 vdd.n11001 vdd.n11000 0.002
R52408 vdd.n10991 vdd.n10990 0.002
R52409 vdd.n10993 vdd.n10992 0.002
R52410 vdd.n10983 vdd.n10982 0.002
R52411 vdd.n10985 vdd.n10984 0.002
R52412 vdd.n11150 vdd.n11149 0.002
R52413 vdd.n11152 vdd.n11151 0.002
R52414 vdd.n11299 vdd.n11298 0.002
R52415 vdd.n11301 vdd.n11300 0.002
R52416 vdd.n11291 vdd.n11290 0.002
R52417 vdd.n11293 vdd.n11292 0.002
R52418 vdd.n11283 vdd.n11282 0.002
R52419 vdd.n11285 vdd.n11284 0.002
R52420 vdd.n11275 vdd.n11274 0.002
R52421 vdd.n11277 vdd.n11276 0.002
R52422 vdd.n11267 vdd.n11266 0.002
R52423 vdd.n11269 vdd.n11268 0.002
R52424 vdd.n11259 vdd.n11258 0.002
R52425 vdd.n11261 vdd.n11260 0.002
R52426 vdd.n11251 vdd.n11250 0.002
R52427 vdd.n11253 vdd.n11252 0.002
R52428 vdd.n11243 vdd.n11242 0.002
R52429 vdd.n11245 vdd.n11244 0.002
R52430 vdd.n11235 vdd.n11234 0.002
R52431 vdd.n11237 vdd.n11236 0.002
R52432 vdd.n11219 vdd.n11218 0.002
R52433 vdd.n11221 vdd.n11220 0.002
R52434 vdd.n11211 vdd.n11210 0.002
R52435 vdd.n11213 vdd.n11212 0.002
R52436 vdd.n11203 vdd.n11202 0.002
R52437 vdd.n11205 vdd.n11204 0.002
R52438 vdd.n11195 vdd.n11194 0.002
R52439 vdd.n11197 vdd.n11196 0.002
R52440 vdd.n11187 vdd.n11186 0.002
R52441 vdd.n11189 vdd.n11188 0.002
R52442 vdd.n11179 vdd.n11178 0.002
R52443 vdd.n11181 vdd.n11180 0.002
R52444 vdd.n11171 vdd.n11170 0.002
R52445 vdd.n11173 vdd.n11172 0.002
R52446 vdd.n11163 vdd.n11162 0.002
R52447 vdd.n11165 vdd.n11164 0.002
R52448 vdd.n11330 vdd.n11329 0.002
R52449 vdd.n11332 vdd.n11331 0.002
R52450 vdd vdd.n13545 0.002
R52451 vdd.n11387 vdd.n11348 0.001
R52452 vdd.n11386 vdd.n11385 0.001
R52453 vdd.n13506 vdd.n13467 0.001
R52454 vdd.n13505 vdd.n13504 0.001
R52455 vdd vdd.n11478 0.001
R52456 vdd.n11359 vdd.n11358 0.001
R52457 vdd.n11415 vdd.n11414 0.001
R52458 vdd.n13478 vdd.n13477 0.001
R52459 vdd.n13534 vdd.n13533 0.001
R52460 vp_n.n3043 vp_n.t19 702.112
R52461 vp_n.n1573 vp_n.t565 702.112
R52462 vp_n.n22 vp_n.t191 702.112
R52463 vp_n.n3229 vp_n.t396 702.112
R52464 vp_n.n3226 vp_n.t595 702.112
R52465 vp_n.n1583 vp_n.t450 702.112
R52466 vp_n.n32 vp_n.t109 702.112
R52467 vp_n.n3239 vp_n.t323 702.112
R52468 vp_n.n3236 vp_n.t518 702.112
R52469 vp_n.n1593 vp_n.t53 702.112
R52470 vp_n.n42 vp_n.t310 702.112
R52471 vp_n.n3249 vp_n.t524 702.112
R52472 vp_n.n3246 vp_n.t114 702.112
R52473 vp_n.n1603 vp_n.t176 702.112
R52474 vp_n.n52 vp_n.t398 702.112
R52475 vp_n.n3259 vp_n.t598 702.112
R52476 vp_n.n3256 vp_n.t196 702.112
R52477 vp_n.n1613 vp_n.t73 702.112
R52478 vp_n.n62 vp_n.t332 702.112
R52479 vp_n.n3269 vp_n.t544 702.112
R52480 vp_n.n3266 vp_n.t135 702.112
R52481 vp_n.n1623 vp_n.t66 702.112
R52482 vp_n.n72 vp_n.t327 702.112
R52483 vp_n.n3279 vp_n.t537 702.112
R52484 vp_n.n3276 vp_n.t129 702.112
R52485 vp_n.n1633 vp_n.t95 702.112
R52486 vp_n.n82 vp_n.t350 702.112
R52487 vp_n.n3289 vp_n.t558 702.112
R52488 vp_n.n3286 vp_n.t152 702.112
R52489 vp_n.n1643 vp_n.t303 702.112
R52490 vp_n.n92 vp_n.t548 702.112
R52491 vp_n.n3299 vp_n.t156 702.112
R52492 vp_n.n3296 vp_n.t354 702.112
R52493 vp_n.n1653 vp_n.t4 702.112
R52494 vp_n.n102 vp_n.t225 702.112
R52495 vp_n.n3309 vp_n.t434 702.112
R52496 vp_n.n3306 vp_n.t27 702.112
R52497 vp_n.n1663 vp_n.t319 702.112
R52498 vp_n.n112 vp_n.t563 702.112
R52499 vp_n.n3319 vp_n.t168 702.112
R52500 vp_n.n3316 vp_n.t367 702.112
R52501 vp_n.n1673 vp_n.t312 702.112
R52502 vp_n.n122 vp_n.t561 702.112
R52503 vp_n.n3329 vp_n.t164 702.112
R52504 vp_n.n3326 vp_n.t364 702.112
R52505 vp_n.n1683 vp_n.t209 702.112
R52506 vp_n.n132 vp_n.t442 702.112
R52507 vp_n.n3339 vp_n.t52 702.112
R52508 vp_n.n3336 vp_n.t248 702.112
R52509 vp_n.n1693 vp_n.t542 702.112
R52510 vp_n.n142 vp_n.t172 702.112
R52511 vp_n.n3349 vp_n.t383 702.112
R52512 vp_n.n3346 vp_n.t579 702.112
R52513 vp_n.n1703 vp_n.t218 702.112
R52514 vp_n.n152 vp_n.t463 702.112
R52515 vp_n.n3359 vp_n.t74 702.112
R52516 vp_n.n3356 vp_n.t270 702.112
R52517 vp_n.n1713 vp_n.t419 702.112
R52518 vp_n.n162 vp_n.t59 702.112
R52519 vp_n.n3369 vp_n.t281 702.112
R52520 vp_n.n3366 vp_n.t471 702.112
R52521 vp_n.n1723 vp_n.t525 702.112
R52522 vp_n.n172 vp_n.t162 702.112
R52523 vp_n.n3379 vp_n.t372 702.112
R52524 vp_n.n3376 vp_n.t567 702.112
R52525 vp_n.n1733 vp_n.t122 702.112
R52526 vp_n.n182 vp_n.t368 702.112
R52527 vp_n.n3389 vp_n.t574 702.112
R52528 vp_n.n3386 vp_n.t169 702.112
R52529 vp_n.n1743 vp_n.t330 702.112
R52530 vp_n.n192 vp_n.t566 702.112
R52531 vp_n.n3399 vp_n.t173 702.112
R52532 vp_n.n3396 vp_n.t371 702.112
R52533 vp_n.n1753 vp_n.t141 702.112
R52534 vp_n.n202 vp_n.t378 702.112
R52535 vp_n.n3409 vp_n.t585 702.112
R52536 vp_n.n3406 vp_n.t179 702.112
R52537 vp_n.n1763 vp_n.t348 702.112
R52538 vp_n.n212 vp_n.t580 702.112
R52539 vp_n.n3419 vp_n.t186 702.112
R52540 vp_n.n3416 vp_n.t384 702.112
R52541 vp_n.n1773 vp_n.t157 702.112
R52542 vp_n.n222 vp_n.t388 702.112
R52543 vp_n.n3429 vp_n.t593 702.112
R52544 vp_n.n3426 vp_n.t189 702.112
R52545 vp_n.n1783 vp_n.t360 702.112
R52546 vp_n.n232 vp_n.t591 702.112
R52547 vp_n.n3439 vp_n.t193 702.112
R52548 vp_n.n3436 vp_n.t394 702.112
R52549 vp_n.n1793 vp_n.t241 702.112
R52550 vp_n.n242 vp_n.t500 702.112
R52551 vp_n.n3449 vp_n.t112 702.112
R52552 vp_n.n3446 vp_n.t307 702.112
R52553 vp_n.n1803 vp_n.t370 702.112
R52554 vp_n.n252 vp_n.t596 702.112
R52555 vp_n.n3459 vp_n.t195 702.112
R52556 vp_n.n3456 vp_n.t397 702.112
R52557 vp_n.n1813 vp_n.t261 702.112
R52558 vp_n.n262 vp_n.t520 702.112
R52559 vp_n.n3469 vp_n.t128 702.112
R52560 vp_n.n3466 vp_n.t326 702.112
R52561 vp_n.n1823 vp_n.t255 702.112
R52562 vp_n.n272 vp_n.t514 702.112
R52563 vp_n.n3479 vp_n.t121 702.112
R52564 vp_n.n3476 vp_n.t318 702.112
R52565 vp_n.n1833 vp_n.t583 702.112
R52566 vp_n.n282 vp_n.t197 702.112
R52567 vp_n.n3489 vp_n.t399 702.112
R52568 vp_n.n3486 vp_n.t599 702.112
R52569 vp_n.n1843 vp_n.t488 702.112
R52570 vp_n.n292 vp_n.t137 702.112
R52571 vp_n.n3499 vp_n.t352 702.112
R52572 vp_n.n3496 vp_n.t547 702.112
R52573 vp_n.n1853 vp_n.t480 702.112
R52574 vp_n.n302 vp_n.t133 702.112
R52575 vp_n.n3509 vp_n.t347 702.112
R52576 vp_n.n3506 vp_n.t541 702.112
R52577 vp_n.n1863 vp_n.t506 702.112
R52578 vp_n.n312 vp_n.t154 702.112
R52579 vp_n.n3519 vp_n.t363 702.112
R52580 vp_n.n3516 vp_n.t560 702.112
R52581 vp_n.n1873 vp_n.t502 702.112
R52582 vp_n.n322 vp_n.t149 702.112
R52583 vp_n.n3529 vp_n.t359 702.112
R52584 vp_n.n3526 vp_n.t556 702.112
R52585 vp_n.n1883 vp_n.t407 702.112
R52586 vp_n.n332 vp_n.t29 702.112
R52587 vp_n.n3539 vp_n.t240 702.112
R52588 vp_n.n3536 vp_n.t438 702.112
R52589 vp_n.n1893 vp_n.t125 702.112
R52590 vp_n.n342 vp_n.t369 702.112
R52591 vp_n.n3549 vp_n.t577 702.112
R52592 vp_n.n3546 vp_n.t170 702.112
R52593 vp_n.n1903 vp_n.t118 702.112
R52594 vp_n.n352 vp_n.t366 702.112
R52595 vp_n.n3559 vp_n.t571 702.112
R52596 vp_n.n3556 vp_n.t165 702.112
R52597 vp_n.n1913 vp_n.t11 702.112
R52598 vp_n.n362 vp_n.t249 702.112
R52599 vp_n.n3569 vp_n.t466 702.112
R52600 vp_n.n3566 vp_n.t54 702.112
R52601 vp_n.n1923 vp_n.t139 702.112
R52602 vp_n.n372 vp_n.t375 702.112
R52603 vp_n.n3579 vp_n.t582 702.112
R52604 vp_n.n3576 vp_n.t177 702.112
R52605 vp_n.n1933 vp_n.t20 702.112
R52606 vp_n.n382 vp_n.t274 702.112
R52607 vp_n.n3589 vp_n.t486 702.112
R52608 vp_n.n3586 vp_n.t80 702.112
R52609 vp_n.n1943 vp_n.t224 702.112
R52610 vp_n.n392 vp_n.t474 702.112
R52611 vp_n.n3599 vp_n.t87 702.112
R52612 vp_n.n3596 vp_n.t284 702.112
R52613 vp_n.n1953 vp_n.t334 702.112
R52614 vp_n.n402 vp_n.t569 702.112
R52615 vp_n.n3609 vp_n.t175 702.112
R52616 vp_n.n3606 vp_n.t373 702.112
R52617 vp_n.n1963 vp_n.t534 702.112
R52618 vp_n.n412 vp_n.t171 702.112
R52619 vp_n.n3619 vp_n.t381 702.112
R52620 vp_n.n3616 vp_n.t576 702.112
R52621 vp_n.n1973 vp_n.t528 702.112
R52622 vp_n.n422 vp_n.t166 702.112
R52623 vp_n.n3629 vp_n.t374 702.112
R52624 vp_n.n3626 vp_n.t570 702.112
R52625 vp_n.n1983 vp_n.t550 702.112
R52626 vp_n.n432 vp_n.t182 702.112
R52627 vp_n.n3639 vp_n.t390 702.112
R52628 vp_n.n3636 vp_n.t587 702.112
R52629 vp_n.n1993 vp_n.t151 702.112
R52630 vp_n.n442 vp_n.t385 702.112
R52631 vp_n.n3649 vp_n.t592 702.112
R52632 vp_n.n3646 vp_n.t187 702.112
R52633 vp_n.n2003 vp_n.t425 702.112
R52634 vp_n.n452 vp_n.t79 702.112
R52635 vp_n.n3659 vp_n.t294 702.112
R52636 vp_n.n3656 vp_n.t487 702.112
R52637 vp_n.n2013 vp_n.t161 702.112
R52638 vp_n.n462 vp_n.t395 702.112
R52639 vp_n.n3669 vp_n.t597 702.112
R52640 vp_n.n3666 vp_n.t194 702.112
R52641 vp_n.n2023 vp_n.t443 702.112
R52642 vp_n.n472 vp_n.t99 702.112
R52643 vp_n.n3679 vp_n.t311 702.112
R52644 vp_n.n3676 vp_n.t505 702.112
R52645 vp_n.n2033 vp_n.t40 702.112
R52646 vp_n.n482 vp_n.t304 702.112
R52647 vp_n.n3689 vp_n.t517 702.112
R52648 vp_n.n3686 vp_n.t108 702.112
R52649 vp_n.n2043 vp_n.t69 702.112
R52650 vp_n.n492 vp_n.t329 702.112
R52651 vp_n.n3699 vp_n.t540 702.112
R52652 vp_n.n3696 vp_n.t132 702.112
R52653 vp_n.n2053 vp_n.t62 702.112
R52654 vp_n.n502 vp_n.t322 702.112
R52655 vp_n.n3709 vp_n.t533 702.112
R52656 vp_n.n3706 vp_n.t124 702.112
R52657 vp_n.n2063 vp_n.t269 702.112
R52658 vp_n.n512 vp_n.t523 702.112
R52659 vp_n.n3719 vp_n.t134 702.112
R52660 vp_n.n3716 vp_n.t331 702.112
R52661 vp_n.n2073 vp_n.t88 702.112
R52662 vp_n.n522 vp_n.t341 702.112
R52663 vp_n.n3729 vp_n.t549 702.112
R52664 vp_n.n3726 vp_n.t144 702.112
R52665 vp_n.n2083 vp_n.t291 702.112
R52666 vp_n.n532 vp_n.t543 702.112
R52667 vp_n.n3739 vp_n.t150 702.112
R52668 vp_n.n3736 vp_n.t349 702.112
R52669 vp_n.n2093 vp_n.t204 702.112
R52670 vp_n.n542 vp_n.t423 702.112
R52671 vp_n.n3749 vp_n.t31 702.112
R52672 vp_n.n3746 vp_n.t227 702.112
R52673 vp_n.n2103 vp_n.t309 702.112
R52674 vp_n.n552 vp_n.t557 702.112
R52675 vp_n.n3759 vp_n.t160 702.112
R52676 vp_n.n3756 vp_n.t361 702.112
R52677 vp_n.n2113 vp_n.t207 702.112
R52678 vp_n.n562 vp_n.t440 702.112
R52679 vp_n.n3769 vp_n.t45 702.112
R52680 vp_n.n3766 vp_n.t245 702.112
R52681 vp_n.n2123 vp_n.t206 702.112
R52682 vp_n.n572 vp_n.t433 702.112
R52683 vp_n.n3779 vp_n.t39 702.112
R52684 vp_n.n3776 vp_n.t237 702.112
R52685 vp_n.n2133 vp_n.t531 702.112
R52686 vp_n.n582 vp_n.t167 702.112
R52687 vp_n.n3789 vp_n.t376 702.112
R52688 vp_n.n3786 vp_n.t573 702.112
R52689 vp_n.n2143 vp_n.t417 702.112
R52690 vp_n.n592 vp_n.t56 702.112
R52691 vp_n.n3799 vp_n.t276 702.112
R52692 vp_n.n3796 vp_n.t469 702.112
R52693 vp_n.n2153 vp_n.t416 702.112
R52694 vp_n.n602 vp_n.t50 702.112
R52695 vp_n.n3809 vp_n.t266 702.112
R52696 vp_n.n3806 vp_n.t462 702.112
R52697 vp_n.n2163 vp_n.t428 702.112
R52698 vp_n.n612 vp_n.t84 702.112
R52699 vp_n.n3819 vp_n.t298 702.112
R52700 vp_n.n3816 vp_n.t491 702.112
R52701 vp_n.n2173 vp_n.t424 702.112
R52702 vp_n.n622 vp_n.t72 702.112
R52703 vp_n.n3829 vp_n.t290 702.112
R52704 vp_n.n3826 vp_n.t483 702.112
R52705 vp_n.n2183 vp_n.t9 702.112
R52706 vp_n.n632 vp_n.t244 702.112
R52707 vp_n.n3839 vp_n.t458 702.112
R52708 vp_n.n3836 vp_n.t46 702.112
R52709 vp_n.n2193 vp_n.t344 702.112
R52710 vp_n.n642 vp_n.t578 702.112
R52711 vp_n.n3849 vp_n.t184 702.112
R52712 vp_n.n3846 vp_n.t382 702.112
R52713 vp_n.n2203 vp_n.t338 702.112
R52714 vp_n.n652 vp_n.t572 702.112
R52715 vp_n.n3859 vp_n.t178 702.112
R52716 vp_n.n3856 vp_n.t377 702.112
R52717 vp_n.n2213 vp_n.t221 702.112
R52718 vp_n.n662 vp_n.t470 702.112
R52719 vp_n.n3869 vp_n.t83 702.112
R52720 vp_n.n3866 vp_n.t278 702.112
R52721 vp_n.n2223 vp_n.t353 702.112
R52722 vp_n.n672 vp_n.t584 702.112
R52723 vp_n.n3879 vp_n.t188 702.112
R52724 vp_n.n3876 vp_n.t387 702.112
R52725 vp_n.n2233 vp_n.t231 702.112
R52726 vp_n.n682 vp_n.t492 702.112
R52727 vp_n.n3889 vp_n.t102 702.112
R52728 vp_n.n3886 vp_n.t297 702.112
R52729 vp_n.n2243 vp_n.t437 702.112
R52730 vp_n.n692 vp_n.t91 702.112
R52731 vp_n.n3899 vp_n.t306 702.112
R52732 vp_n.n3896 vp_n.t499 702.112
R52733 vp_n.n2253 vp_n.t251 702.112
R52734 vp_n.n702 vp_n.t510 702.112
R52735 vp_n.n3909 vp_n.t117 702.112
R52736 vp_n.n3906 vp_n.t314 702.112
R52737 vp_n.n2263 vp_n.t454 702.112
R52738 vp_n.n712 vp_n.t111 702.112
R52739 vp_n.n3919 vp_n.t325 702.112
R52740 vp_n.n3916 vp_n.t519 702.112
R52741 vp_n.n2273 vp_n.t277 702.112
R52742 vp_n.n722 vp_n.t527 702.112
R52743 vp_n.n3929 vp_n.t138 702.112
R52744 vp_n.n3926 vp_n.t336 702.112
R52745 vp_n.n2283 vp_n.t476 702.112
R52746 vp_n.n732 vp_n.t127 702.112
R52747 vp_n.n3939 vp_n.t343 702.112
R52748 vp_n.n3936 vp_n.t536 702.112
R52749 vp_n.n2293 vp_n.t77 702.112
R52750 vp_n.n742 vp_n.t333 702.112
R52751 vp_n.n3949 vp_n.t545 702.112
R52752 vp_n.n3946 vp_n.t136 702.112
R52753 vp_n.n2303 vp_n.t498 702.112
R52754 vp_n.n752 vp_n.t146 702.112
R52755 vp_n.n3959 vp_n.t356 702.112
R52756 vp_n.n3956 vp_n.t553 702.112
R52757 vp_n.n2313 vp_n.t98 702.112
R52758 vp_n.n762 vp_n.t351 702.112
R52759 vp_n.n3969 vp_n.t559 702.112
R52760 vp_n.n3966 vp_n.t153 702.112
R52761 vp_n.n2323 vp_n.t404 702.112
R52762 vp_n.n772 vp_n.t22 702.112
R52763 vp_n.n3979 vp_n.t230 702.112
R52764 vp_n.n3976 vp_n.t427 702.112
R52765 vp_n.n2333 vp_n.t115 702.112
R52766 vp_n.n782 vp_n.t362 702.112
R52767 vp_n.n3989 vp_n.t568 702.112
R52768 vp_n.n3986 vp_n.t163 702.112
R52769 vp_n.n2343 vp_n.t10 702.112
R52770 vp_n.n792 vp_n.t247 702.112
R52771 vp_n.n3999 vp_n.t461 702.112
R52772 vp_n.n3996 vp_n.t49 702.112
R52773 vp_n.n2353 vp_n.t7 702.112
R52774 vp_n.n802 vp_n.t239 702.112
R52775 vp_n.n4009 vp_n.t453 702.112
R52776 vp_n.n4006 vp_n.t42 702.112
R52777 vp_n.n2363 vp_n.t339 702.112
R52778 vp_n.n812 vp_n.t575 702.112
R52779 vp_n.n4019 vp_n.t181 702.112
R52780 vp_n.n4016 vp_n.t379 702.112
R52781 vp_n.n2373 vp_n.t16 702.112
R52782 vp_n.n822 vp_n.t260 702.112
R52783 vp_n.n4029 vp_n.t475 702.112
R52784 vp_n.n4026 vp_n.t65 702.112
R52785 vp_n.n2383 vp_n.t219 702.112
R52786 vp_n.n832 vp_n.t464 702.112
R52787 vp_n.n4039 vp_n.t76 702.112
R52788 vp_n.n4036 vp_n.t272 702.112
R52789 vp_n.n2393 vp_n.t234 702.112
R52790 vp_n.n842 vp_n.t496 702.112
R52791 vp_n.n4049 vp_n.t105 702.112
R52792 vp_n.n4046 vp_n.t302 702.112
R52793 vp_n.n2403 vp_n.t229 702.112
R52794 vp_n.n852 vp_n.t485 702.112
R52795 vp_n.n4059 vp_n.t96 702.112
R52796 vp_n.n4056 vp_n.t293 702.112
R52797 vp_n.n2413 vp_n.t415 702.112
R52798 vp_n.n862 vp_n.t51 702.112
R52799 vp_n.n4069 vp_n.t268 702.112
R52800 vp_n.n4066 vp_n.t460 702.112
R52801 vp_n.n2423 vp_n.t546 702.112
R52802 vp_n.n872 vp_n.t174 702.112
R52803 vp_n.n4079 vp_n.t386 702.112
R52804 vp_n.n4076 vp_n.t581 702.112
R52805 vp_n.n2433 vp_n.t142 702.112
R52806 vp_n.n882 vp_n.t380 702.112
R52807 vp_n.n4089 vp_n.t586 702.112
R52808 vp_n.n4086 vp_n.t180 702.112
R52809 vp_n.n2443 vp_n.t24 702.112
R52810 vp_n.n892 vp_n.t280 702.112
R52811 vp_n.n4099 vp_n.t495 702.112
R52812 vp_n.n4096 vp_n.t86 702.112
R52813 vp_n.n2453 vp_n.t158 702.112
R52814 vp_n.n902 vp_n.t389 702.112
R52815 vp_n.n4109 vp_n.t594 702.112
R52816 vp_n.n4106 vp_n.t190 702.112
R52817 vp_n.n2463 vp_n.t36 702.112
R52818 vp_n.n912 vp_n.t301 702.112
R52819 vp_n.n4119 vp_n.t513 702.112
R52820 vp_n.n4116 vp_n.t106 702.112
R52821 vp_n.n2473 vp_n.t33 702.112
R52822 vp_n.n922 vp_n.t292 702.112
R52823 vp_n.n4129 vp_n.t504 702.112
R52824 vp_n.n4126 vp_n.t97 702.112
R52825 vp_n.n2483 vp_n.t57 702.112
R52826 vp_n.n932 vp_n.t317 702.112
R52827 vp_n.n4139 vp_n.t530 702.112
R52828 vp_n.n4136 vp_n.t120 702.112
R52829 vp_n.n2493 vp_n.t263 702.112
R52830 vp_n.n942 vp_n.t521 702.112
R52831 vp_n.n4149 vp_n.t131 702.112
R52832 vp_n.n4146 vp_n.t328 702.112
R52833 vp_n.n2503 vp_n.t257 702.112
R52834 vp_n.n952 vp_n.t515 702.112
R52835 vp_n.n4159 vp_n.t123 702.112
R52836 vp_n.n4156 vp_n.t320 702.112
R52837 vp_n.n2513 vp_n.t286 702.112
R52838 vp_n.n962 vp_n.t539 702.112
R52839 vp_n.n4169 vp_n.t148 702.112
R52840 vp_n.n4166 vp_n.t346 702.112
R52841 vp_n.n2523 vp_n.t282 702.112
R52842 vp_n.n972 vp_n.t532 702.112
R52843 vp_n.n4179 vp_n.t143 702.112
R52844 vp_n.n4176 vp_n.t340 702.112
R52845 vp_n.n2533 vp_n.t202 702.112
R52846 vp_n.n982 vp_n.t418 702.112
R52847 vp_n.n4189 vp_n.t25 702.112
R52848 vp_n.n4186 vp_n.t222 702.112
R52849 vp_n.n2543 vp_n.t507 702.112
R52850 vp_n.n992 vp_n.t155 702.112
R52851 vp_n.n4199 vp_n.t365 702.112
R52852 vp_n.n4196 vp_n.t562 702.112
R52853 vp_n.n2553 vp_n.t205 702.112
R52854 vp_n.n1002 vp_n.t431 702.112
R52855 vp_n.n4209 vp_n.t37 702.112
R52856 vp_n.n4206 vp_n.t235 702.112
R52857 vp_n.n2563 vp_n.t408 702.112
R52858 vp_n.n1012 vp_n.t30 702.112
R52859 vp_n.n4219 vp_n.t243 702.112
R52860 vp_n.n4216 vp_n.t439 702.112
R52861 vp_n.n2573 vp_n.t212 702.112
R52862 vp_n.n1022 vp_n.t447 702.112
R52863 vp_n.n4229 vp_n.t58 702.112
R52864 vp_n.n4226 vp_n.t254 702.112
R52865 vp_n.n2583 vp_n.t413 702.112
R52866 vp_n.n1032 vp_n.t44 702.112
R52867 vp_n.n4239 vp_n.t262 702.112
R52868 vp_n.n4236 vp_n.t456 702.112
R52869 vp_n.n2593 vp_n.t12 702.112
R52870 vp_n.n1042 vp_n.t250 702.112
R52871 vp_n.n4249 vp_n.t467 702.112
R52872 vp_n.n4246 vp_n.t55 702.112
R52873 vp_n.n2603 vp_n.t422 702.112
R52874 vp_n.n1052 vp_n.t67 702.112
R52875 vp_n.n4259 vp_n.t285 702.112
R52876 vp_n.n4256 vp_n.t478 702.112
R52877 vp_n.n2613 vp_n.t21 702.112
R52878 vp_n.n1062 vp_n.t275 702.112
R52879 vp_n.n4269 vp_n.t489 702.112
R52880 vp_n.n4266 vp_n.t81 702.112
R52881 vp_n.n2623 vp_n.t400 702.112
R52882 vp_n.n1072 vp_n.t0 702.112
R52883 vp_n.n4279 vp_n.t201 702.112
R52884 vp_n.n4276 vp_n.t402 702.112
R52885 vp_n.n2633 vp_n.t34 702.112
R52886 vp_n.n1082 vp_n.t296 702.112
R52887 vp_n.n4289 vp_n.t508 702.112
R52888 vp_n.n4286 vp_n.t100 702.112
R52889 vp_n.n2643 vp_n.t220 702.112
R52890 vp_n.n1092 vp_n.t465 702.112
R52891 vp_n.n4299 vp_n.t78 702.112
R52892 vp_n.n4296 vp_n.t273 702.112
R52893 vp_n.n2653 vp_n.t215 702.112
R52894 vp_n.n1102 vp_n.t457 702.112
R52895 vp_n.n4309 vp_n.t68 702.112
R52896 vp_n.n4306 vp_n.t264 702.112
R52897 vp_n.n2663 vp_n.t552 702.112
R52898 vp_n.n1112 vp_n.t183 702.112
R52899 vp_n.n4319 vp_n.t391 702.112
R52900 vp_n.n4316 vp_n.t588 702.112
R52901 vp_n.n2673 vp_n.t226 702.112
R52902 vp_n.n1122 vp_n.t479 702.112
R52903 vp_n.n4329 vp_n.t92 702.112
R52904 vp_n.n4326 vp_n.t287 702.112
R52905 vp_n.n2683 vp_n.t426 702.112
R52906 vp_n.n1132 vp_n.t82 702.112
R52907 vp_n.n4339 vp_n.t295 702.112
R52908 vp_n.n4336 vp_n.t490 702.112
R52909 vp_n.n2693 vp_n.t449 702.112
R52910 vp_n.n1142 vp_n.t107 702.112
R52911 vp_n.n4349 vp_n.t321 702.112
R52912 vp_n.n4346 vp_n.t516 702.112
R52913 vp_n.n2703 vp_n.t444 702.112
R52914 vp_n.n1152 vp_n.t101 702.112
R52915 vp_n.n4359 vp_n.t313 702.112
R52916 vp_n.n4356 vp_n.t509 702.112
R52917 vp_n.n2713 vp_n.t401 702.112
R52918 vp_n.n1162 vp_n.t5 702.112
R52919 vp_n.n4369 vp_n.t210 702.112
R52920 vp_n.n4366 vp_n.t409 702.112
R52921 vp_n.n2723 vp_n.t468 702.112
R52922 vp_n.n1172 vp_n.t116 702.112
R52923 vp_n.n4379 vp_n.t335 702.112
R52924 vp_n.n4376 vp_n.t526 702.112
R52925 vp_n.n2733 vp_n.t63 702.112
R52926 vp_n.n1182 vp_n.t324 702.112
R52927 vp_n.n4389 vp_n.t535 702.112
R52928 vp_n.n4386 vp_n.t126 702.112
R52929 vp_n.n2743 vp_n.t1 702.112
R52930 vp_n.n1192 vp_n.t213 702.112
R52931 vp_n.n4399 vp_n.t420 702.112
R52932 vp_n.n4396 vp_n.t14 702.112
R52933 vp_n.n2753 vp_n.t90 702.112
R52934 vp_n.n1202 vp_n.t342 702.112
R52935 vp_n.n4409 vp_n.t551 702.112
R52936 vp_n.n4406 vp_n.t145 702.112
R52937 vp_n.n2763 vp_n.t2 702.112
R52938 vp_n.n1212 vp_n.t223 702.112
R52939 vp_n.n4419 vp_n.t432 702.112
R52940 vp_n.n4416 vp_n.t26 702.112
R52941 vp_n.n2773 vp_n.t110 702.112
R52942 vp_n.n1222 vp_n.t355 702.112
R52943 vp_n.n4429 vp_n.t564 702.112
R52944 vp_n.n4426 vp_n.t159 702.112
R52945 vp_n.n2783 vp_n.t6 702.112
R52946 vp_n.n1232 vp_n.t236 702.112
R52947 vp_n.n4439 vp_n.t448 702.112
R52948 vp_n.n4436 vp_n.t38 702.112
R52949 vp_n.n2793 vp_n.t208 702.112
R52950 vp_n.n1242 vp_n.t441 702.112
R52951 vp_n.n4449 vp_n.t47 702.112
R52952 vp_n.n4446 vp_n.t246 702.112
R52953 vp_n.n2803 vp_n.t15 702.112
R52954 vp_n.n1252 vp_n.t256 702.112
R52955 vp_n.n4459 vp_n.t472 702.112
R52956 vp_n.n4456 vp_n.t60 702.112
R52957 vp_n.n2813 vp_n.t216 702.112
R52958 vp_n.n1262 vp_n.t459 702.112
R52959 vp_n.n4469 vp_n.t70 702.112
R52960 vp_n.n4466 vp_n.t265 702.112
R52961 vp_n.n2823 vp_n.t214 702.112
R52962 vp_n.n1272 vp_n.t452 702.112
R52963 vp_n.n4479 vp_n.t64 702.112
R52964 vp_n.n4476 vp_n.t258 702.112
R52965 vp_n.n2833 vp_n.t228 702.112
R52966 vp_n.n1282 vp_n.t481 702.112
R52967 vp_n.n4489 vp_n.t93 702.112
R52968 vp_n.n4486 vp_n.t288 702.112
R52969 vp_n.n2843 vp_n.t429 702.112
R52970 vp_n.n1292 vp_n.t85 702.112
R52971 vp_n.n4499 vp_n.t299 702.112
R52972 vp_n.n4496 vp_n.t493 702.112
R52973 vp_n.n2853 vp_n.t198 702.112
R52974 vp_n.n1302 vp_n.t403 702.112
R52975 vp_n.n4509 vp_n.t3 702.112
R52976 vp_n.n4506 vp_n.t203 702.112
R52977 vp_n.n2863 vp_n.t445 702.112
R52978 vp_n.n1312 vp_n.t103 702.112
R52979 vp_n.n4519 vp_n.t315 702.112
R52980 vp_n.n4516 vp_n.t511 702.112
R52981 vp_n.n2873 vp_n.t421 702.112
R52982 vp_n.n1322 vp_n.t61 702.112
R52983 vp_n.n4529 vp_n.t283 702.112
R52984 vp_n.n4526 vp_n.t473 702.112
R52985 vp_n.n2883 vp_n.t18 702.112
R52986 vp_n.n1332 vp_n.t267 702.112
R52987 vp_n.n4539 vp_n.t482 702.112
R52988 vp_n.n4536 vp_n.t71 702.112
R52989 vp_n.n2893 vp_n.t357 702.112
R52990 vp_n.n1342 vp_n.t590 702.112
R52991 vp_n.n4549 vp_n.t192 702.112
R52992 vp_n.n4546 vp_n.t393 702.112
R52993 vp_n.n2903 vp_n.t32 702.112
R52994 vp_n.n1352 vp_n.t289 702.112
R52995 vp_n.n4559 vp_n.t503 702.112
R52996 vp_n.n4556 vp_n.t94 702.112
R52997 vp_n.n2913 vp_n.t232 702.112
R52998 vp_n.n1362 vp_n.t494 702.112
R52999 vp_n.n4569 vp_n.t104 702.112
R53000 vp_n.n4566 vp_n.t300 702.112
R53001 vp_n.n2923 vp_n.t48 702.112
R53002 vp_n.n1372 vp_n.t308 702.112
R53003 vp_n.n4579 vp_n.t522 702.112
R53004 vp_n.n4576 vp_n.t113 702.112
R53005 vp_n.n2933 vp_n.t252 702.112
R53006 vp_n.n1382 vp_n.t512 702.112
R53007 vp_n.n4589 vp_n.t119 702.112
R53008 vp_n.n4586 vp_n.t316 702.112
R53009 vp_n.n2943 vp_n.t199 702.112
R53010 vp_n.n1392 vp_n.t410 702.112
R53011 vp_n.n4599 vp_n.t13 702.112
R53012 vp_n.n4596 vp_n.t211 702.112
R53013 vp_n.n2953 vp_n.t279 702.112
R53014 vp_n.n1402 vp_n.t529 702.112
R53015 vp_n.n4609 vp_n.t140 702.112
R53016 vp_n.n4606 vp_n.t337 702.112
R53017 vp_n.n2963 vp_n.t477 702.112
R53018 vp_n.n1412 vp_n.t130 702.112
R53019 vp_n.n4619 vp_n.t345 702.112
R53020 vp_n.n4616 vp_n.t538 702.112
R53021 vp_n.n2973 vp_n.t200 702.112
R53022 vp_n.n1422 vp_n.t414 702.112
R53023 vp_n.n4629 vp_n.t17 702.112
R53024 vp_n.n4626 vp_n.t217 702.112
R53025 vp_n.n2983 vp_n.t501 702.112
R53026 vp_n.n1432 vp_n.t147 702.112
R53027 vp_n.n4639 vp_n.t358 702.112
R53028 vp_n.n4636 vp_n.t555 702.112
R53029 vp_n.n2993 vp_n.t406 702.112
R53030 vp_n.n1442 vp_n.t28 702.112
R53031 vp_n.n4649 vp_n.t238 702.112
R53032 vp_n.n4646 vp_n.t436 702.112
R53033 vp_n.n3003 vp_n.t405 702.112
R53034 vp_n.n1452 vp_n.t23 702.112
R53035 vp_n.n4659 vp_n.t233 702.112
R53036 vp_n.n4656 vp_n.t430 702.112
R53037 vp_n.n3013 vp_n.t412 702.112
R53038 vp_n.n1462 vp_n.t41 702.112
R53039 vp_n.n4669 vp_n.t259 702.112
R53040 vp_n.n4666 vp_n.t451 702.112
R53041 vp_n.n3023 vp_n.t411 702.112
R53042 vp_n.n1472 vp_n.t35 702.112
R53043 vp_n.n4679 vp_n.t253 702.112
R53044 vp_n.n4676 vp_n.t446 702.112
R53045 vp_n.n3033 vp_n.t8 702.112
R53046 vp_n.n1482 vp_n.t242 702.112
R53047 vp_n.n4689 vp_n.t455 702.112
R53048 vp_n.n4686 vp_n.t43 702.112
R53049 vp_n.n4699 vp_n.t484 702.112
R53050 vp_n.n4696 vp_n.t75 702.112
R53051 vp_n.n1492 vp_n.t271 702.112
R53052 vp_n.n1563 vp_n.t435 702.112
R53053 vp_n.n12 vp_n.t89 702.112
R53054 vp_n.n3216 vp_n.t497 702.112
R53055 vp_n.n3219 vp_n.t305 702.112
R53056 vp_n.n3209 vp_n.t392 702.112
R53057 vp_n.n3206 vp_n.t589 702.112
R53058 vp_n.n2 vp_n.t185 702.112
R53059 vp_n.n1553 vp_n.t554 702.112
R53060 vp_n.n1574 vp_n.n1573 13.653
R53061 vp_n.n3227 vp_n.n3226 13.653
R53062 vp_n.n23 vp_n.n22 13.653
R53063 vp_n.n1587 vp_n.n1586 13.653
R53064 vp_n.n3240 vp_n.n3239 13.653
R53065 vp_n.n36 vp_n.n35 13.653
R53066 vp_n.n33 vp_n.n32 13.653
R53067 vp_n.n1594 vp_n.n1593 13.653
R53068 vp_n.n3247 vp_n.n3246 13.653
R53069 vp_n.n43 vp_n.n42 13.653
R53070 vp_n.n1607 vp_n.n1606 13.653
R53071 vp_n.n3260 vp_n.n3259 13.653
R53072 vp_n.n56 vp_n.n55 13.653
R53073 vp_n.n53 vp_n.n52 13.653
R53074 vp_n.n1614 vp_n.n1613 13.653
R53075 vp_n.n3267 vp_n.n3266 13.653
R53076 vp_n.n63 vp_n.n62 13.653
R53077 vp_n.n1627 vp_n.n1626 13.653
R53078 vp_n.n3280 vp_n.n3279 13.653
R53079 vp_n.n76 vp_n.n75 13.653
R53080 vp_n.n73 vp_n.n72 13.653
R53081 vp_n.n1634 vp_n.n1633 13.653
R53082 vp_n.n3287 vp_n.n3286 13.653
R53083 vp_n.n83 vp_n.n82 13.653
R53084 vp_n.n1647 vp_n.n1646 13.653
R53085 vp_n.n3300 vp_n.n3299 13.653
R53086 vp_n.n96 vp_n.n95 13.653
R53087 vp_n.n93 vp_n.n92 13.653
R53088 vp_n.n1654 vp_n.n1653 13.653
R53089 vp_n.n3307 vp_n.n3306 13.653
R53090 vp_n.n103 vp_n.n102 13.653
R53091 vp_n.n1667 vp_n.n1666 13.653
R53092 vp_n.n3320 vp_n.n3319 13.653
R53093 vp_n.n116 vp_n.n115 13.653
R53094 vp_n.n113 vp_n.n112 13.653
R53095 vp_n.n1674 vp_n.n1673 13.653
R53096 vp_n.n3327 vp_n.n3326 13.653
R53097 vp_n.n123 vp_n.n122 13.653
R53098 vp_n.n1687 vp_n.n1686 13.653
R53099 vp_n.n3340 vp_n.n3339 13.653
R53100 vp_n.n136 vp_n.n135 13.653
R53101 vp_n.n133 vp_n.n132 13.653
R53102 vp_n.n1694 vp_n.n1693 13.653
R53103 vp_n.n3347 vp_n.n3346 13.653
R53104 vp_n.n143 vp_n.n142 13.653
R53105 vp_n.n1707 vp_n.n1706 13.653
R53106 vp_n.n3360 vp_n.n3359 13.653
R53107 vp_n.n156 vp_n.n155 13.653
R53108 vp_n.n153 vp_n.n152 13.653
R53109 vp_n.n1714 vp_n.n1713 13.653
R53110 vp_n.n3367 vp_n.n3366 13.653
R53111 vp_n.n163 vp_n.n162 13.653
R53112 vp_n.n1727 vp_n.n1726 13.653
R53113 vp_n.n3380 vp_n.n3379 13.653
R53114 vp_n.n176 vp_n.n175 13.653
R53115 vp_n.n173 vp_n.n172 13.653
R53116 vp_n.n1734 vp_n.n1733 13.653
R53117 vp_n.n3387 vp_n.n3386 13.653
R53118 vp_n.n183 vp_n.n182 13.653
R53119 vp_n.n1747 vp_n.n1746 13.653
R53120 vp_n.n3400 vp_n.n3399 13.653
R53121 vp_n.n196 vp_n.n195 13.653
R53122 vp_n.n193 vp_n.n192 13.653
R53123 vp_n.n1754 vp_n.n1753 13.653
R53124 vp_n.n3407 vp_n.n3406 13.653
R53125 vp_n.n203 vp_n.n202 13.653
R53126 vp_n.n1767 vp_n.n1766 13.653
R53127 vp_n.n3420 vp_n.n3419 13.653
R53128 vp_n.n216 vp_n.n215 13.653
R53129 vp_n.n213 vp_n.n212 13.653
R53130 vp_n.n1774 vp_n.n1773 13.653
R53131 vp_n.n3427 vp_n.n3426 13.653
R53132 vp_n.n223 vp_n.n222 13.653
R53133 vp_n.n1787 vp_n.n1786 13.653
R53134 vp_n.n3440 vp_n.n3439 13.653
R53135 vp_n.n236 vp_n.n235 13.653
R53136 vp_n.n233 vp_n.n232 13.653
R53137 vp_n.n1794 vp_n.n1793 13.653
R53138 vp_n.n3447 vp_n.n3446 13.653
R53139 vp_n.n243 vp_n.n242 13.653
R53140 vp_n.n1807 vp_n.n1806 13.653
R53141 vp_n.n3460 vp_n.n3459 13.653
R53142 vp_n.n256 vp_n.n255 13.653
R53143 vp_n.n253 vp_n.n252 13.653
R53144 vp_n.n1814 vp_n.n1813 13.653
R53145 vp_n.n3467 vp_n.n3466 13.653
R53146 vp_n.n263 vp_n.n262 13.653
R53147 vp_n.n1827 vp_n.n1826 13.653
R53148 vp_n.n3480 vp_n.n3479 13.653
R53149 vp_n.n276 vp_n.n275 13.653
R53150 vp_n.n273 vp_n.n272 13.653
R53151 vp_n.n1834 vp_n.n1833 13.653
R53152 vp_n.n3487 vp_n.n3486 13.653
R53153 vp_n.n283 vp_n.n282 13.653
R53154 vp_n.n1847 vp_n.n1846 13.653
R53155 vp_n.n3500 vp_n.n3499 13.653
R53156 vp_n.n296 vp_n.n295 13.653
R53157 vp_n.n293 vp_n.n292 13.653
R53158 vp_n.n1854 vp_n.n1853 13.653
R53159 vp_n.n3507 vp_n.n3506 13.653
R53160 vp_n.n303 vp_n.n302 13.653
R53161 vp_n.n1867 vp_n.n1866 13.653
R53162 vp_n.n3520 vp_n.n3519 13.653
R53163 vp_n.n316 vp_n.n315 13.653
R53164 vp_n.n313 vp_n.n312 13.653
R53165 vp_n.n1874 vp_n.n1873 13.653
R53166 vp_n.n3527 vp_n.n3526 13.653
R53167 vp_n.n323 vp_n.n322 13.653
R53168 vp_n.n1887 vp_n.n1886 13.653
R53169 vp_n.n3540 vp_n.n3539 13.653
R53170 vp_n.n336 vp_n.n335 13.653
R53171 vp_n.n333 vp_n.n332 13.653
R53172 vp_n.n1894 vp_n.n1893 13.653
R53173 vp_n.n3547 vp_n.n3546 13.653
R53174 vp_n.n343 vp_n.n342 13.653
R53175 vp_n.n1907 vp_n.n1906 13.653
R53176 vp_n.n3560 vp_n.n3559 13.653
R53177 vp_n.n356 vp_n.n355 13.653
R53178 vp_n.n353 vp_n.n352 13.653
R53179 vp_n.n1914 vp_n.n1913 13.653
R53180 vp_n.n3567 vp_n.n3566 13.653
R53181 vp_n.n363 vp_n.n362 13.653
R53182 vp_n.n1927 vp_n.n1926 13.653
R53183 vp_n.n3580 vp_n.n3579 13.653
R53184 vp_n.n376 vp_n.n375 13.653
R53185 vp_n.n373 vp_n.n372 13.653
R53186 vp_n.n1934 vp_n.n1933 13.653
R53187 vp_n.n3587 vp_n.n3586 13.653
R53188 vp_n.n383 vp_n.n382 13.653
R53189 vp_n.n1947 vp_n.n1946 13.653
R53190 vp_n.n3600 vp_n.n3599 13.653
R53191 vp_n.n396 vp_n.n395 13.653
R53192 vp_n.n393 vp_n.n392 13.653
R53193 vp_n.n1954 vp_n.n1953 13.653
R53194 vp_n.n3607 vp_n.n3606 13.653
R53195 vp_n.n403 vp_n.n402 13.653
R53196 vp_n.n1967 vp_n.n1966 13.653
R53197 vp_n.n3620 vp_n.n3619 13.653
R53198 vp_n.n416 vp_n.n415 13.653
R53199 vp_n.n413 vp_n.n412 13.653
R53200 vp_n.n1974 vp_n.n1973 13.653
R53201 vp_n.n3627 vp_n.n3626 13.653
R53202 vp_n.n423 vp_n.n422 13.653
R53203 vp_n.n1987 vp_n.n1986 13.653
R53204 vp_n.n3640 vp_n.n3639 13.653
R53205 vp_n.n436 vp_n.n435 13.653
R53206 vp_n.n433 vp_n.n432 13.653
R53207 vp_n.n1994 vp_n.n1993 13.653
R53208 vp_n.n3647 vp_n.n3646 13.653
R53209 vp_n.n443 vp_n.n442 13.653
R53210 vp_n.n2007 vp_n.n2006 13.653
R53211 vp_n.n3660 vp_n.n3659 13.653
R53212 vp_n.n456 vp_n.n455 13.653
R53213 vp_n.n453 vp_n.n452 13.653
R53214 vp_n.n2014 vp_n.n2013 13.653
R53215 vp_n.n3667 vp_n.n3666 13.653
R53216 vp_n.n463 vp_n.n462 13.653
R53217 vp_n.n2027 vp_n.n2026 13.653
R53218 vp_n.n3680 vp_n.n3679 13.653
R53219 vp_n.n476 vp_n.n475 13.653
R53220 vp_n.n473 vp_n.n472 13.653
R53221 vp_n.n2034 vp_n.n2033 13.653
R53222 vp_n.n3687 vp_n.n3686 13.653
R53223 vp_n.n483 vp_n.n482 13.653
R53224 vp_n.n2047 vp_n.n2046 13.653
R53225 vp_n.n3700 vp_n.n3699 13.653
R53226 vp_n.n496 vp_n.n495 13.653
R53227 vp_n.n493 vp_n.n492 13.653
R53228 vp_n.n2054 vp_n.n2053 13.653
R53229 vp_n.n3707 vp_n.n3706 13.653
R53230 vp_n.n503 vp_n.n502 13.653
R53231 vp_n.n2067 vp_n.n2066 13.653
R53232 vp_n.n3720 vp_n.n3719 13.653
R53233 vp_n.n516 vp_n.n515 13.653
R53234 vp_n.n513 vp_n.n512 13.653
R53235 vp_n.n2074 vp_n.n2073 13.653
R53236 vp_n.n3727 vp_n.n3726 13.653
R53237 vp_n.n523 vp_n.n522 13.653
R53238 vp_n.n2087 vp_n.n2086 13.653
R53239 vp_n.n3740 vp_n.n3739 13.653
R53240 vp_n.n536 vp_n.n535 13.653
R53241 vp_n.n533 vp_n.n532 13.653
R53242 vp_n.n2094 vp_n.n2093 13.653
R53243 vp_n.n3747 vp_n.n3746 13.653
R53244 vp_n.n543 vp_n.n542 13.653
R53245 vp_n.n2107 vp_n.n2106 13.653
R53246 vp_n.n3760 vp_n.n3759 13.653
R53247 vp_n.n556 vp_n.n555 13.653
R53248 vp_n.n553 vp_n.n552 13.653
R53249 vp_n.n2114 vp_n.n2113 13.653
R53250 vp_n.n3767 vp_n.n3766 13.653
R53251 vp_n.n563 vp_n.n562 13.653
R53252 vp_n.n2127 vp_n.n2126 13.653
R53253 vp_n.n3780 vp_n.n3779 13.653
R53254 vp_n.n576 vp_n.n575 13.653
R53255 vp_n.n573 vp_n.n572 13.653
R53256 vp_n.n2134 vp_n.n2133 13.653
R53257 vp_n.n3787 vp_n.n3786 13.653
R53258 vp_n.n583 vp_n.n582 13.653
R53259 vp_n.n2147 vp_n.n2146 13.653
R53260 vp_n.n3800 vp_n.n3799 13.653
R53261 vp_n.n596 vp_n.n595 13.653
R53262 vp_n.n593 vp_n.n592 13.653
R53263 vp_n.n2154 vp_n.n2153 13.653
R53264 vp_n.n3807 vp_n.n3806 13.653
R53265 vp_n.n603 vp_n.n602 13.653
R53266 vp_n.n2167 vp_n.n2166 13.653
R53267 vp_n.n3820 vp_n.n3819 13.653
R53268 vp_n.n616 vp_n.n615 13.653
R53269 vp_n.n613 vp_n.n612 13.653
R53270 vp_n.n2174 vp_n.n2173 13.653
R53271 vp_n.n3827 vp_n.n3826 13.653
R53272 vp_n.n623 vp_n.n622 13.653
R53273 vp_n.n2187 vp_n.n2186 13.653
R53274 vp_n.n3840 vp_n.n3839 13.653
R53275 vp_n.n636 vp_n.n635 13.653
R53276 vp_n.n633 vp_n.n632 13.653
R53277 vp_n.n2194 vp_n.n2193 13.653
R53278 vp_n.n3847 vp_n.n3846 13.653
R53279 vp_n.n643 vp_n.n642 13.653
R53280 vp_n.n2207 vp_n.n2206 13.653
R53281 vp_n.n3860 vp_n.n3859 13.653
R53282 vp_n.n656 vp_n.n655 13.653
R53283 vp_n.n653 vp_n.n652 13.653
R53284 vp_n.n2214 vp_n.n2213 13.653
R53285 vp_n.n3867 vp_n.n3866 13.653
R53286 vp_n.n663 vp_n.n662 13.653
R53287 vp_n.n2227 vp_n.n2226 13.653
R53288 vp_n.n3880 vp_n.n3879 13.653
R53289 vp_n.n676 vp_n.n675 13.653
R53290 vp_n.n673 vp_n.n672 13.653
R53291 vp_n.n2234 vp_n.n2233 13.653
R53292 vp_n.n3887 vp_n.n3886 13.653
R53293 vp_n.n683 vp_n.n682 13.653
R53294 vp_n.n2247 vp_n.n2246 13.653
R53295 vp_n.n3900 vp_n.n3899 13.653
R53296 vp_n.n696 vp_n.n695 13.653
R53297 vp_n.n693 vp_n.n692 13.653
R53298 vp_n.n2254 vp_n.n2253 13.653
R53299 vp_n.n3907 vp_n.n3906 13.653
R53300 vp_n.n703 vp_n.n702 13.653
R53301 vp_n.n2267 vp_n.n2266 13.653
R53302 vp_n.n3920 vp_n.n3919 13.653
R53303 vp_n.n716 vp_n.n715 13.653
R53304 vp_n.n713 vp_n.n712 13.653
R53305 vp_n.n2274 vp_n.n2273 13.653
R53306 vp_n.n3927 vp_n.n3926 13.653
R53307 vp_n.n723 vp_n.n722 13.653
R53308 vp_n.n2287 vp_n.n2286 13.653
R53309 vp_n.n3940 vp_n.n3939 13.653
R53310 vp_n.n736 vp_n.n735 13.653
R53311 vp_n.n733 vp_n.n732 13.653
R53312 vp_n.n2294 vp_n.n2293 13.653
R53313 vp_n.n3947 vp_n.n3946 13.653
R53314 vp_n.n743 vp_n.n742 13.653
R53315 vp_n.n2307 vp_n.n2306 13.653
R53316 vp_n.n3960 vp_n.n3959 13.653
R53317 vp_n.n756 vp_n.n755 13.653
R53318 vp_n.n753 vp_n.n752 13.653
R53319 vp_n.n2314 vp_n.n2313 13.653
R53320 vp_n.n3967 vp_n.n3966 13.653
R53321 vp_n.n763 vp_n.n762 13.653
R53322 vp_n.n2327 vp_n.n2326 13.653
R53323 vp_n.n3980 vp_n.n3979 13.653
R53324 vp_n.n776 vp_n.n775 13.653
R53325 vp_n.n773 vp_n.n772 13.653
R53326 vp_n.n2334 vp_n.n2333 13.653
R53327 vp_n.n3987 vp_n.n3986 13.653
R53328 vp_n.n783 vp_n.n782 13.653
R53329 vp_n.n2347 vp_n.n2346 13.653
R53330 vp_n.n4000 vp_n.n3999 13.653
R53331 vp_n.n796 vp_n.n795 13.653
R53332 vp_n.n793 vp_n.n792 13.653
R53333 vp_n.n2354 vp_n.n2353 13.653
R53334 vp_n.n4007 vp_n.n4006 13.653
R53335 vp_n.n803 vp_n.n802 13.653
R53336 vp_n.n2367 vp_n.n2366 13.653
R53337 vp_n.n4020 vp_n.n4019 13.653
R53338 vp_n.n816 vp_n.n815 13.653
R53339 vp_n.n813 vp_n.n812 13.653
R53340 vp_n.n2374 vp_n.n2373 13.653
R53341 vp_n.n4027 vp_n.n4026 13.653
R53342 vp_n.n823 vp_n.n822 13.653
R53343 vp_n.n2387 vp_n.n2386 13.653
R53344 vp_n.n4040 vp_n.n4039 13.653
R53345 vp_n.n836 vp_n.n835 13.653
R53346 vp_n.n833 vp_n.n832 13.653
R53347 vp_n.n2394 vp_n.n2393 13.653
R53348 vp_n.n4047 vp_n.n4046 13.653
R53349 vp_n.n843 vp_n.n842 13.653
R53350 vp_n.n2407 vp_n.n2406 13.653
R53351 vp_n.n4060 vp_n.n4059 13.653
R53352 vp_n.n856 vp_n.n855 13.653
R53353 vp_n.n853 vp_n.n852 13.653
R53354 vp_n.n2414 vp_n.n2413 13.653
R53355 vp_n.n4067 vp_n.n4066 13.653
R53356 vp_n.n863 vp_n.n862 13.653
R53357 vp_n.n2427 vp_n.n2426 13.653
R53358 vp_n.n4080 vp_n.n4079 13.653
R53359 vp_n.n876 vp_n.n875 13.653
R53360 vp_n.n873 vp_n.n872 13.653
R53361 vp_n.n2434 vp_n.n2433 13.653
R53362 vp_n.n4087 vp_n.n4086 13.653
R53363 vp_n.n883 vp_n.n882 13.653
R53364 vp_n.n2447 vp_n.n2446 13.653
R53365 vp_n.n4100 vp_n.n4099 13.653
R53366 vp_n.n896 vp_n.n895 13.653
R53367 vp_n.n893 vp_n.n892 13.653
R53368 vp_n.n2454 vp_n.n2453 13.653
R53369 vp_n.n4107 vp_n.n4106 13.653
R53370 vp_n.n903 vp_n.n902 13.653
R53371 vp_n.n2467 vp_n.n2466 13.653
R53372 vp_n.n4120 vp_n.n4119 13.653
R53373 vp_n.n916 vp_n.n915 13.653
R53374 vp_n.n913 vp_n.n912 13.653
R53375 vp_n.n2474 vp_n.n2473 13.653
R53376 vp_n.n4127 vp_n.n4126 13.653
R53377 vp_n.n923 vp_n.n922 13.653
R53378 vp_n.n2487 vp_n.n2486 13.653
R53379 vp_n.n4140 vp_n.n4139 13.653
R53380 vp_n.n936 vp_n.n935 13.653
R53381 vp_n.n933 vp_n.n932 13.653
R53382 vp_n.n2494 vp_n.n2493 13.653
R53383 vp_n.n4147 vp_n.n4146 13.653
R53384 vp_n.n943 vp_n.n942 13.653
R53385 vp_n.n2507 vp_n.n2506 13.653
R53386 vp_n.n4160 vp_n.n4159 13.653
R53387 vp_n.n956 vp_n.n955 13.653
R53388 vp_n.n953 vp_n.n952 13.653
R53389 vp_n.n2514 vp_n.n2513 13.653
R53390 vp_n.n4167 vp_n.n4166 13.653
R53391 vp_n.n963 vp_n.n962 13.653
R53392 vp_n.n2527 vp_n.n2526 13.653
R53393 vp_n.n4180 vp_n.n4179 13.653
R53394 vp_n.n976 vp_n.n975 13.653
R53395 vp_n.n973 vp_n.n972 13.653
R53396 vp_n.n2534 vp_n.n2533 13.653
R53397 vp_n.n4187 vp_n.n4186 13.653
R53398 vp_n.n983 vp_n.n982 13.653
R53399 vp_n.n2547 vp_n.n2546 13.653
R53400 vp_n.n4200 vp_n.n4199 13.653
R53401 vp_n.n996 vp_n.n995 13.653
R53402 vp_n.n993 vp_n.n992 13.653
R53403 vp_n.n2554 vp_n.n2553 13.653
R53404 vp_n.n4207 vp_n.n4206 13.653
R53405 vp_n.n1003 vp_n.n1002 13.653
R53406 vp_n.n2567 vp_n.n2566 13.653
R53407 vp_n.n4220 vp_n.n4219 13.653
R53408 vp_n.n1016 vp_n.n1015 13.653
R53409 vp_n.n1013 vp_n.n1012 13.653
R53410 vp_n.n2574 vp_n.n2573 13.653
R53411 vp_n.n4227 vp_n.n4226 13.653
R53412 vp_n.n1023 vp_n.n1022 13.653
R53413 vp_n.n2587 vp_n.n2586 13.653
R53414 vp_n.n4240 vp_n.n4239 13.653
R53415 vp_n.n1036 vp_n.n1035 13.653
R53416 vp_n.n1033 vp_n.n1032 13.653
R53417 vp_n.n2594 vp_n.n2593 13.653
R53418 vp_n.n4247 vp_n.n4246 13.653
R53419 vp_n.n1043 vp_n.n1042 13.653
R53420 vp_n.n2607 vp_n.n2606 13.653
R53421 vp_n.n4260 vp_n.n4259 13.653
R53422 vp_n.n1056 vp_n.n1055 13.653
R53423 vp_n.n1053 vp_n.n1052 13.653
R53424 vp_n.n2614 vp_n.n2613 13.653
R53425 vp_n.n4267 vp_n.n4266 13.653
R53426 vp_n.n1063 vp_n.n1062 13.653
R53427 vp_n.n2627 vp_n.n2626 13.653
R53428 vp_n.n4280 vp_n.n4279 13.653
R53429 vp_n.n1076 vp_n.n1075 13.653
R53430 vp_n.n1073 vp_n.n1072 13.653
R53431 vp_n.n2634 vp_n.n2633 13.653
R53432 vp_n.n4287 vp_n.n4286 13.653
R53433 vp_n.n1083 vp_n.n1082 13.653
R53434 vp_n.n2647 vp_n.n2646 13.653
R53435 vp_n.n4300 vp_n.n4299 13.653
R53436 vp_n.n1096 vp_n.n1095 13.653
R53437 vp_n.n1093 vp_n.n1092 13.653
R53438 vp_n.n2654 vp_n.n2653 13.653
R53439 vp_n.n4307 vp_n.n4306 13.653
R53440 vp_n.n1103 vp_n.n1102 13.653
R53441 vp_n.n2667 vp_n.n2666 13.653
R53442 vp_n.n4320 vp_n.n4319 13.653
R53443 vp_n.n1116 vp_n.n1115 13.653
R53444 vp_n.n1113 vp_n.n1112 13.653
R53445 vp_n.n2674 vp_n.n2673 13.653
R53446 vp_n.n4327 vp_n.n4326 13.653
R53447 vp_n.n1123 vp_n.n1122 13.653
R53448 vp_n.n2687 vp_n.n2686 13.653
R53449 vp_n.n4340 vp_n.n4339 13.653
R53450 vp_n.n1136 vp_n.n1135 13.653
R53451 vp_n.n1133 vp_n.n1132 13.653
R53452 vp_n.n2694 vp_n.n2693 13.653
R53453 vp_n.n4347 vp_n.n4346 13.653
R53454 vp_n.n1143 vp_n.n1142 13.653
R53455 vp_n.n2707 vp_n.n2706 13.653
R53456 vp_n.n4360 vp_n.n4359 13.653
R53457 vp_n.n1156 vp_n.n1155 13.653
R53458 vp_n.n1153 vp_n.n1152 13.653
R53459 vp_n.n2714 vp_n.n2713 13.653
R53460 vp_n.n4367 vp_n.n4366 13.653
R53461 vp_n.n1163 vp_n.n1162 13.653
R53462 vp_n.n2727 vp_n.n2726 13.653
R53463 vp_n.n4380 vp_n.n4379 13.653
R53464 vp_n.n1176 vp_n.n1175 13.653
R53465 vp_n.n1173 vp_n.n1172 13.653
R53466 vp_n.n2734 vp_n.n2733 13.653
R53467 vp_n.n4387 vp_n.n4386 13.653
R53468 vp_n.n1183 vp_n.n1182 13.653
R53469 vp_n.n2747 vp_n.n2746 13.653
R53470 vp_n.n4400 vp_n.n4399 13.653
R53471 vp_n.n1196 vp_n.n1195 13.653
R53472 vp_n.n1193 vp_n.n1192 13.653
R53473 vp_n.n2754 vp_n.n2753 13.653
R53474 vp_n.n4407 vp_n.n4406 13.653
R53475 vp_n.n1203 vp_n.n1202 13.653
R53476 vp_n.n2767 vp_n.n2766 13.653
R53477 vp_n.n4420 vp_n.n4419 13.653
R53478 vp_n.n1216 vp_n.n1215 13.653
R53479 vp_n.n1213 vp_n.n1212 13.653
R53480 vp_n.n2774 vp_n.n2773 13.653
R53481 vp_n.n4427 vp_n.n4426 13.653
R53482 vp_n.n1223 vp_n.n1222 13.653
R53483 vp_n.n2787 vp_n.n2786 13.653
R53484 vp_n.n4440 vp_n.n4439 13.653
R53485 vp_n.n1236 vp_n.n1235 13.653
R53486 vp_n.n1233 vp_n.n1232 13.653
R53487 vp_n.n2794 vp_n.n2793 13.653
R53488 vp_n.n4447 vp_n.n4446 13.653
R53489 vp_n.n1243 vp_n.n1242 13.653
R53490 vp_n.n2807 vp_n.n2806 13.653
R53491 vp_n.n4460 vp_n.n4459 13.653
R53492 vp_n.n1256 vp_n.n1255 13.653
R53493 vp_n.n1253 vp_n.n1252 13.653
R53494 vp_n.n2814 vp_n.n2813 13.653
R53495 vp_n.n4467 vp_n.n4466 13.653
R53496 vp_n.n1263 vp_n.n1262 13.653
R53497 vp_n.n2827 vp_n.n2826 13.653
R53498 vp_n.n4480 vp_n.n4479 13.653
R53499 vp_n.n1276 vp_n.n1275 13.653
R53500 vp_n.n1273 vp_n.n1272 13.653
R53501 vp_n.n2834 vp_n.n2833 13.653
R53502 vp_n.n4487 vp_n.n4486 13.653
R53503 vp_n.n1283 vp_n.n1282 13.653
R53504 vp_n.n2847 vp_n.n2846 13.653
R53505 vp_n.n4500 vp_n.n4499 13.653
R53506 vp_n.n1296 vp_n.n1295 13.653
R53507 vp_n.n1293 vp_n.n1292 13.653
R53508 vp_n.n2854 vp_n.n2853 13.653
R53509 vp_n.n4507 vp_n.n4506 13.653
R53510 vp_n.n1303 vp_n.n1302 13.653
R53511 vp_n.n2867 vp_n.n2866 13.653
R53512 vp_n.n4520 vp_n.n4519 13.653
R53513 vp_n.n1316 vp_n.n1315 13.653
R53514 vp_n.n1313 vp_n.n1312 13.653
R53515 vp_n.n2874 vp_n.n2873 13.653
R53516 vp_n.n4527 vp_n.n4526 13.653
R53517 vp_n.n1323 vp_n.n1322 13.653
R53518 vp_n.n2887 vp_n.n2886 13.653
R53519 vp_n.n4540 vp_n.n4539 13.653
R53520 vp_n.n1336 vp_n.n1335 13.653
R53521 vp_n.n1333 vp_n.n1332 13.653
R53522 vp_n.n2894 vp_n.n2893 13.653
R53523 vp_n.n4547 vp_n.n4546 13.653
R53524 vp_n.n1343 vp_n.n1342 13.653
R53525 vp_n.n2907 vp_n.n2906 13.653
R53526 vp_n.n4560 vp_n.n4559 13.653
R53527 vp_n.n1356 vp_n.n1355 13.653
R53528 vp_n.n1353 vp_n.n1352 13.653
R53529 vp_n.n2914 vp_n.n2913 13.653
R53530 vp_n.n4567 vp_n.n4566 13.653
R53531 vp_n.n1363 vp_n.n1362 13.653
R53532 vp_n.n2927 vp_n.n2926 13.653
R53533 vp_n.n4580 vp_n.n4579 13.653
R53534 vp_n.n1376 vp_n.n1375 13.653
R53535 vp_n.n1373 vp_n.n1372 13.653
R53536 vp_n.n2934 vp_n.n2933 13.653
R53537 vp_n.n4587 vp_n.n4586 13.653
R53538 vp_n.n1383 vp_n.n1382 13.653
R53539 vp_n.n2947 vp_n.n2946 13.653
R53540 vp_n.n4600 vp_n.n4599 13.653
R53541 vp_n.n1396 vp_n.n1395 13.653
R53542 vp_n.n1393 vp_n.n1392 13.653
R53543 vp_n.n2954 vp_n.n2953 13.653
R53544 vp_n.n4607 vp_n.n4606 13.653
R53545 vp_n.n1403 vp_n.n1402 13.653
R53546 vp_n.n2967 vp_n.n2966 13.653
R53547 vp_n.n4620 vp_n.n4619 13.653
R53548 vp_n.n1416 vp_n.n1415 13.653
R53549 vp_n.n1413 vp_n.n1412 13.653
R53550 vp_n.n2974 vp_n.n2973 13.653
R53551 vp_n.n4627 vp_n.n4626 13.653
R53552 vp_n.n1423 vp_n.n1422 13.653
R53553 vp_n.n2987 vp_n.n2986 13.653
R53554 vp_n.n4640 vp_n.n4639 13.653
R53555 vp_n.n1436 vp_n.n1435 13.653
R53556 vp_n.n1433 vp_n.n1432 13.653
R53557 vp_n.n2994 vp_n.n2993 13.653
R53558 vp_n.n4647 vp_n.n4646 13.653
R53559 vp_n.n1443 vp_n.n1442 13.653
R53560 vp_n.n3007 vp_n.n3006 13.653
R53561 vp_n.n4660 vp_n.n4659 13.653
R53562 vp_n.n1456 vp_n.n1455 13.653
R53563 vp_n.n1453 vp_n.n1452 13.653
R53564 vp_n.n3014 vp_n.n3013 13.653
R53565 vp_n.n4667 vp_n.n4666 13.653
R53566 vp_n.n1463 vp_n.n1462 13.653
R53567 vp_n.n3027 vp_n.n3026 13.653
R53568 vp_n.n4680 vp_n.n4679 13.653
R53569 vp_n.n1476 vp_n.n1475 13.653
R53570 vp_n.n1473 vp_n.n1472 13.653
R53571 vp_n.n3034 vp_n.n3033 13.653
R53572 vp_n.n4687 vp_n.n4686 13.653
R53573 vp_n.n1483 vp_n.n1482 13.653
R53574 vp_n.n26 vp_n.n25 13.653
R53575 vp_n.n46 vp_n.n45 13.653
R53576 vp_n.n66 vp_n.n65 13.653
R53577 vp_n.n86 vp_n.n85 13.653
R53578 vp_n.n106 vp_n.n105 13.653
R53579 vp_n.n126 vp_n.n125 13.653
R53580 vp_n.n146 vp_n.n145 13.653
R53581 vp_n.n166 vp_n.n165 13.653
R53582 vp_n.n186 vp_n.n185 13.653
R53583 vp_n.n206 vp_n.n205 13.653
R53584 vp_n.n226 vp_n.n225 13.653
R53585 vp_n.n246 vp_n.n245 13.653
R53586 vp_n.n266 vp_n.n265 13.653
R53587 vp_n.n286 vp_n.n285 13.653
R53588 vp_n.n306 vp_n.n305 13.653
R53589 vp_n.n326 vp_n.n325 13.653
R53590 vp_n.n346 vp_n.n345 13.653
R53591 vp_n.n366 vp_n.n365 13.653
R53592 vp_n.n386 vp_n.n385 13.653
R53593 vp_n.n406 vp_n.n405 13.653
R53594 vp_n.n426 vp_n.n425 13.653
R53595 vp_n.n446 vp_n.n445 13.653
R53596 vp_n.n466 vp_n.n465 13.653
R53597 vp_n.n486 vp_n.n485 13.653
R53598 vp_n.n506 vp_n.n505 13.653
R53599 vp_n.n526 vp_n.n525 13.653
R53600 vp_n.n546 vp_n.n545 13.653
R53601 vp_n.n566 vp_n.n565 13.653
R53602 vp_n.n586 vp_n.n585 13.653
R53603 vp_n.n606 vp_n.n605 13.653
R53604 vp_n.n626 vp_n.n625 13.653
R53605 vp_n.n646 vp_n.n645 13.653
R53606 vp_n.n666 vp_n.n665 13.653
R53607 vp_n.n686 vp_n.n685 13.653
R53608 vp_n.n706 vp_n.n705 13.653
R53609 vp_n.n726 vp_n.n725 13.653
R53610 vp_n.n746 vp_n.n745 13.653
R53611 vp_n.n766 vp_n.n765 13.653
R53612 vp_n.n786 vp_n.n785 13.653
R53613 vp_n.n806 vp_n.n805 13.653
R53614 vp_n.n826 vp_n.n825 13.653
R53615 vp_n.n846 vp_n.n845 13.653
R53616 vp_n.n866 vp_n.n865 13.653
R53617 vp_n.n886 vp_n.n885 13.653
R53618 vp_n.n906 vp_n.n905 13.653
R53619 vp_n.n926 vp_n.n925 13.653
R53620 vp_n.n946 vp_n.n945 13.653
R53621 vp_n.n966 vp_n.n965 13.653
R53622 vp_n.n986 vp_n.n985 13.653
R53623 vp_n.n1006 vp_n.n1005 13.653
R53624 vp_n.n1026 vp_n.n1025 13.653
R53625 vp_n.n1046 vp_n.n1045 13.653
R53626 vp_n.n1066 vp_n.n1065 13.653
R53627 vp_n.n1086 vp_n.n1085 13.653
R53628 vp_n.n1106 vp_n.n1105 13.653
R53629 vp_n.n1126 vp_n.n1125 13.653
R53630 vp_n.n1146 vp_n.n1145 13.653
R53631 vp_n.n1166 vp_n.n1165 13.653
R53632 vp_n.n1186 vp_n.n1185 13.653
R53633 vp_n.n1206 vp_n.n1205 13.653
R53634 vp_n.n1226 vp_n.n1225 13.653
R53635 vp_n.n1246 vp_n.n1245 13.653
R53636 vp_n.n1266 vp_n.n1265 13.653
R53637 vp_n.n1286 vp_n.n1285 13.653
R53638 vp_n.n1306 vp_n.n1305 13.653
R53639 vp_n.n1326 vp_n.n1325 13.653
R53640 vp_n.n1346 vp_n.n1345 13.653
R53641 vp_n.n1366 vp_n.n1365 13.653
R53642 vp_n.n1386 vp_n.n1385 13.653
R53643 vp_n.n1406 vp_n.n1405 13.653
R53644 vp_n.n1426 vp_n.n1425 13.653
R53645 vp_n.n1446 vp_n.n1445 13.653
R53646 vp_n.n1466 vp_n.n1465 13.653
R53647 vp_n.n1486 vp_n.n1485 13.653
R53648 vp_n.n4697 vp_n.n4696 13.653
R53649 vp_n.n1496 vp_n.n1495 13.653
R53650 vp_n.n1493 vp_n.n1492 13.653
R53651 vp_n.n3047 vp_n.n3046 13.653
R53652 vp_n.n1577 vp_n.n1576 13.653
R53653 vp_n.n1584 vp_n.n1583 13.653
R53654 vp_n.n1597 vp_n.n1596 13.653
R53655 vp_n.n1604 vp_n.n1603 13.653
R53656 vp_n.n1617 vp_n.n1616 13.653
R53657 vp_n.n1624 vp_n.n1623 13.653
R53658 vp_n.n1637 vp_n.n1636 13.653
R53659 vp_n.n1644 vp_n.n1643 13.653
R53660 vp_n.n1657 vp_n.n1656 13.653
R53661 vp_n.n1664 vp_n.n1663 13.653
R53662 vp_n.n1677 vp_n.n1676 13.653
R53663 vp_n.n1684 vp_n.n1683 13.653
R53664 vp_n.n1697 vp_n.n1696 13.653
R53665 vp_n.n1704 vp_n.n1703 13.653
R53666 vp_n.n1717 vp_n.n1716 13.653
R53667 vp_n.n1724 vp_n.n1723 13.653
R53668 vp_n.n1737 vp_n.n1736 13.653
R53669 vp_n.n1744 vp_n.n1743 13.653
R53670 vp_n.n1757 vp_n.n1756 13.653
R53671 vp_n.n1764 vp_n.n1763 13.653
R53672 vp_n.n1777 vp_n.n1776 13.653
R53673 vp_n.n1784 vp_n.n1783 13.653
R53674 vp_n.n1797 vp_n.n1796 13.653
R53675 vp_n.n1804 vp_n.n1803 13.653
R53676 vp_n.n1817 vp_n.n1816 13.653
R53677 vp_n.n1824 vp_n.n1823 13.653
R53678 vp_n.n1837 vp_n.n1836 13.653
R53679 vp_n.n1844 vp_n.n1843 13.653
R53680 vp_n.n1857 vp_n.n1856 13.653
R53681 vp_n.n1864 vp_n.n1863 13.653
R53682 vp_n.n1877 vp_n.n1876 13.653
R53683 vp_n.n1884 vp_n.n1883 13.653
R53684 vp_n.n1897 vp_n.n1896 13.653
R53685 vp_n.n1904 vp_n.n1903 13.653
R53686 vp_n.n1917 vp_n.n1916 13.653
R53687 vp_n.n1924 vp_n.n1923 13.653
R53688 vp_n.n1937 vp_n.n1936 13.653
R53689 vp_n.n1944 vp_n.n1943 13.653
R53690 vp_n.n1957 vp_n.n1956 13.653
R53691 vp_n.n1964 vp_n.n1963 13.653
R53692 vp_n.n1977 vp_n.n1976 13.653
R53693 vp_n.n1984 vp_n.n1983 13.653
R53694 vp_n.n1997 vp_n.n1996 13.653
R53695 vp_n.n2004 vp_n.n2003 13.653
R53696 vp_n.n2017 vp_n.n2016 13.653
R53697 vp_n.n2024 vp_n.n2023 13.653
R53698 vp_n.n2037 vp_n.n2036 13.653
R53699 vp_n.n2044 vp_n.n2043 13.653
R53700 vp_n.n2057 vp_n.n2056 13.653
R53701 vp_n.n2064 vp_n.n2063 13.653
R53702 vp_n.n2077 vp_n.n2076 13.653
R53703 vp_n.n2084 vp_n.n2083 13.653
R53704 vp_n.n2097 vp_n.n2096 13.653
R53705 vp_n.n2104 vp_n.n2103 13.653
R53706 vp_n.n2117 vp_n.n2116 13.653
R53707 vp_n.n2124 vp_n.n2123 13.653
R53708 vp_n.n2137 vp_n.n2136 13.653
R53709 vp_n.n2144 vp_n.n2143 13.653
R53710 vp_n.n2157 vp_n.n2156 13.653
R53711 vp_n.n2164 vp_n.n2163 13.653
R53712 vp_n.n2177 vp_n.n2176 13.653
R53713 vp_n.n2184 vp_n.n2183 13.653
R53714 vp_n.n2197 vp_n.n2196 13.653
R53715 vp_n.n2204 vp_n.n2203 13.653
R53716 vp_n.n2217 vp_n.n2216 13.653
R53717 vp_n.n2224 vp_n.n2223 13.653
R53718 vp_n.n2237 vp_n.n2236 13.653
R53719 vp_n.n2244 vp_n.n2243 13.653
R53720 vp_n.n2257 vp_n.n2256 13.653
R53721 vp_n.n2264 vp_n.n2263 13.653
R53722 vp_n.n2277 vp_n.n2276 13.653
R53723 vp_n.n2284 vp_n.n2283 13.653
R53724 vp_n.n2297 vp_n.n2296 13.653
R53725 vp_n.n2304 vp_n.n2303 13.653
R53726 vp_n.n2317 vp_n.n2316 13.653
R53727 vp_n.n2324 vp_n.n2323 13.653
R53728 vp_n.n2337 vp_n.n2336 13.653
R53729 vp_n.n2344 vp_n.n2343 13.653
R53730 vp_n.n2357 vp_n.n2356 13.653
R53731 vp_n.n2364 vp_n.n2363 13.653
R53732 vp_n.n2377 vp_n.n2376 13.653
R53733 vp_n.n2384 vp_n.n2383 13.653
R53734 vp_n.n2397 vp_n.n2396 13.653
R53735 vp_n.n2404 vp_n.n2403 13.653
R53736 vp_n.n2417 vp_n.n2416 13.653
R53737 vp_n.n2424 vp_n.n2423 13.653
R53738 vp_n.n2437 vp_n.n2436 13.653
R53739 vp_n.n2444 vp_n.n2443 13.653
R53740 vp_n.n2457 vp_n.n2456 13.653
R53741 vp_n.n2464 vp_n.n2463 13.653
R53742 vp_n.n2477 vp_n.n2476 13.653
R53743 vp_n.n2484 vp_n.n2483 13.653
R53744 vp_n.n2497 vp_n.n2496 13.653
R53745 vp_n.n2504 vp_n.n2503 13.653
R53746 vp_n.n2517 vp_n.n2516 13.653
R53747 vp_n.n2524 vp_n.n2523 13.653
R53748 vp_n.n2537 vp_n.n2536 13.653
R53749 vp_n.n2544 vp_n.n2543 13.653
R53750 vp_n.n2557 vp_n.n2556 13.653
R53751 vp_n.n2564 vp_n.n2563 13.653
R53752 vp_n.n2577 vp_n.n2576 13.653
R53753 vp_n.n2584 vp_n.n2583 13.653
R53754 vp_n.n2597 vp_n.n2596 13.653
R53755 vp_n.n2604 vp_n.n2603 13.653
R53756 vp_n.n2617 vp_n.n2616 13.653
R53757 vp_n.n2624 vp_n.n2623 13.653
R53758 vp_n.n2637 vp_n.n2636 13.653
R53759 vp_n.n2644 vp_n.n2643 13.653
R53760 vp_n.n2657 vp_n.n2656 13.653
R53761 vp_n.n2664 vp_n.n2663 13.653
R53762 vp_n.n2677 vp_n.n2676 13.653
R53763 vp_n.n2684 vp_n.n2683 13.653
R53764 vp_n.n2697 vp_n.n2696 13.653
R53765 vp_n.n2704 vp_n.n2703 13.653
R53766 vp_n.n2717 vp_n.n2716 13.653
R53767 vp_n.n2724 vp_n.n2723 13.653
R53768 vp_n.n2737 vp_n.n2736 13.653
R53769 vp_n.n2744 vp_n.n2743 13.653
R53770 vp_n.n2757 vp_n.n2756 13.653
R53771 vp_n.n2764 vp_n.n2763 13.653
R53772 vp_n.n2777 vp_n.n2776 13.653
R53773 vp_n.n2784 vp_n.n2783 13.653
R53774 vp_n.n2797 vp_n.n2796 13.653
R53775 vp_n.n2804 vp_n.n2803 13.653
R53776 vp_n.n2817 vp_n.n2816 13.653
R53777 vp_n.n2824 vp_n.n2823 13.653
R53778 vp_n.n2837 vp_n.n2836 13.653
R53779 vp_n.n2844 vp_n.n2843 13.653
R53780 vp_n.n2857 vp_n.n2856 13.653
R53781 vp_n.n2864 vp_n.n2863 13.653
R53782 vp_n.n2877 vp_n.n2876 13.653
R53783 vp_n.n2884 vp_n.n2883 13.653
R53784 vp_n.n2897 vp_n.n2896 13.653
R53785 vp_n.n2904 vp_n.n2903 13.653
R53786 vp_n.n2917 vp_n.n2916 13.653
R53787 vp_n.n2924 vp_n.n2923 13.653
R53788 vp_n.n2937 vp_n.n2936 13.653
R53789 vp_n.n2944 vp_n.n2943 13.653
R53790 vp_n.n2957 vp_n.n2956 13.653
R53791 vp_n.n2964 vp_n.n2963 13.653
R53792 vp_n.n2977 vp_n.n2976 13.653
R53793 vp_n.n2984 vp_n.n2983 13.653
R53794 vp_n.n2997 vp_n.n2996 13.653
R53795 vp_n.n3004 vp_n.n3003 13.653
R53796 vp_n.n3017 vp_n.n3016 13.653
R53797 vp_n.n3024 vp_n.n3023 13.653
R53798 vp_n.n3037 vp_n.n3036 13.653
R53799 vp_n.n3044 vp_n.n3043 13.653
R53800 vp_n.n1567 vp_n.n1566 13.653
R53801 vp_n.n1564 vp_n.n1563 13.653
R53802 vp_n.n13 vp_n.n12 13.653
R53803 vp_n.n16 vp_n.n15 13.653
R53804 vp_n.n3220 vp_n.n3219 13.653
R53805 vp_n.n3217 vp_n.n3216 13.653
R53806 vp_n.n4700 vp_n.n4699 13.653
R53807 vp_n.n4690 vp_n.n4689 13.653
R53808 vp_n.n4677 vp_n.n4676 13.653
R53809 vp_n.n4670 vp_n.n4669 13.653
R53810 vp_n.n4657 vp_n.n4656 13.653
R53811 vp_n.n4650 vp_n.n4649 13.653
R53812 vp_n.n4637 vp_n.n4636 13.653
R53813 vp_n.n4630 vp_n.n4629 13.653
R53814 vp_n.n4617 vp_n.n4616 13.653
R53815 vp_n.n4610 vp_n.n4609 13.653
R53816 vp_n.n4597 vp_n.n4596 13.653
R53817 vp_n.n4590 vp_n.n4589 13.653
R53818 vp_n.n4577 vp_n.n4576 13.653
R53819 vp_n.n4570 vp_n.n4569 13.653
R53820 vp_n.n4557 vp_n.n4556 13.653
R53821 vp_n.n4550 vp_n.n4549 13.653
R53822 vp_n.n4537 vp_n.n4536 13.653
R53823 vp_n.n4530 vp_n.n4529 13.653
R53824 vp_n.n4517 vp_n.n4516 13.653
R53825 vp_n.n4510 vp_n.n4509 13.653
R53826 vp_n.n4497 vp_n.n4496 13.653
R53827 vp_n.n4490 vp_n.n4489 13.653
R53828 vp_n.n4477 vp_n.n4476 13.653
R53829 vp_n.n4470 vp_n.n4469 13.653
R53830 vp_n.n4457 vp_n.n4456 13.653
R53831 vp_n.n4450 vp_n.n4449 13.653
R53832 vp_n.n4437 vp_n.n4436 13.653
R53833 vp_n.n4430 vp_n.n4429 13.653
R53834 vp_n.n4417 vp_n.n4416 13.653
R53835 vp_n.n4410 vp_n.n4409 13.653
R53836 vp_n.n4397 vp_n.n4396 13.653
R53837 vp_n.n4390 vp_n.n4389 13.653
R53838 vp_n.n4377 vp_n.n4376 13.653
R53839 vp_n.n4370 vp_n.n4369 13.653
R53840 vp_n.n4357 vp_n.n4356 13.653
R53841 vp_n.n4350 vp_n.n4349 13.653
R53842 vp_n.n4337 vp_n.n4336 13.653
R53843 vp_n.n4330 vp_n.n4329 13.653
R53844 vp_n.n4317 vp_n.n4316 13.653
R53845 vp_n.n4310 vp_n.n4309 13.653
R53846 vp_n.n4297 vp_n.n4296 13.653
R53847 vp_n.n4290 vp_n.n4289 13.653
R53848 vp_n.n4277 vp_n.n4276 13.653
R53849 vp_n.n4270 vp_n.n4269 13.653
R53850 vp_n.n4257 vp_n.n4256 13.653
R53851 vp_n.n4250 vp_n.n4249 13.653
R53852 vp_n.n4237 vp_n.n4236 13.653
R53853 vp_n.n4230 vp_n.n4229 13.653
R53854 vp_n.n4217 vp_n.n4216 13.653
R53855 vp_n.n4210 vp_n.n4209 13.653
R53856 vp_n.n4197 vp_n.n4196 13.653
R53857 vp_n.n4190 vp_n.n4189 13.653
R53858 vp_n.n4177 vp_n.n4176 13.653
R53859 vp_n.n4170 vp_n.n4169 13.653
R53860 vp_n.n4157 vp_n.n4156 13.653
R53861 vp_n.n4150 vp_n.n4149 13.653
R53862 vp_n.n4137 vp_n.n4136 13.653
R53863 vp_n.n4130 vp_n.n4129 13.653
R53864 vp_n.n4117 vp_n.n4116 13.653
R53865 vp_n.n4110 vp_n.n4109 13.653
R53866 vp_n.n4097 vp_n.n4096 13.653
R53867 vp_n.n4090 vp_n.n4089 13.653
R53868 vp_n.n4077 vp_n.n4076 13.653
R53869 vp_n.n4070 vp_n.n4069 13.653
R53870 vp_n.n4057 vp_n.n4056 13.653
R53871 vp_n.n4050 vp_n.n4049 13.653
R53872 vp_n.n4037 vp_n.n4036 13.653
R53873 vp_n.n4030 vp_n.n4029 13.653
R53874 vp_n.n4017 vp_n.n4016 13.653
R53875 vp_n.n4010 vp_n.n4009 13.653
R53876 vp_n.n3997 vp_n.n3996 13.653
R53877 vp_n.n3990 vp_n.n3989 13.653
R53878 vp_n.n3977 vp_n.n3976 13.653
R53879 vp_n.n3970 vp_n.n3969 13.653
R53880 vp_n.n3957 vp_n.n3956 13.653
R53881 vp_n.n3950 vp_n.n3949 13.653
R53882 vp_n.n3937 vp_n.n3936 13.653
R53883 vp_n.n3930 vp_n.n3929 13.653
R53884 vp_n.n3917 vp_n.n3916 13.653
R53885 vp_n.n3910 vp_n.n3909 13.653
R53886 vp_n.n3897 vp_n.n3896 13.653
R53887 vp_n.n3890 vp_n.n3889 13.653
R53888 vp_n.n3877 vp_n.n3876 13.653
R53889 vp_n.n3870 vp_n.n3869 13.653
R53890 vp_n.n3857 vp_n.n3856 13.653
R53891 vp_n.n3850 vp_n.n3849 13.653
R53892 vp_n.n3837 vp_n.n3836 13.653
R53893 vp_n.n3830 vp_n.n3829 13.653
R53894 vp_n.n3817 vp_n.n3816 13.653
R53895 vp_n.n3810 vp_n.n3809 13.653
R53896 vp_n.n3797 vp_n.n3796 13.653
R53897 vp_n.n3790 vp_n.n3789 13.653
R53898 vp_n.n3777 vp_n.n3776 13.653
R53899 vp_n.n3770 vp_n.n3769 13.653
R53900 vp_n.n3757 vp_n.n3756 13.653
R53901 vp_n.n3750 vp_n.n3749 13.653
R53902 vp_n.n3737 vp_n.n3736 13.653
R53903 vp_n.n3730 vp_n.n3729 13.653
R53904 vp_n.n3717 vp_n.n3716 13.653
R53905 vp_n.n3710 vp_n.n3709 13.653
R53906 vp_n.n3697 vp_n.n3696 13.653
R53907 vp_n.n3690 vp_n.n3689 13.653
R53908 vp_n.n3677 vp_n.n3676 13.653
R53909 vp_n.n3670 vp_n.n3669 13.653
R53910 vp_n.n3657 vp_n.n3656 13.653
R53911 vp_n.n3650 vp_n.n3649 13.653
R53912 vp_n.n3637 vp_n.n3636 13.653
R53913 vp_n.n3630 vp_n.n3629 13.653
R53914 vp_n.n3617 vp_n.n3616 13.653
R53915 vp_n.n3610 vp_n.n3609 13.653
R53916 vp_n.n3597 vp_n.n3596 13.653
R53917 vp_n.n3590 vp_n.n3589 13.653
R53918 vp_n.n3577 vp_n.n3576 13.653
R53919 vp_n.n3570 vp_n.n3569 13.653
R53920 vp_n.n3557 vp_n.n3556 13.653
R53921 vp_n.n3550 vp_n.n3549 13.653
R53922 vp_n.n3537 vp_n.n3536 13.653
R53923 vp_n.n3530 vp_n.n3529 13.653
R53924 vp_n.n3517 vp_n.n3516 13.653
R53925 vp_n.n3510 vp_n.n3509 13.653
R53926 vp_n.n3497 vp_n.n3496 13.653
R53927 vp_n.n3490 vp_n.n3489 13.653
R53928 vp_n.n3477 vp_n.n3476 13.653
R53929 vp_n.n3470 vp_n.n3469 13.653
R53930 vp_n.n3457 vp_n.n3456 13.653
R53931 vp_n.n3450 vp_n.n3449 13.653
R53932 vp_n.n3437 vp_n.n3436 13.653
R53933 vp_n.n3430 vp_n.n3429 13.653
R53934 vp_n.n3417 vp_n.n3416 13.653
R53935 vp_n.n3410 vp_n.n3409 13.653
R53936 vp_n.n3397 vp_n.n3396 13.653
R53937 vp_n.n3390 vp_n.n3389 13.653
R53938 vp_n.n3377 vp_n.n3376 13.653
R53939 vp_n.n3370 vp_n.n3369 13.653
R53940 vp_n.n3357 vp_n.n3356 13.653
R53941 vp_n.n3350 vp_n.n3349 13.653
R53942 vp_n.n3337 vp_n.n3336 13.653
R53943 vp_n.n3330 vp_n.n3329 13.653
R53944 vp_n.n3317 vp_n.n3316 13.653
R53945 vp_n.n3310 vp_n.n3309 13.653
R53946 vp_n.n3297 vp_n.n3296 13.653
R53947 vp_n.n3290 vp_n.n3289 13.653
R53948 vp_n.n3277 vp_n.n3276 13.653
R53949 vp_n.n3270 vp_n.n3269 13.653
R53950 vp_n.n3257 vp_n.n3256 13.653
R53951 vp_n.n3250 vp_n.n3249 13.653
R53952 vp_n.n3237 vp_n.n3236 13.653
R53953 vp_n.n3230 vp_n.n3229 13.653
R53954 vp_n.n3207 vp_n.n3206 13.653
R53955 vp_n.n3210 vp_n.n3209 13.653
R53956 vp_n.n3 vp_n.n2 13.653
R53957 vp_n.n6 vp_n.n5 13.653
R53958 vp_n.n1554 vp_n.n1553 13.653
R53959 vp_n.n1557 vp_n.n1556 13.653
R53960 vp_n.n1559 vp_n.n1558 12.877
R53961 vp_n.n8 vp_n.n7 12.877
R53962 vp_n.n18 vp_n.n17 12.877
R53963 vp_n.n1579 vp_n.n1578 12.877
R53964 vp_n.n3232 vp_n.n3231 12.877
R53965 vp_n.n28 vp_n.n27 12.877
R53966 vp_n.n1589 vp_n.n1588 12.877
R53967 vp_n.n3242 vp_n.n3241 12.877
R53968 vp_n.n38 vp_n.n37 12.877
R53969 vp_n.n1599 vp_n.n1598 12.877
R53970 vp_n.n3252 vp_n.n3251 12.877
R53971 vp_n.n48 vp_n.n47 12.877
R53972 vp_n.n1609 vp_n.n1608 12.877
R53973 vp_n.n3262 vp_n.n3261 12.877
R53974 vp_n.n58 vp_n.n57 12.877
R53975 vp_n.n1619 vp_n.n1618 12.877
R53976 vp_n.n3272 vp_n.n3271 12.877
R53977 vp_n.n68 vp_n.n67 12.877
R53978 vp_n.n1629 vp_n.n1628 12.877
R53979 vp_n.n3282 vp_n.n3281 12.877
R53980 vp_n.n78 vp_n.n77 12.877
R53981 vp_n.n1639 vp_n.n1638 12.877
R53982 vp_n.n3292 vp_n.n3291 12.877
R53983 vp_n.n88 vp_n.n87 12.877
R53984 vp_n.n1649 vp_n.n1648 12.877
R53985 vp_n.n3302 vp_n.n3301 12.877
R53986 vp_n.n98 vp_n.n97 12.877
R53987 vp_n.n1659 vp_n.n1658 12.877
R53988 vp_n.n3312 vp_n.n3311 12.877
R53989 vp_n.n108 vp_n.n107 12.877
R53990 vp_n.n1669 vp_n.n1668 12.877
R53991 vp_n.n3322 vp_n.n3321 12.877
R53992 vp_n.n118 vp_n.n117 12.877
R53993 vp_n.n1679 vp_n.n1678 12.877
R53994 vp_n.n3332 vp_n.n3331 12.877
R53995 vp_n.n128 vp_n.n127 12.877
R53996 vp_n.n1689 vp_n.n1688 12.877
R53997 vp_n.n3342 vp_n.n3341 12.877
R53998 vp_n.n138 vp_n.n137 12.877
R53999 vp_n.n1699 vp_n.n1698 12.877
R54000 vp_n.n3352 vp_n.n3351 12.877
R54001 vp_n.n148 vp_n.n147 12.877
R54002 vp_n.n1709 vp_n.n1708 12.877
R54003 vp_n.n3362 vp_n.n3361 12.877
R54004 vp_n.n158 vp_n.n157 12.877
R54005 vp_n.n1719 vp_n.n1718 12.877
R54006 vp_n.n3372 vp_n.n3371 12.877
R54007 vp_n.n168 vp_n.n167 12.877
R54008 vp_n.n1729 vp_n.n1728 12.877
R54009 vp_n.n3382 vp_n.n3381 12.877
R54010 vp_n.n178 vp_n.n177 12.877
R54011 vp_n.n1739 vp_n.n1738 12.877
R54012 vp_n.n3392 vp_n.n3391 12.877
R54013 vp_n.n188 vp_n.n187 12.877
R54014 vp_n.n1749 vp_n.n1748 12.877
R54015 vp_n.n3402 vp_n.n3401 12.877
R54016 vp_n.n198 vp_n.n197 12.877
R54017 vp_n.n1759 vp_n.n1758 12.877
R54018 vp_n.n3412 vp_n.n3411 12.877
R54019 vp_n.n208 vp_n.n207 12.877
R54020 vp_n.n1769 vp_n.n1768 12.877
R54021 vp_n.n3422 vp_n.n3421 12.877
R54022 vp_n.n218 vp_n.n217 12.877
R54023 vp_n.n1779 vp_n.n1778 12.877
R54024 vp_n.n3432 vp_n.n3431 12.877
R54025 vp_n.n228 vp_n.n227 12.877
R54026 vp_n.n1789 vp_n.n1788 12.877
R54027 vp_n.n3442 vp_n.n3441 12.877
R54028 vp_n.n238 vp_n.n237 12.877
R54029 vp_n.n1799 vp_n.n1798 12.877
R54030 vp_n.n3452 vp_n.n3451 12.877
R54031 vp_n.n248 vp_n.n247 12.877
R54032 vp_n.n1809 vp_n.n1808 12.877
R54033 vp_n.n3462 vp_n.n3461 12.877
R54034 vp_n.n258 vp_n.n257 12.877
R54035 vp_n.n1819 vp_n.n1818 12.877
R54036 vp_n.n3472 vp_n.n3471 12.877
R54037 vp_n.n268 vp_n.n267 12.877
R54038 vp_n.n1829 vp_n.n1828 12.877
R54039 vp_n.n3482 vp_n.n3481 12.877
R54040 vp_n.n278 vp_n.n277 12.877
R54041 vp_n.n1839 vp_n.n1838 12.877
R54042 vp_n.n3492 vp_n.n3491 12.877
R54043 vp_n.n288 vp_n.n287 12.877
R54044 vp_n.n1849 vp_n.n1848 12.877
R54045 vp_n.n3502 vp_n.n3501 12.877
R54046 vp_n.n298 vp_n.n297 12.877
R54047 vp_n.n1859 vp_n.n1858 12.877
R54048 vp_n.n3512 vp_n.n3511 12.877
R54049 vp_n.n308 vp_n.n307 12.877
R54050 vp_n.n1869 vp_n.n1868 12.877
R54051 vp_n.n3522 vp_n.n3521 12.877
R54052 vp_n.n318 vp_n.n317 12.877
R54053 vp_n.n1879 vp_n.n1878 12.877
R54054 vp_n.n3532 vp_n.n3531 12.877
R54055 vp_n.n328 vp_n.n327 12.877
R54056 vp_n.n1889 vp_n.n1888 12.877
R54057 vp_n.n3542 vp_n.n3541 12.877
R54058 vp_n.n338 vp_n.n337 12.877
R54059 vp_n.n1899 vp_n.n1898 12.877
R54060 vp_n.n3552 vp_n.n3551 12.877
R54061 vp_n.n348 vp_n.n347 12.877
R54062 vp_n.n1909 vp_n.n1908 12.877
R54063 vp_n.n3562 vp_n.n3561 12.877
R54064 vp_n.n358 vp_n.n357 12.877
R54065 vp_n.n1919 vp_n.n1918 12.877
R54066 vp_n.n3572 vp_n.n3571 12.877
R54067 vp_n.n368 vp_n.n367 12.877
R54068 vp_n.n1929 vp_n.n1928 12.877
R54069 vp_n.n3582 vp_n.n3581 12.877
R54070 vp_n.n378 vp_n.n377 12.877
R54071 vp_n.n1939 vp_n.n1938 12.877
R54072 vp_n.n3592 vp_n.n3591 12.877
R54073 vp_n.n388 vp_n.n387 12.877
R54074 vp_n.n1949 vp_n.n1948 12.877
R54075 vp_n.n3602 vp_n.n3601 12.877
R54076 vp_n.n398 vp_n.n397 12.877
R54077 vp_n.n1959 vp_n.n1958 12.877
R54078 vp_n.n3612 vp_n.n3611 12.877
R54079 vp_n.n408 vp_n.n407 12.877
R54080 vp_n.n1969 vp_n.n1968 12.877
R54081 vp_n.n3622 vp_n.n3621 12.877
R54082 vp_n.n418 vp_n.n417 12.877
R54083 vp_n.n1979 vp_n.n1978 12.877
R54084 vp_n.n3632 vp_n.n3631 12.877
R54085 vp_n.n428 vp_n.n427 12.877
R54086 vp_n.n1989 vp_n.n1988 12.877
R54087 vp_n.n3642 vp_n.n3641 12.877
R54088 vp_n.n438 vp_n.n437 12.877
R54089 vp_n.n1999 vp_n.n1998 12.877
R54090 vp_n.n3652 vp_n.n3651 12.877
R54091 vp_n.n448 vp_n.n447 12.877
R54092 vp_n.n2009 vp_n.n2008 12.877
R54093 vp_n.n3662 vp_n.n3661 12.877
R54094 vp_n.n458 vp_n.n457 12.877
R54095 vp_n.n2019 vp_n.n2018 12.877
R54096 vp_n.n3672 vp_n.n3671 12.877
R54097 vp_n.n468 vp_n.n467 12.877
R54098 vp_n.n2029 vp_n.n2028 12.877
R54099 vp_n.n3682 vp_n.n3681 12.877
R54100 vp_n.n478 vp_n.n477 12.877
R54101 vp_n.n2039 vp_n.n2038 12.877
R54102 vp_n.n3692 vp_n.n3691 12.877
R54103 vp_n.n488 vp_n.n487 12.877
R54104 vp_n.n2049 vp_n.n2048 12.877
R54105 vp_n.n3702 vp_n.n3701 12.877
R54106 vp_n.n498 vp_n.n497 12.877
R54107 vp_n.n2059 vp_n.n2058 12.877
R54108 vp_n.n3712 vp_n.n3711 12.877
R54109 vp_n.n508 vp_n.n507 12.877
R54110 vp_n.n2069 vp_n.n2068 12.877
R54111 vp_n.n3722 vp_n.n3721 12.877
R54112 vp_n.n518 vp_n.n517 12.877
R54113 vp_n.n2079 vp_n.n2078 12.877
R54114 vp_n.n3732 vp_n.n3731 12.877
R54115 vp_n.n528 vp_n.n527 12.877
R54116 vp_n.n2089 vp_n.n2088 12.877
R54117 vp_n.n3742 vp_n.n3741 12.877
R54118 vp_n.n538 vp_n.n537 12.877
R54119 vp_n.n2099 vp_n.n2098 12.877
R54120 vp_n.n3752 vp_n.n3751 12.877
R54121 vp_n.n548 vp_n.n547 12.877
R54122 vp_n.n2109 vp_n.n2108 12.877
R54123 vp_n.n3762 vp_n.n3761 12.877
R54124 vp_n.n558 vp_n.n557 12.877
R54125 vp_n.n2119 vp_n.n2118 12.877
R54126 vp_n.n3772 vp_n.n3771 12.877
R54127 vp_n.n568 vp_n.n567 12.877
R54128 vp_n.n2129 vp_n.n2128 12.877
R54129 vp_n.n3782 vp_n.n3781 12.877
R54130 vp_n.n578 vp_n.n577 12.877
R54131 vp_n.n2139 vp_n.n2138 12.877
R54132 vp_n.n3792 vp_n.n3791 12.877
R54133 vp_n.n588 vp_n.n587 12.877
R54134 vp_n.n2149 vp_n.n2148 12.877
R54135 vp_n.n3802 vp_n.n3801 12.877
R54136 vp_n.n598 vp_n.n597 12.877
R54137 vp_n.n2159 vp_n.n2158 12.877
R54138 vp_n.n3812 vp_n.n3811 12.877
R54139 vp_n.n608 vp_n.n607 12.877
R54140 vp_n.n2169 vp_n.n2168 12.877
R54141 vp_n.n3822 vp_n.n3821 12.877
R54142 vp_n.n618 vp_n.n617 12.877
R54143 vp_n.n2179 vp_n.n2178 12.877
R54144 vp_n.n3832 vp_n.n3831 12.877
R54145 vp_n.n628 vp_n.n627 12.877
R54146 vp_n.n2189 vp_n.n2188 12.877
R54147 vp_n.n3842 vp_n.n3841 12.877
R54148 vp_n.n638 vp_n.n637 12.877
R54149 vp_n.n2199 vp_n.n2198 12.877
R54150 vp_n.n3852 vp_n.n3851 12.877
R54151 vp_n.n648 vp_n.n647 12.877
R54152 vp_n.n2209 vp_n.n2208 12.877
R54153 vp_n.n3862 vp_n.n3861 12.877
R54154 vp_n.n658 vp_n.n657 12.877
R54155 vp_n.n2219 vp_n.n2218 12.877
R54156 vp_n.n3872 vp_n.n3871 12.877
R54157 vp_n.n668 vp_n.n667 12.877
R54158 vp_n.n2229 vp_n.n2228 12.877
R54159 vp_n.n3882 vp_n.n3881 12.877
R54160 vp_n.n678 vp_n.n677 12.877
R54161 vp_n.n2239 vp_n.n2238 12.877
R54162 vp_n.n3892 vp_n.n3891 12.877
R54163 vp_n.n688 vp_n.n687 12.877
R54164 vp_n.n2249 vp_n.n2248 12.877
R54165 vp_n.n3902 vp_n.n3901 12.877
R54166 vp_n.n698 vp_n.n697 12.877
R54167 vp_n.n2259 vp_n.n2258 12.877
R54168 vp_n.n3912 vp_n.n3911 12.877
R54169 vp_n.n708 vp_n.n707 12.877
R54170 vp_n.n2269 vp_n.n2268 12.877
R54171 vp_n.n3922 vp_n.n3921 12.877
R54172 vp_n.n718 vp_n.n717 12.877
R54173 vp_n.n2279 vp_n.n2278 12.877
R54174 vp_n.n3932 vp_n.n3931 12.877
R54175 vp_n.n728 vp_n.n727 12.877
R54176 vp_n.n2289 vp_n.n2288 12.877
R54177 vp_n.n3942 vp_n.n3941 12.877
R54178 vp_n.n738 vp_n.n737 12.877
R54179 vp_n.n2299 vp_n.n2298 12.877
R54180 vp_n.n3952 vp_n.n3951 12.877
R54181 vp_n.n748 vp_n.n747 12.877
R54182 vp_n.n2309 vp_n.n2308 12.877
R54183 vp_n.n3962 vp_n.n3961 12.877
R54184 vp_n.n758 vp_n.n757 12.877
R54185 vp_n.n2319 vp_n.n2318 12.877
R54186 vp_n.n3972 vp_n.n3971 12.877
R54187 vp_n.n768 vp_n.n767 12.877
R54188 vp_n.n2329 vp_n.n2328 12.877
R54189 vp_n.n3982 vp_n.n3981 12.877
R54190 vp_n.n778 vp_n.n777 12.877
R54191 vp_n.n2339 vp_n.n2338 12.877
R54192 vp_n.n3992 vp_n.n3991 12.877
R54193 vp_n.n788 vp_n.n787 12.877
R54194 vp_n.n2349 vp_n.n2348 12.877
R54195 vp_n.n4002 vp_n.n4001 12.877
R54196 vp_n.n798 vp_n.n797 12.877
R54197 vp_n.n2359 vp_n.n2358 12.877
R54198 vp_n.n4012 vp_n.n4011 12.877
R54199 vp_n.n808 vp_n.n807 12.877
R54200 vp_n.n2369 vp_n.n2368 12.877
R54201 vp_n.n4022 vp_n.n4021 12.877
R54202 vp_n.n818 vp_n.n817 12.877
R54203 vp_n.n2379 vp_n.n2378 12.877
R54204 vp_n.n4032 vp_n.n4031 12.877
R54205 vp_n.n828 vp_n.n827 12.877
R54206 vp_n.n2389 vp_n.n2388 12.877
R54207 vp_n.n4042 vp_n.n4041 12.877
R54208 vp_n.n838 vp_n.n837 12.877
R54209 vp_n.n2399 vp_n.n2398 12.877
R54210 vp_n.n4052 vp_n.n4051 12.877
R54211 vp_n.n848 vp_n.n847 12.877
R54212 vp_n.n2409 vp_n.n2408 12.877
R54213 vp_n.n4062 vp_n.n4061 12.877
R54214 vp_n.n858 vp_n.n857 12.877
R54215 vp_n.n2419 vp_n.n2418 12.877
R54216 vp_n.n4072 vp_n.n4071 12.877
R54217 vp_n.n868 vp_n.n867 12.877
R54218 vp_n.n2429 vp_n.n2428 12.877
R54219 vp_n.n4082 vp_n.n4081 12.877
R54220 vp_n.n878 vp_n.n877 12.877
R54221 vp_n.n2439 vp_n.n2438 12.877
R54222 vp_n.n4092 vp_n.n4091 12.877
R54223 vp_n.n888 vp_n.n887 12.877
R54224 vp_n.n2449 vp_n.n2448 12.877
R54225 vp_n.n4102 vp_n.n4101 12.877
R54226 vp_n.n898 vp_n.n897 12.877
R54227 vp_n.n2459 vp_n.n2458 12.877
R54228 vp_n.n4112 vp_n.n4111 12.877
R54229 vp_n.n908 vp_n.n907 12.877
R54230 vp_n.n2469 vp_n.n2468 12.877
R54231 vp_n.n4122 vp_n.n4121 12.877
R54232 vp_n.n918 vp_n.n917 12.877
R54233 vp_n.n2479 vp_n.n2478 12.877
R54234 vp_n.n4132 vp_n.n4131 12.877
R54235 vp_n.n928 vp_n.n927 12.877
R54236 vp_n.n2489 vp_n.n2488 12.877
R54237 vp_n.n4142 vp_n.n4141 12.877
R54238 vp_n.n938 vp_n.n937 12.877
R54239 vp_n.n2499 vp_n.n2498 12.877
R54240 vp_n.n4152 vp_n.n4151 12.877
R54241 vp_n.n948 vp_n.n947 12.877
R54242 vp_n.n2509 vp_n.n2508 12.877
R54243 vp_n.n4162 vp_n.n4161 12.877
R54244 vp_n.n958 vp_n.n957 12.877
R54245 vp_n.n2519 vp_n.n2518 12.877
R54246 vp_n.n4172 vp_n.n4171 12.877
R54247 vp_n.n968 vp_n.n967 12.877
R54248 vp_n.n2529 vp_n.n2528 12.877
R54249 vp_n.n4182 vp_n.n4181 12.877
R54250 vp_n.n978 vp_n.n977 12.877
R54251 vp_n.n2539 vp_n.n2538 12.877
R54252 vp_n.n4192 vp_n.n4191 12.877
R54253 vp_n.n988 vp_n.n987 12.877
R54254 vp_n.n2549 vp_n.n2548 12.877
R54255 vp_n.n4202 vp_n.n4201 12.877
R54256 vp_n.n998 vp_n.n997 12.877
R54257 vp_n.n2559 vp_n.n2558 12.877
R54258 vp_n.n4212 vp_n.n4211 12.877
R54259 vp_n.n1008 vp_n.n1007 12.877
R54260 vp_n.n2569 vp_n.n2568 12.877
R54261 vp_n.n4222 vp_n.n4221 12.877
R54262 vp_n.n1018 vp_n.n1017 12.877
R54263 vp_n.n2579 vp_n.n2578 12.877
R54264 vp_n.n4232 vp_n.n4231 12.877
R54265 vp_n.n1028 vp_n.n1027 12.877
R54266 vp_n.n2589 vp_n.n2588 12.877
R54267 vp_n.n4242 vp_n.n4241 12.877
R54268 vp_n.n1038 vp_n.n1037 12.877
R54269 vp_n.n2599 vp_n.n2598 12.877
R54270 vp_n.n4252 vp_n.n4251 12.877
R54271 vp_n.n1048 vp_n.n1047 12.877
R54272 vp_n.n2609 vp_n.n2608 12.877
R54273 vp_n.n4262 vp_n.n4261 12.877
R54274 vp_n.n1058 vp_n.n1057 12.877
R54275 vp_n.n2619 vp_n.n2618 12.877
R54276 vp_n.n4272 vp_n.n4271 12.877
R54277 vp_n.n1068 vp_n.n1067 12.877
R54278 vp_n.n2629 vp_n.n2628 12.877
R54279 vp_n.n4282 vp_n.n4281 12.877
R54280 vp_n.n1078 vp_n.n1077 12.877
R54281 vp_n.n2639 vp_n.n2638 12.877
R54282 vp_n.n4292 vp_n.n4291 12.877
R54283 vp_n.n1088 vp_n.n1087 12.877
R54284 vp_n.n2649 vp_n.n2648 12.877
R54285 vp_n.n4302 vp_n.n4301 12.877
R54286 vp_n.n1098 vp_n.n1097 12.877
R54287 vp_n.n2659 vp_n.n2658 12.877
R54288 vp_n.n4312 vp_n.n4311 12.877
R54289 vp_n.n1108 vp_n.n1107 12.877
R54290 vp_n.n2669 vp_n.n2668 12.877
R54291 vp_n.n4322 vp_n.n4321 12.877
R54292 vp_n.n1118 vp_n.n1117 12.877
R54293 vp_n.n2679 vp_n.n2678 12.877
R54294 vp_n.n4332 vp_n.n4331 12.877
R54295 vp_n.n1128 vp_n.n1127 12.877
R54296 vp_n.n2689 vp_n.n2688 12.877
R54297 vp_n.n4342 vp_n.n4341 12.877
R54298 vp_n.n1138 vp_n.n1137 12.877
R54299 vp_n.n2699 vp_n.n2698 12.877
R54300 vp_n.n4352 vp_n.n4351 12.877
R54301 vp_n.n1148 vp_n.n1147 12.877
R54302 vp_n.n2709 vp_n.n2708 12.877
R54303 vp_n.n4362 vp_n.n4361 12.877
R54304 vp_n.n1158 vp_n.n1157 12.877
R54305 vp_n.n2719 vp_n.n2718 12.877
R54306 vp_n.n4372 vp_n.n4371 12.877
R54307 vp_n.n1168 vp_n.n1167 12.877
R54308 vp_n.n2729 vp_n.n2728 12.877
R54309 vp_n.n4382 vp_n.n4381 12.877
R54310 vp_n.n1178 vp_n.n1177 12.877
R54311 vp_n.n2739 vp_n.n2738 12.877
R54312 vp_n.n4392 vp_n.n4391 12.877
R54313 vp_n.n1188 vp_n.n1187 12.877
R54314 vp_n.n2749 vp_n.n2748 12.877
R54315 vp_n.n4402 vp_n.n4401 12.877
R54316 vp_n.n1198 vp_n.n1197 12.877
R54317 vp_n.n2759 vp_n.n2758 12.877
R54318 vp_n.n4412 vp_n.n4411 12.877
R54319 vp_n.n1208 vp_n.n1207 12.877
R54320 vp_n.n2769 vp_n.n2768 12.877
R54321 vp_n.n4422 vp_n.n4421 12.877
R54322 vp_n.n1218 vp_n.n1217 12.877
R54323 vp_n.n2779 vp_n.n2778 12.877
R54324 vp_n.n4432 vp_n.n4431 12.877
R54325 vp_n.n1228 vp_n.n1227 12.877
R54326 vp_n.n2789 vp_n.n2788 12.877
R54327 vp_n.n4442 vp_n.n4441 12.877
R54328 vp_n.n1238 vp_n.n1237 12.877
R54329 vp_n.n2799 vp_n.n2798 12.877
R54330 vp_n.n4452 vp_n.n4451 12.877
R54331 vp_n.n1248 vp_n.n1247 12.877
R54332 vp_n.n2809 vp_n.n2808 12.877
R54333 vp_n.n4462 vp_n.n4461 12.877
R54334 vp_n.n1258 vp_n.n1257 12.877
R54335 vp_n.n2819 vp_n.n2818 12.877
R54336 vp_n.n4472 vp_n.n4471 12.877
R54337 vp_n.n1268 vp_n.n1267 12.877
R54338 vp_n.n2829 vp_n.n2828 12.877
R54339 vp_n.n4482 vp_n.n4481 12.877
R54340 vp_n.n1278 vp_n.n1277 12.877
R54341 vp_n.n2839 vp_n.n2838 12.877
R54342 vp_n.n4492 vp_n.n4491 12.877
R54343 vp_n.n1288 vp_n.n1287 12.877
R54344 vp_n.n2849 vp_n.n2848 12.877
R54345 vp_n.n4502 vp_n.n4501 12.877
R54346 vp_n.n1298 vp_n.n1297 12.877
R54347 vp_n.n2859 vp_n.n2858 12.877
R54348 vp_n.n4512 vp_n.n4511 12.877
R54349 vp_n.n1308 vp_n.n1307 12.877
R54350 vp_n.n2869 vp_n.n2868 12.877
R54351 vp_n.n4522 vp_n.n4521 12.877
R54352 vp_n.n1318 vp_n.n1317 12.877
R54353 vp_n.n2879 vp_n.n2878 12.877
R54354 vp_n.n4532 vp_n.n4531 12.877
R54355 vp_n.n1328 vp_n.n1327 12.877
R54356 vp_n.n2889 vp_n.n2888 12.877
R54357 vp_n.n4542 vp_n.n4541 12.877
R54358 vp_n.n1338 vp_n.n1337 12.877
R54359 vp_n.n2899 vp_n.n2898 12.877
R54360 vp_n.n4552 vp_n.n4551 12.877
R54361 vp_n.n1348 vp_n.n1347 12.877
R54362 vp_n.n2909 vp_n.n2908 12.877
R54363 vp_n.n4562 vp_n.n4561 12.877
R54364 vp_n.n1358 vp_n.n1357 12.877
R54365 vp_n.n2919 vp_n.n2918 12.877
R54366 vp_n.n4572 vp_n.n4571 12.877
R54367 vp_n.n1368 vp_n.n1367 12.877
R54368 vp_n.n2929 vp_n.n2928 12.877
R54369 vp_n.n4582 vp_n.n4581 12.877
R54370 vp_n.n1378 vp_n.n1377 12.877
R54371 vp_n.n2939 vp_n.n2938 12.877
R54372 vp_n.n4592 vp_n.n4591 12.877
R54373 vp_n.n1388 vp_n.n1387 12.877
R54374 vp_n.n2949 vp_n.n2948 12.877
R54375 vp_n.n4602 vp_n.n4601 12.877
R54376 vp_n.n1398 vp_n.n1397 12.877
R54377 vp_n.n2959 vp_n.n2958 12.877
R54378 vp_n.n4612 vp_n.n4611 12.877
R54379 vp_n.n1408 vp_n.n1407 12.877
R54380 vp_n.n2969 vp_n.n2968 12.877
R54381 vp_n.n4622 vp_n.n4621 12.877
R54382 vp_n.n1418 vp_n.n1417 12.877
R54383 vp_n.n2979 vp_n.n2978 12.877
R54384 vp_n.n4632 vp_n.n4631 12.877
R54385 vp_n.n1428 vp_n.n1427 12.877
R54386 vp_n.n2989 vp_n.n2988 12.877
R54387 vp_n.n4642 vp_n.n4641 12.877
R54388 vp_n.n1438 vp_n.n1437 12.877
R54389 vp_n.n2999 vp_n.n2998 12.877
R54390 vp_n.n4652 vp_n.n4651 12.877
R54391 vp_n.n1448 vp_n.n1447 12.877
R54392 vp_n.n3009 vp_n.n3008 12.877
R54393 vp_n.n4662 vp_n.n4661 12.877
R54394 vp_n.n1458 vp_n.n1457 12.877
R54395 vp_n.n3019 vp_n.n3018 12.877
R54396 vp_n.n4672 vp_n.n4671 12.877
R54397 vp_n.n1468 vp_n.n1467 12.877
R54398 vp_n.n3029 vp_n.n3028 12.877
R54399 vp_n.n4682 vp_n.n4681 12.877
R54400 vp_n.n1478 vp_n.n1477 12.877
R54401 vp_n.n3039 vp_n.n3038 12.877
R54402 vp_n.n4692 vp_n.n4691 12.877
R54403 vp_n.n1488 vp_n.n1487 12.877
R54404 vp_n.n1498 vp_n.n1497 12.877
R54405 vp_n.n4702 vp_n.n4701 12.877
R54406 vp_n.n3049 vp_n.n3048 12.877
R54407 vp_n.n1569 vp_n.n1568 12.877
R54408 vp_n.n3222 vp_n.n3221 12.877
R54409 vp_n.n3212 vp_n.n3211 12.877
R54410 vp_n.n1559 vp_n.n1555 12.538
R54411 vp_n.n8 vp_n.n4 12.538
R54412 vp_n.n18 vp_n.n14 12.538
R54413 vp_n.n1579 vp_n.n1575 12.538
R54414 vp_n.n3232 vp_n.n3228 12.538
R54415 vp_n.n28 vp_n.n24 12.538
R54416 vp_n.n1589 vp_n.n1585 12.538
R54417 vp_n.n3242 vp_n.n3238 12.538
R54418 vp_n.n38 vp_n.n34 12.538
R54419 vp_n.n1599 vp_n.n1595 12.538
R54420 vp_n.n3252 vp_n.n3248 12.538
R54421 vp_n.n48 vp_n.n44 12.538
R54422 vp_n.n1609 vp_n.n1605 12.538
R54423 vp_n.n3262 vp_n.n3258 12.538
R54424 vp_n.n58 vp_n.n54 12.538
R54425 vp_n.n1619 vp_n.n1615 12.538
R54426 vp_n.n3272 vp_n.n3268 12.538
R54427 vp_n.n68 vp_n.n64 12.538
R54428 vp_n.n1629 vp_n.n1625 12.538
R54429 vp_n.n3282 vp_n.n3278 12.538
R54430 vp_n.n78 vp_n.n74 12.538
R54431 vp_n.n1639 vp_n.n1635 12.538
R54432 vp_n.n3292 vp_n.n3288 12.538
R54433 vp_n.n88 vp_n.n84 12.538
R54434 vp_n.n1649 vp_n.n1645 12.538
R54435 vp_n.n3302 vp_n.n3298 12.538
R54436 vp_n.n98 vp_n.n94 12.538
R54437 vp_n.n1659 vp_n.n1655 12.538
R54438 vp_n.n3312 vp_n.n3308 12.538
R54439 vp_n.n108 vp_n.n104 12.538
R54440 vp_n.n1669 vp_n.n1665 12.538
R54441 vp_n.n3322 vp_n.n3318 12.538
R54442 vp_n.n118 vp_n.n114 12.538
R54443 vp_n.n1679 vp_n.n1675 12.538
R54444 vp_n.n3332 vp_n.n3328 12.538
R54445 vp_n.n128 vp_n.n124 12.538
R54446 vp_n.n1689 vp_n.n1685 12.538
R54447 vp_n.n3342 vp_n.n3338 12.538
R54448 vp_n.n138 vp_n.n134 12.538
R54449 vp_n.n1699 vp_n.n1695 12.538
R54450 vp_n.n3352 vp_n.n3348 12.538
R54451 vp_n.n148 vp_n.n144 12.538
R54452 vp_n.n1709 vp_n.n1705 12.538
R54453 vp_n.n3362 vp_n.n3358 12.538
R54454 vp_n.n158 vp_n.n154 12.538
R54455 vp_n.n1719 vp_n.n1715 12.538
R54456 vp_n.n3372 vp_n.n3368 12.538
R54457 vp_n.n168 vp_n.n164 12.538
R54458 vp_n.n1729 vp_n.n1725 12.538
R54459 vp_n.n3382 vp_n.n3378 12.538
R54460 vp_n.n178 vp_n.n174 12.538
R54461 vp_n.n1739 vp_n.n1735 12.538
R54462 vp_n.n3392 vp_n.n3388 12.538
R54463 vp_n.n188 vp_n.n184 12.538
R54464 vp_n.n1749 vp_n.n1745 12.538
R54465 vp_n.n3402 vp_n.n3398 12.538
R54466 vp_n.n198 vp_n.n194 12.538
R54467 vp_n.n1759 vp_n.n1755 12.538
R54468 vp_n.n3412 vp_n.n3408 12.538
R54469 vp_n.n208 vp_n.n204 12.538
R54470 vp_n.n1769 vp_n.n1765 12.538
R54471 vp_n.n3422 vp_n.n3418 12.538
R54472 vp_n.n218 vp_n.n214 12.538
R54473 vp_n.n1779 vp_n.n1775 12.538
R54474 vp_n.n3432 vp_n.n3428 12.538
R54475 vp_n.n228 vp_n.n224 12.538
R54476 vp_n.n1789 vp_n.n1785 12.538
R54477 vp_n.n3442 vp_n.n3438 12.538
R54478 vp_n.n238 vp_n.n234 12.538
R54479 vp_n.n1799 vp_n.n1795 12.538
R54480 vp_n.n3452 vp_n.n3448 12.538
R54481 vp_n.n248 vp_n.n244 12.538
R54482 vp_n.n1809 vp_n.n1805 12.538
R54483 vp_n.n3462 vp_n.n3458 12.538
R54484 vp_n.n258 vp_n.n254 12.538
R54485 vp_n.n1819 vp_n.n1815 12.538
R54486 vp_n.n3472 vp_n.n3468 12.538
R54487 vp_n.n268 vp_n.n264 12.538
R54488 vp_n.n1829 vp_n.n1825 12.538
R54489 vp_n.n3482 vp_n.n3478 12.538
R54490 vp_n.n278 vp_n.n274 12.538
R54491 vp_n.n1839 vp_n.n1835 12.538
R54492 vp_n.n3492 vp_n.n3488 12.538
R54493 vp_n.n288 vp_n.n284 12.538
R54494 vp_n.n1849 vp_n.n1845 12.538
R54495 vp_n.n3502 vp_n.n3498 12.538
R54496 vp_n.n298 vp_n.n294 12.538
R54497 vp_n.n1859 vp_n.n1855 12.538
R54498 vp_n.n3512 vp_n.n3508 12.538
R54499 vp_n.n308 vp_n.n304 12.538
R54500 vp_n.n1869 vp_n.n1865 12.538
R54501 vp_n.n3522 vp_n.n3518 12.538
R54502 vp_n.n318 vp_n.n314 12.538
R54503 vp_n.n1879 vp_n.n1875 12.538
R54504 vp_n.n3532 vp_n.n3528 12.538
R54505 vp_n.n328 vp_n.n324 12.538
R54506 vp_n.n1889 vp_n.n1885 12.538
R54507 vp_n.n3542 vp_n.n3538 12.538
R54508 vp_n.n338 vp_n.n334 12.538
R54509 vp_n.n1899 vp_n.n1895 12.538
R54510 vp_n.n3552 vp_n.n3548 12.538
R54511 vp_n.n348 vp_n.n344 12.538
R54512 vp_n.n1909 vp_n.n1905 12.538
R54513 vp_n.n3562 vp_n.n3558 12.538
R54514 vp_n.n358 vp_n.n354 12.538
R54515 vp_n.n1919 vp_n.n1915 12.538
R54516 vp_n.n3572 vp_n.n3568 12.538
R54517 vp_n.n368 vp_n.n364 12.538
R54518 vp_n.n1929 vp_n.n1925 12.538
R54519 vp_n.n3582 vp_n.n3578 12.538
R54520 vp_n.n378 vp_n.n374 12.538
R54521 vp_n.n1939 vp_n.n1935 12.538
R54522 vp_n.n3592 vp_n.n3588 12.538
R54523 vp_n.n388 vp_n.n384 12.538
R54524 vp_n.n1949 vp_n.n1945 12.538
R54525 vp_n.n3602 vp_n.n3598 12.538
R54526 vp_n.n398 vp_n.n394 12.538
R54527 vp_n.n1959 vp_n.n1955 12.538
R54528 vp_n.n3612 vp_n.n3608 12.538
R54529 vp_n.n408 vp_n.n404 12.538
R54530 vp_n.n1969 vp_n.n1965 12.538
R54531 vp_n.n3622 vp_n.n3618 12.538
R54532 vp_n.n418 vp_n.n414 12.538
R54533 vp_n.n1979 vp_n.n1975 12.538
R54534 vp_n.n3632 vp_n.n3628 12.538
R54535 vp_n.n428 vp_n.n424 12.538
R54536 vp_n.n1989 vp_n.n1985 12.538
R54537 vp_n.n3642 vp_n.n3638 12.538
R54538 vp_n.n438 vp_n.n434 12.538
R54539 vp_n.n1999 vp_n.n1995 12.538
R54540 vp_n.n3652 vp_n.n3648 12.538
R54541 vp_n.n448 vp_n.n444 12.538
R54542 vp_n.n2009 vp_n.n2005 12.538
R54543 vp_n.n3662 vp_n.n3658 12.538
R54544 vp_n.n458 vp_n.n454 12.538
R54545 vp_n.n2019 vp_n.n2015 12.538
R54546 vp_n.n3672 vp_n.n3668 12.538
R54547 vp_n.n468 vp_n.n464 12.538
R54548 vp_n.n2029 vp_n.n2025 12.538
R54549 vp_n.n3682 vp_n.n3678 12.538
R54550 vp_n.n478 vp_n.n474 12.538
R54551 vp_n.n2039 vp_n.n2035 12.538
R54552 vp_n.n3692 vp_n.n3688 12.538
R54553 vp_n.n488 vp_n.n484 12.538
R54554 vp_n.n2049 vp_n.n2045 12.538
R54555 vp_n.n3702 vp_n.n3698 12.538
R54556 vp_n.n498 vp_n.n494 12.538
R54557 vp_n.n2059 vp_n.n2055 12.538
R54558 vp_n.n3712 vp_n.n3708 12.538
R54559 vp_n.n508 vp_n.n504 12.538
R54560 vp_n.n2069 vp_n.n2065 12.538
R54561 vp_n.n3722 vp_n.n3718 12.538
R54562 vp_n.n518 vp_n.n514 12.538
R54563 vp_n.n2079 vp_n.n2075 12.538
R54564 vp_n.n3732 vp_n.n3728 12.538
R54565 vp_n.n528 vp_n.n524 12.538
R54566 vp_n.n2089 vp_n.n2085 12.538
R54567 vp_n.n3742 vp_n.n3738 12.538
R54568 vp_n.n538 vp_n.n534 12.538
R54569 vp_n.n2099 vp_n.n2095 12.538
R54570 vp_n.n3752 vp_n.n3748 12.538
R54571 vp_n.n548 vp_n.n544 12.538
R54572 vp_n.n2109 vp_n.n2105 12.538
R54573 vp_n.n3762 vp_n.n3758 12.538
R54574 vp_n.n558 vp_n.n554 12.538
R54575 vp_n.n2119 vp_n.n2115 12.538
R54576 vp_n.n3772 vp_n.n3768 12.538
R54577 vp_n.n568 vp_n.n564 12.538
R54578 vp_n.n2129 vp_n.n2125 12.538
R54579 vp_n.n3782 vp_n.n3778 12.538
R54580 vp_n.n578 vp_n.n574 12.538
R54581 vp_n.n2139 vp_n.n2135 12.538
R54582 vp_n.n3792 vp_n.n3788 12.538
R54583 vp_n.n588 vp_n.n584 12.538
R54584 vp_n.n2149 vp_n.n2145 12.538
R54585 vp_n.n3802 vp_n.n3798 12.538
R54586 vp_n.n598 vp_n.n594 12.538
R54587 vp_n.n2159 vp_n.n2155 12.538
R54588 vp_n.n3812 vp_n.n3808 12.538
R54589 vp_n.n608 vp_n.n604 12.538
R54590 vp_n.n2169 vp_n.n2165 12.538
R54591 vp_n.n3822 vp_n.n3818 12.538
R54592 vp_n.n618 vp_n.n614 12.538
R54593 vp_n.n2179 vp_n.n2175 12.538
R54594 vp_n.n3832 vp_n.n3828 12.538
R54595 vp_n.n628 vp_n.n624 12.538
R54596 vp_n.n2189 vp_n.n2185 12.538
R54597 vp_n.n3842 vp_n.n3838 12.538
R54598 vp_n.n638 vp_n.n634 12.538
R54599 vp_n.n2199 vp_n.n2195 12.538
R54600 vp_n.n3852 vp_n.n3848 12.538
R54601 vp_n.n648 vp_n.n644 12.538
R54602 vp_n.n2209 vp_n.n2205 12.538
R54603 vp_n.n3862 vp_n.n3858 12.538
R54604 vp_n.n658 vp_n.n654 12.538
R54605 vp_n.n2219 vp_n.n2215 12.538
R54606 vp_n.n3872 vp_n.n3868 12.538
R54607 vp_n.n668 vp_n.n664 12.538
R54608 vp_n.n2229 vp_n.n2225 12.538
R54609 vp_n.n3882 vp_n.n3878 12.538
R54610 vp_n.n678 vp_n.n674 12.538
R54611 vp_n.n2239 vp_n.n2235 12.538
R54612 vp_n.n3892 vp_n.n3888 12.538
R54613 vp_n.n688 vp_n.n684 12.538
R54614 vp_n.n2249 vp_n.n2245 12.538
R54615 vp_n.n3902 vp_n.n3898 12.538
R54616 vp_n.n698 vp_n.n694 12.538
R54617 vp_n.n2259 vp_n.n2255 12.538
R54618 vp_n.n3912 vp_n.n3908 12.538
R54619 vp_n.n708 vp_n.n704 12.538
R54620 vp_n.n2269 vp_n.n2265 12.538
R54621 vp_n.n3922 vp_n.n3918 12.538
R54622 vp_n.n718 vp_n.n714 12.538
R54623 vp_n.n2279 vp_n.n2275 12.538
R54624 vp_n.n3932 vp_n.n3928 12.538
R54625 vp_n.n728 vp_n.n724 12.538
R54626 vp_n.n2289 vp_n.n2285 12.538
R54627 vp_n.n3942 vp_n.n3938 12.538
R54628 vp_n.n738 vp_n.n734 12.538
R54629 vp_n.n2299 vp_n.n2295 12.538
R54630 vp_n.n3952 vp_n.n3948 12.538
R54631 vp_n.n748 vp_n.n744 12.538
R54632 vp_n.n2309 vp_n.n2305 12.538
R54633 vp_n.n3962 vp_n.n3958 12.538
R54634 vp_n.n758 vp_n.n754 12.538
R54635 vp_n.n2319 vp_n.n2315 12.538
R54636 vp_n.n3972 vp_n.n3968 12.538
R54637 vp_n.n768 vp_n.n764 12.538
R54638 vp_n.n2329 vp_n.n2325 12.538
R54639 vp_n.n3982 vp_n.n3978 12.538
R54640 vp_n.n778 vp_n.n774 12.538
R54641 vp_n.n2339 vp_n.n2335 12.538
R54642 vp_n.n3992 vp_n.n3988 12.538
R54643 vp_n.n788 vp_n.n784 12.538
R54644 vp_n.n2349 vp_n.n2345 12.538
R54645 vp_n.n4002 vp_n.n3998 12.538
R54646 vp_n.n798 vp_n.n794 12.538
R54647 vp_n.n2359 vp_n.n2355 12.538
R54648 vp_n.n4012 vp_n.n4008 12.538
R54649 vp_n.n808 vp_n.n804 12.538
R54650 vp_n.n2369 vp_n.n2365 12.538
R54651 vp_n.n4022 vp_n.n4018 12.538
R54652 vp_n.n818 vp_n.n814 12.538
R54653 vp_n.n2379 vp_n.n2375 12.538
R54654 vp_n.n4032 vp_n.n4028 12.538
R54655 vp_n.n828 vp_n.n824 12.538
R54656 vp_n.n2389 vp_n.n2385 12.538
R54657 vp_n.n4042 vp_n.n4038 12.538
R54658 vp_n.n838 vp_n.n834 12.538
R54659 vp_n.n2399 vp_n.n2395 12.538
R54660 vp_n.n4052 vp_n.n4048 12.538
R54661 vp_n.n848 vp_n.n844 12.538
R54662 vp_n.n2409 vp_n.n2405 12.538
R54663 vp_n.n4062 vp_n.n4058 12.538
R54664 vp_n.n858 vp_n.n854 12.538
R54665 vp_n.n2419 vp_n.n2415 12.538
R54666 vp_n.n4072 vp_n.n4068 12.538
R54667 vp_n.n868 vp_n.n864 12.538
R54668 vp_n.n2429 vp_n.n2425 12.538
R54669 vp_n.n4082 vp_n.n4078 12.538
R54670 vp_n.n878 vp_n.n874 12.538
R54671 vp_n.n2439 vp_n.n2435 12.538
R54672 vp_n.n4092 vp_n.n4088 12.538
R54673 vp_n.n888 vp_n.n884 12.538
R54674 vp_n.n2449 vp_n.n2445 12.538
R54675 vp_n.n4102 vp_n.n4098 12.538
R54676 vp_n.n898 vp_n.n894 12.538
R54677 vp_n.n2459 vp_n.n2455 12.538
R54678 vp_n.n4112 vp_n.n4108 12.538
R54679 vp_n.n908 vp_n.n904 12.538
R54680 vp_n.n2469 vp_n.n2465 12.538
R54681 vp_n.n4122 vp_n.n4118 12.538
R54682 vp_n.n918 vp_n.n914 12.538
R54683 vp_n.n2479 vp_n.n2475 12.538
R54684 vp_n.n4132 vp_n.n4128 12.538
R54685 vp_n.n928 vp_n.n924 12.538
R54686 vp_n.n2489 vp_n.n2485 12.538
R54687 vp_n.n4142 vp_n.n4138 12.538
R54688 vp_n.n938 vp_n.n934 12.538
R54689 vp_n.n2499 vp_n.n2495 12.538
R54690 vp_n.n4152 vp_n.n4148 12.538
R54691 vp_n.n948 vp_n.n944 12.538
R54692 vp_n.n2509 vp_n.n2505 12.538
R54693 vp_n.n4162 vp_n.n4158 12.538
R54694 vp_n.n958 vp_n.n954 12.538
R54695 vp_n.n2519 vp_n.n2515 12.538
R54696 vp_n.n4172 vp_n.n4168 12.538
R54697 vp_n.n968 vp_n.n964 12.538
R54698 vp_n.n2529 vp_n.n2525 12.538
R54699 vp_n.n4182 vp_n.n4178 12.538
R54700 vp_n.n978 vp_n.n974 12.538
R54701 vp_n.n2539 vp_n.n2535 12.538
R54702 vp_n.n4192 vp_n.n4188 12.538
R54703 vp_n.n988 vp_n.n984 12.538
R54704 vp_n.n2549 vp_n.n2545 12.538
R54705 vp_n.n4202 vp_n.n4198 12.538
R54706 vp_n.n998 vp_n.n994 12.538
R54707 vp_n.n2559 vp_n.n2555 12.538
R54708 vp_n.n4212 vp_n.n4208 12.538
R54709 vp_n.n1008 vp_n.n1004 12.538
R54710 vp_n.n2569 vp_n.n2565 12.538
R54711 vp_n.n4222 vp_n.n4218 12.538
R54712 vp_n.n1018 vp_n.n1014 12.538
R54713 vp_n.n2579 vp_n.n2575 12.538
R54714 vp_n.n4232 vp_n.n4228 12.538
R54715 vp_n.n1028 vp_n.n1024 12.538
R54716 vp_n.n2589 vp_n.n2585 12.538
R54717 vp_n.n4242 vp_n.n4238 12.538
R54718 vp_n.n1038 vp_n.n1034 12.538
R54719 vp_n.n2599 vp_n.n2595 12.538
R54720 vp_n.n4252 vp_n.n4248 12.538
R54721 vp_n.n1048 vp_n.n1044 12.538
R54722 vp_n.n2609 vp_n.n2605 12.538
R54723 vp_n.n4262 vp_n.n4258 12.538
R54724 vp_n.n1058 vp_n.n1054 12.538
R54725 vp_n.n2619 vp_n.n2615 12.538
R54726 vp_n.n4272 vp_n.n4268 12.538
R54727 vp_n.n1068 vp_n.n1064 12.538
R54728 vp_n.n2629 vp_n.n2625 12.538
R54729 vp_n.n4282 vp_n.n4278 12.538
R54730 vp_n.n1078 vp_n.n1074 12.538
R54731 vp_n.n2639 vp_n.n2635 12.538
R54732 vp_n.n4292 vp_n.n4288 12.538
R54733 vp_n.n1088 vp_n.n1084 12.538
R54734 vp_n.n2649 vp_n.n2645 12.538
R54735 vp_n.n4302 vp_n.n4298 12.538
R54736 vp_n.n1098 vp_n.n1094 12.538
R54737 vp_n.n2659 vp_n.n2655 12.538
R54738 vp_n.n4312 vp_n.n4308 12.538
R54739 vp_n.n1108 vp_n.n1104 12.538
R54740 vp_n.n2669 vp_n.n2665 12.538
R54741 vp_n.n4322 vp_n.n4318 12.538
R54742 vp_n.n1118 vp_n.n1114 12.538
R54743 vp_n.n2679 vp_n.n2675 12.538
R54744 vp_n.n4332 vp_n.n4328 12.538
R54745 vp_n.n1128 vp_n.n1124 12.538
R54746 vp_n.n2689 vp_n.n2685 12.538
R54747 vp_n.n4342 vp_n.n4338 12.538
R54748 vp_n.n1138 vp_n.n1134 12.538
R54749 vp_n.n2699 vp_n.n2695 12.538
R54750 vp_n.n4352 vp_n.n4348 12.538
R54751 vp_n.n1148 vp_n.n1144 12.538
R54752 vp_n.n2709 vp_n.n2705 12.538
R54753 vp_n.n4362 vp_n.n4358 12.538
R54754 vp_n.n1158 vp_n.n1154 12.538
R54755 vp_n.n2719 vp_n.n2715 12.538
R54756 vp_n.n4372 vp_n.n4368 12.538
R54757 vp_n.n1168 vp_n.n1164 12.538
R54758 vp_n.n2729 vp_n.n2725 12.538
R54759 vp_n.n4382 vp_n.n4378 12.538
R54760 vp_n.n1178 vp_n.n1174 12.538
R54761 vp_n.n2739 vp_n.n2735 12.538
R54762 vp_n.n4392 vp_n.n4388 12.538
R54763 vp_n.n1188 vp_n.n1184 12.538
R54764 vp_n.n2749 vp_n.n2745 12.538
R54765 vp_n.n4402 vp_n.n4398 12.538
R54766 vp_n.n1198 vp_n.n1194 12.538
R54767 vp_n.n2759 vp_n.n2755 12.538
R54768 vp_n.n4412 vp_n.n4408 12.538
R54769 vp_n.n1208 vp_n.n1204 12.538
R54770 vp_n.n2769 vp_n.n2765 12.538
R54771 vp_n.n4422 vp_n.n4418 12.538
R54772 vp_n.n1218 vp_n.n1214 12.538
R54773 vp_n.n2779 vp_n.n2775 12.538
R54774 vp_n.n4432 vp_n.n4428 12.538
R54775 vp_n.n1228 vp_n.n1224 12.538
R54776 vp_n.n2789 vp_n.n2785 12.538
R54777 vp_n.n4442 vp_n.n4438 12.538
R54778 vp_n.n1238 vp_n.n1234 12.538
R54779 vp_n.n2799 vp_n.n2795 12.538
R54780 vp_n.n4452 vp_n.n4448 12.538
R54781 vp_n.n1248 vp_n.n1244 12.538
R54782 vp_n.n2809 vp_n.n2805 12.538
R54783 vp_n.n4462 vp_n.n4458 12.538
R54784 vp_n.n1258 vp_n.n1254 12.538
R54785 vp_n.n2819 vp_n.n2815 12.538
R54786 vp_n.n4472 vp_n.n4468 12.538
R54787 vp_n.n1268 vp_n.n1264 12.538
R54788 vp_n.n2829 vp_n.n2825 12.538
R54789 vp_n.n4482 vp_n.n4478 12.538
R54790 vp_n.n1278 vp_n.n1274 12.538
R54791 vp_n.n2839 vp_n.n2835 12.538
R54792 vp_n.n4492 vp_n.n4488 12.538
R54793 vp_n.n1288 vp_n.n1284 12.538
R54794 vp_n.n2849 vp_n.n2845 12.538
R54795 vp_n.n4502 vp_n.n4498 12.538
R54796 vp_n.n1298 vp_n.n1294 12.538
R54797 vp_n.n2859 vp_n.n2855 12.538
R54798 vp_n.n4512 vp_n.n4508 12.538
R54799 vp_n.n1308 vp_n.n1304 12.538
R54800 vp_n.n2869 vp_n.n2865 12.538
R54801 vp_n.n4522 vp_n.n4518 12.538
R54802 vp_n.n1318 vp_n.n1314 12.538
R54803 vp_n.n2879 vp_n.n2875 12.538
R54804 vp_n.n4532 vp_n.n4528 12.538
R54805 vp_n.n1328 vp_n.n1324 12.538
R54806 vp_n.n2889 vp_n.n2885 12.538
R54807 vp_n.n4542 vp_n.n4538 12.538
R54808 vp_n.n1338 vp_n.n1334 12.538
R54809 vp_n.n2899 vp_n.n2895 12.538
R54810 vp_n.n4552 vp_n.n4548 12.538
R54811 vp_n.n1348 vp_n.n1344 12.538
R54812 vp_n.n2909 vp_n.n2905 12.538
R54813 vp_n.n4562 vp_n.n4558 12.538
R54814 vp_n.n1358 vp_n.n1354 12.538
R54815 vp_n.n2919 vp_n.n2915 12.538
R54816 vp_n.n4572 vp_n.n4568 12.538
R54817 vp_n.n1368 vp_n.n1364 12.538
R54818 vp_n.n2929 vp_n.n2925 12.538
R54819 vp_n.n4582 vp_n.n4578 12.538
R54820 vp_n.n1378 vp_n.n1374 12.538
R54821 vp_n.n2939 vp_n.n2935 12.538
R54822 vp_n.n4592 vp_n.n4588 12.538
R54823 vp_n.n1388 vp_n.n1384 12.538
R54824 vp_n.n2949 vp_n.n2945 12.538
R54825 vp_n.n4602 vp_n.n4598 12.538
R54826 vp_n.n1398 vp_n.n1394 12.538
R54827 vp_n.n2959 vp_n.n2955 12.538
R54828 vp_n.n4612 vp_n.n4608 12.538
R54829 vp_n.n1408 vp_n.n1404 12.538
R54830 vp_n.n2969 vp_n.n2965 12.538
R54831 vp_n.n4622 vp_n.n4618 12.538
R54832 vp_n.n1418 vp_n.n1414 12.538
R54833 vp_n.n2979 vp_n.n2975 12.538
R54834 vp_n.n4632 vp_n.n4628 12.538
R54835 vp_n.n1428 vp_n.n1424 12.538
R54836 vp_n.n2989 vp_n.n2985 12.538
R54837 vp_n.n4642 vp_n.n4638 12.538
R54838 vp_n.n1438 vp_n.n1434 12.538
R54839 vp_n.n2999 vp_n.n2995 12.538
R54840 vp_n.n4652 vp_n.n4648 12.538
R54841 vp_n.n1448 vp_n.n1444 12.538
R54842 vp_n.n3009 vp_n.n3005 12.538
R54843 vp_n.n4662 vp_n.n4658 12.538
R54844 vp_n.n1458 vp_n.n1454 12.538
R54845 vp_n.n3019 vp_n.n3015 12.538
R54846 vp_n.n4672 vp_n.n4668 12.538
R54847 vp_n.n1468 vp_n.n1464 12.538
R54848 vp_n.n3029 vp_n.n3025 12.538
R54849 vp_n.n4682 vp_n.n4678 12.538
R54850 vp_n.n1478 vp_n.n1474 12.538
R54851 vp_n.n3039 vp_n.n3035 12.538
R54852 vp_n.n4692 vp_n.n4688 12.538
R54853 vp_n.n1488 vp_n.n1484 12.538
R54854 vp_n.n1498 vp_n.n1494 12.538
R54855 vp_n.n4702 vp_n.n4698 12.538
R54856 vp_n.n3049 vp_n.n3045 12.538
R54857 vp_n.n1569 vp_n.n1565 12.538
R54858 vp_n.n3222 vp_n.n3218 12.538
R54859 vp_n.n3212 vp_n.n3208 12.538
R54860 vp_n.n1555 vp_n.n1554 5.761
R54861 vp_n.n4 vp_n.n3 5.761
R54862 vp_n.n14 vp_n.n13 5.761
R54863 vp_n.n1575 vp_n.n1574 5.761
R54864 vp_n.n3228 vp_n.n3227 5.761
R54865 vp_n.n24 vp_n.n23 5.761
R54866 vp_n.n1585 vp_n.n1584 5.761
R54867 vp_n.n3238 vp_n.n3237 5.761
R54868 vp_n.n34 vp_n.n33 5.761
R54869 vp_n.n1595 vp_n.n1594 5.761
R54870 vp_n.n3248 vp_n.n3247 5.761
R54871 vp_n.n44 vp_n.n43 5.761
R54872 vp_n.n1605 vp_n.n1604 5.761
R54873 vp_n.n3258 vp_n.n3257 5.761
R54874 vp_n.n54 vp_n.n53 5.761
R54875 vp_n.n1615 vp_n.n1614 5.761
R54876 vp_n.n3268 vp_n.n3267 5.761
R54877 vp_n.n64 vp_n.n63 5.761
R54878 vp_n.n1625 vp_n.n1624 5.761
R54879 vp_n.n3278 vp_n.n3277 5.761
R54880 vp_n.n74 vp_n.n73 5.761
R54881 vp_n.n1635 vp_n.n1634 5.761
R54882 vp_n.n3288 vp_n.n3287 5.761
R54883 vp_n.n84 vp_n.n83 5.761
R54884 vp_n.n1645 vp_n.n1644 5.761
R54885 vp_n.n3298 vp_n.n3297 5.761
R54886 vp_n.n94 vp_n.n93 5.761
R54887 vp_n.n1655 vp_n.n1654 5.761
R54888 vp_n.n3308 vp_n.n3307 5.761
R54889 vp_n.n104 vp_n.n103 5.761
R54890 vp_n.n1665 vp_n.n1664 5.761
R54891 vp_n.n3318 vp_n.n3317 5.761
R54892 vp_n.n114 vp_n.n113 5.761
R54893 vp_n.n1675 vp_n.n1674 5.761
R54894 vp_n.n3328 vp_n.n3327 5.761
R54895 vp_n.n124 vp_n.n123 5.761
R54896 vp_n.n1685 vp_n.n1684 5.761
R54897 vp_n.n3338 vp_n.n3337 5.761
R54898 vp_n.n134 vp_n.n133 5.761
R54899 vp_n.n1695 vp_n.n1694 5.761
R54900 vp_n.n3348 vp_n.n3347 5.761
R54901 vp_n.n144 vp_n.n143 5.761
R54902 vp_n.n1705 vp_n.n1704 5.761
R54903 vp_n.n3358 vp_n.n3357 5.761
R54904 vp_n.n154 vp_n.n153 5.761
R54905 vp_n.n1715 vp_n.n1714 5.761
R54906 vp_n.n3368 vp_n.n3367 5.761
R54907 vp_n.n164 vp_n.n163 5.761
R54908 vp_n.n1725 vp_n.n1724 5.761
R54909 vp_n.n3378 vp_n.n3377 5.761
R54910 vp_n.n174 vp_n.n173 5.761
R54911 vp_n.n1735 vp_n.n1734 5.761
R54912 vp_n.n3388 vp_n.n3387 5.761
R54913 vp_n.n184 vp_n.n183 5.761
R54914 vp_n.n1745 vp_n.n1744 5.761
R54915 vp_n.n3398 vp_n.n3397 5.761
R54916 vp_n.n194 vp_n.n193 5.761
R54917 vp_n.n1755 vp_n.n1754 5.761
R54918 vp_n.n3408 vp_n.n3407 5.761
R54919 vp_n.n204 vp_n.n203 5.761
R54920 vp_n.n1765 vp_n.n1764 5.761
R54921 vp_n.n3418 vp_n.n3417 5.761
R54922 vp_n.n214 vp_n.n213 5.761
R54923 vp_n.n1775 vp_n.n1774 5.761
R54924 vp_n.n3428 vp_n.n3427 5.761
R54925 vp_n.n224 vp_n.n223 5.761
R54926 vp_n.n1785 vp_n.n1784 5.761
R54927 vp_n.n3438 vp_n.n3437 5.761
R54928 vp_n.n234 vp_n.n233 5.761
R54929 vp_n.n1795 vp_n.n1794 5.761
R54930 vp_n.n3448 vp_n.n3447 5.761
R54931 vp_n.n244 vp_n.n243 5.761
R54932 vp_n.n1805 vp_n.n1804 5.761
R54933 vp_n.n3458 vp_n.n3457 5.761
R54934 vp_n.n254 vp_n.n253 5.761
R54935 vp_n.n1815 vp_n.n1814 5.761
R54936 vp_n.n3468 vp_n.n3467 5.761
R54937 vp_n.n264 vp_n.n263 5.761
R54938 vp_n.n1825 vp_n.n1824 5.761
R54939 vp_n.n3478 vp_n.n3477 5.761
R54940 vp_n.n274 vp_n.n273 5.761
R54941 vp_n.n1835 vp_n.n1834 5.761
R54942 vp_n.n3488 vp_n.n3487 5.761
R54943 vp_n.n284 vp_n.n283 5.761
R54944 vp_n.n1845 vp_n.n1844 5.761
R54945 vp_n.n3498 vp_n.n3497 5.761
R54946 vp_n.n294 vp_n.n293 5.761
R54947 vp_n.n1855 vp_n.n1854 5.761
R54948 vp_n.n3508 vp_n.n3507 5.761
R54949 vp_n.n304 vp_n.n303 5.761
R54950 vp_n.n1865 vp_n.n1864 5.761
R54951 vp_n.n3518 vp_n.n3517 5.761
R54952 vp_n.n314 vp_n.n313 5.761
R54953 vp_n.n1875 vp_n.n1874 5.761
R54954 vp_n.n3528 vp_n.n3527 5.761
R54955 vp_n.n324 vp_n.n323 5.761
R54956 vp_n.n1885 vp_n.n1884 5.761
R54957 vp_n.n3538 vp_n.n3537 5.761
R54958 vp_n.n334 vp_n.n333 5.761
R54959 vp_n.n1895 vp_n.n1894 5.761
R54960 vp_n.n3548 vp_n.n3547 5.761
R54961 vp_n.n344 vp_n.n343 5.761
R54962 vp_n.n1905 vp_n.n1904 5.761
R54963 vp_n.n3558 vp_n.n3557 5.761
R54964 vp_n.n354 vp_n.n353 5.761
R54965 vp_n.n1915 vp_n.n1914 5.761
R54966 vp_n.n3568 vp_n.n3567 5.761
R54967 vp_n.n364 vp_n.n363 5.761
R54968 vp_n.n1925 vp_n.n1924 5.761
R54969 vp_n.n3578 vp_n.n3577 5.761
R54970 vp_n.n374 vp_n.n373 5.761
R54971 vp_n.n1935 vp_n.n1934 5.761
R54972 vp_n.n3588 vp_n.n3587 5.761
R54973 vp_n.n384 vp_n.n383 5.761
R54974 vp_n.n1945 vp_n.n1944 5.761
R54975 vp_n.n3598 vp_n.n3597 5.761
R54976 vp_n.n394 vp_n.n393 5.761
R54977 vp_n.n1955 vp_n.n1954 5.761
R54978 vp_n.n3608 vp_n.n3607 5.761
R54979 vp_n.n404 vp_n.n403 5.761
R54980 vp_n.n1965 vp_n.n1964 5.761
R54981 vp_n.n3618 vp_n.n3617 5.761
R54982 vp_n.n414 vp_n.n413 5.761
R54983 vp_n.n1975 vp_n.n1974 5.761
R54984 vp_n.n3628 vp_n.n3627 5.761
R54985 vp_n.n424 vp_n.n423 5.761
R54986 vp_n.n1985 vp_n.n1984 5.761
R54987 vp_n.n3638 vp_n.n3637 5.761
R54988 vp_n.n434 vp_n.n433 5.761
R54989 vp_n.n1995 vp_n.n1994 5.761
R54990 vp_n.n3648 vp_n.n3647 5.761
R54991 vp_n.n444 vp_n.n443 5.761
R54992 vp_n.n2005 vp_n.n2004 5.761
R54993 vp_n.n3658 vp_n.n3657 5.761
R54994 vp_n.n454 vp_n.n453 5.761
R54995 vp_n.n2015 vp_n.n2014 5.761
R54996 vp_n.n3668 vp_n.n3667 5.761
R54997 vp_n.n464 vp_n.n463 5.761
R54998 vp_n.n2025 vp_n.n2024 5.761
R54999 vp_n.n3678 vp_n.n3677 5.761
R55000 vp_n.n474 vp_n.n473 5.761
R55001 vp_n.n2035 vp_n.n2034 5.761
R55002 vp_n.n3688 vp_n.n3687 5.761
R55003 vp_n.n484 vp_n.n483 5.761
R55004 vp_n.n2045 vp_n.n2044 5.761
R55005 vp_n.n3698 vp_n.n3697 5.761
R55006 vp_n.n494 vp_n.n493 5.761
R55007 vp_n.n2055 vp_n.n2054 5.761
R55008 vp_n.n3708 vp_n.n3707 5.761
R55009 vp_n.n504 vp_n.n503 5.761
R55010 vp_n.n2065 vp_n.n2064 5.761
R55011 vp_n.n3718 vp_n.n3717 5.761
R55012 vp_n.n514 vp_n.n513 5.761
R55013 vp_n.n2075 vp_n.n2074 5.761
R55014 vp_n.n3728 vp_n.n3727 5.761
R55015 vp_n.n524 vp_n.n523 5.761
R55016 vp_n.n2085 vp_n.n2084 5.761
R55017 vp_n.n3738 vp_n.n3737 5.761
R55018 vp_n.n534 vp_n.n533 5.761
R55019 vp_n.n2095 vp_n.n2094 5.761
R55020 vp_n.n3748 vp_n.n3747 5.761
R55021 vp_n.n544 vp_n.n543 5.761
R55022 vp_n.n2105 vp_n.n2104 5.761
R55023 vp_n.n3758 vp_n.n3757 5.761
R55024 vp_n.n554 vp_n.n553 5.761
R55025 vp_n.n2115 vp_n.n2114 5.761
R55026 vp_n.n3768 vp_n.n3767 5.761
R55027 vp_n.n564 vp_n.n563 5.761
R55028 vp_n.n2125 vp_n.n2124 5.761
R55029 vp_n.n3778 vp_n.n3777 5.761
R55030 vp_n.n574 vp_n.n573 5.761
R55031 vp_n.n2135 vp_n.n2134 5.761
R55032 vp_n.n3788 vp_n.n3787 5.761
R55033 vp_n.n584 vp_n.n583 5.761
R55034 vp_n.n2145 vp_n.n2144 5.761
R55035 vp_n.n3798 vp_n.n3797 5.761
R55036 vp_n.n594 vp_n.n593 5.761
R55037 vp_n.n2155 vp_n.n2154 5.761
R55038 vp_n.n3808 vp_n.n3807 5.761
R55039 vp_n.n604 vp_n.n603 5.761
R55040 vp_n.n2165 vp_n.n2164 5.761
R55041 vp_n.n3818 vp_n.n3817 5.761
R55042 vp_n.n614 vp_n.n613 5.761
R55043 vp_n.n2175 vp_n.n2174 5.761
R55044 vp_n.n3828 vp_n.n3827 5.761
R55045 vp_n.n624 vp_n.n623 5.761
R55046 vp_n.n2185 vp_n.n2184 5.761
R55047 vp_n.n3838 vp_n.n3837 5.761
R55048 vp_n.n634 vp_n.n633 5.761
R55049 vp_n.n2195 vp_n.n2194 5.761
R55050 vp_n.n3848 vp_n.n3847 5.761
R55051 vp_n.n644 vp_n.n643 5.761
R55052 vp_n.n2205 vp_n.n2204 5.761
R55053 vp_n.n3858 vp_n.n3857 5.761
R55054 vp_n.n654 vp_n.n653 5.761
R55055 vp_n.n2215 vp_n.n2214 5.761
R55056 vp_n.n3868 vp_n.n3867 5.761
R55057 vp_n.n664 vp_n.n663 5.761
R55058 vp_n.n2225 vp_n.n2224 5.761
R55059 vp_n.n3878 vp_n.n3877 5.761
R55060 vp_n.n674 vp_n.n673 5.761
R55061 vp_n.n2235 vp_n.n2234 5.761
R55062 vp_n.n3888 vp_n.n3887 5.761
R55063 vp_n.n684 vp_n.n683 5.761
R55064 vp_n.n2245 vp_n.n2244 5.761
R55065 vp_n.n3898 vp_n.n3897 5.761
R55066 vp_n.n694 vp_n.n693 5.761
R55067 vp_n.n2255 vp_n.n2254 5.761
R55068 vp_n.n3908 vp_n.n3907 5.761
R55069 vp_n.n704 vp_n.n703 5.761
R55070 vp_n.n2265 vp_n.n2264 5.761
R55071 vp_n.n3918 vp_n.n3917 5.761
R55072 vp_n.n714 vp_n.n713 5.761
R55073 vp_n.n2275 vp_n.n2274 5.761
R55074 vp_n.n3928 vp_n.n3927 5.761
R55075 vp_n.n724 vp_n.n723 5.761
R55076 vp_n.n2285 vp_n.n2284 5.761
R55077 vp_n.n3938 vp_n.n3937 5.761
R55078 vp_n.n734 vp_n.n733 5.761
R55079 vp_n.n2295 vp_n.n2294 5.761
R55080 vp_n.n3948 vp_n.n3947 5.761
R55081 vp_n.n744 vp_n.n743 5.761
R55082 vp_n.n2305 vp_n.n2304 5.761
R55083 vp_n.n3958 vp_n.n3957 5.761
R55084 vp_n.n754 vp_n.n753 5.761
R55085 vp_n.n2315 vp_n.n2314 5.761
R55086 vp_n.n3968 vp_n.n3967 5.761
R55087 vp_n.n764 vp_n.n763 5.761
R55088 vp_n.n2325 vp_n.n2324 5.761
R55089 vp_n.n3978 vp_n.n3977 5.761
R55090 vp_n.n774 vp_n.n773 5.761
R55091 vp_n.n2335 vp_n.n2334 5.761
R55092 vp_n.n3988 vp_n.n3987 5.761
R55093 vp_n.n784 vp_n.n783 5.761
R55094 vp_n.n2345 vp_n.n2344 5.761
R55095 vp_n.n3998 vp_n.n3997 5.761
R55096 vp_n.n794 vp_n.n793 5.761
R55097 vp_n.n2355 vp_n.n2354 5.761
R55098 vp_n.n4008 vp_n.n4007 5.761
R55099 vp_n.n804 vp_n.n803 5.761
R55100 vp_n.n2365 vp_n.n2364 5.761
R55101 vp_n.n4018 vp_n.n4017 5.761
R55102 vp_n.n814 vp_n.n813 5.761
R55103 vp_n.n2375 vp_n.n2374 5.761
R55104 vp_n.n4028 vp_n.n4027 5.761
R55105 vp_n.n824 vp_n.n823 5.761
R55106 vp_n.n2385 vp_n.n2384 5.761
R55107 vp_n.n4038 vp_n.n4037 5.761
R55108 vp_n.n834 vp_n.n833 5.761
R55109 vp_n.n2395 vp_n.n2394 5.761
R55110 vp_n.n4048 vp_n.n4047 5.761
R55111 vp_n.n844 vp_n.n843 5.761
R55112 vp_n.n2405 vp_n.n2404 5.761
R55113 vp_n.n4058 vp_n.n4057 5.761
R55114 vp_n.n854 vp_n.n853 5.761
R55115 vp_n.n2415 vp_n.n2414 5.761
R55116 vp_n.n4068 vp_n.n4067 5.761
R55117 vp_n.n864 vp_n.n863 5.761
R55118 vp_n.n2425 vp_n.n2424 5.761
R55119 vp_n.n4078 vp_n.n4077 5.761
R55120 vp_n.n874 vp_n.n873 5.761
R55121 vp_n.n2435 vp_n.n2434 5.761
R55122 vp_n.n4088 vp_n.n4087 5.761
R55123 vp_n.n884 vp_n.n883 5.761
R55124 vp_n.n2445 vp_n.n2444 5.761
R55125 vp_n.n4098 vp_n.n4097 5.761
R55126 vp_n.n894 vp_n.n893 5.761
R55127 vp_n.n2455 vp_n.n2454 5.761
R55128 vp_n.n4108 vp_n.n4107 5.761
R55129 vp_n.n904 vp_n.n903 5.761
R55130 vp_n.n2465 vp_n.n2464 5.761
R55131 vp_n.n4118 vp_n.n4117 5.761
R55132 vp_n.n914 vp_n.n913 5.761
R55133 vp_n.n2475 vp_n.n2474 5.761
R55134 vp_n.n4128 vp_n.n4127 5.761
R55135 vp_n.n924 vp_n.n923 5.761
R55136 vp_n.n2485 vp_n.n2484 5.761
R55137 vp_n.n4138 vp_n.n4137 5.761
R55138 vp_n.n934 vp_n.n933 5.761
R55139 vp_n.n2495 vp_n.n2494 5.761
R55140 vp_n.n4148 vp_n.n4147 5.761
R55141 vp_n.n944 vp_n.n943 5.761
R55142 vp_n.n2505 vp_n.n2504 5.761
R55143 vp_n.n4158 vp_n.n4157 5.761
R55144 vp_n.n954 vp_n.n953 5.761
R55145 vp_n.n2515 vp_n.n2514 5.761
R55146 vp_n.n4168 vp_n.n4167 5.761
R55147 vp_n.n964 vp_n.n963 5.761
R55148 vp_n.n2525 vp_n.n2524 5.761
R55149 vp_n.n4178 vp_n.n4177 5.761
R55150 vp_n.n974 vp_n.n973 5.761
R55151 vp_n.n2535 vp_n.n2534 5.761
R55152 vp_n.n4188 vp_n.n4187 5.761
R55153 vp_n.n984 vp_n.n983 5.761
R55154 vp_n.n2545 vp_n.n2544 5.761
R55155 vp_n.n4198 vp_n.n4197 5.761
R55156 vp_n.n994 vp_n.n993 5.761
R55157 vp_n.n2555 vp_n.n2554 5.761
R55158 vp_n.n4208 vp_n.n4207 5.761
R55159 vp_n.n1004 vp_n.n1003 5.761
R55160 vp_n.n2565 vp_n.n2564 5.761
R55161 vp_n.n4218 vp_n.n4217 5.761
R55162 vp_n.n1014 vp_n.n1013 5.761
R55163 vp_n.n2575 vp_n.n2574 5.761
R55164 vp_n.n4228 vp_n.n4227 5.761
R55165 vp_n.n1024 vp_n.n1023 5.761
R55166 vp_n.n2585 vp_n.n2584 5.761
R55167 vp_n.n4238 vp_n.n4237 5.761
R55168 vp_n.n1034 vp_n.n1033 5.761
R55169 vp_n.n2595 vp_n.n2594 5.761
R55170 vp_n.n4248 vp_n.n4247 5.761
R55171 vp_n.n1044 vp_n.n1043 5.761
R55172 vp_n.n2605 vp_n.n2604 5.761
R55173 vp_n.n4258 vp_n.n4257 5.761
R55174 vp_n.n1054 vp_n.n1053 5.761
R55175 vp_n.n2615 vp_n.n2614 5.761
R55176 vp_n.n4268 vp_n.n4267 5.761
R55177 vp_n.n1064 vp_n.n1063 5.761
R55178 vp_n.n2625 vp_n.n2624 5.761
R55179 vp_n.n4278 vp_n.n4277 5.761
R55180 vp_n.n1074 vp_n.n1073 5.761
R55181 vp_n.n2635 vp_n.n2634 5.761
R55182 vp_n.n4288 vp_n.n4287 5.761
R55183 vp_n.n1084 vp_n.n1083 5.761
R55184 vp_n.n2645 vp_n.n2644 5.761
R55185 vp_n.n4298 vp_n.n4297 5.761
R55186 vp_n.n1094 vp_n.n1093 5.761
R55187 vp_n.n2655 vp_n.n2654 5.761
R55188 vp_n.n4308 vp_n.n4307 5.761
R55189 vp_n.n1104 vp_n.n1103 5.761
R55190 vp_n.n2665 vp_n.n2664 5.761
R55191 vp_n.n4318 vp_n.n4317 5.761
R55192 vp_n.n1114 vp_n.n1113 5.761
R55193 vp_n.n2675 vp_n.n2674 5.761
R55194 vp_n.n4328 vp_n.n4327 5.761
R55195 vp_n.n1124 vp_n.n1123 5.761
R55196 vp_n.n2685 vp_n.n2684 5.761
R55197 vp_n.n4338 vp_n.n4337 5.761
R55198 vp_n.n1134 vp_n.n1133 5.761
R55199 vp_n.n2695 vp_n.n2694 5.761
R55200 vp_n.n4348 vp_n.n4347 5.761
R55201 vp_n.n1144 vp_n.n1143 5.761
R55202 vp_n.n2705 vp_n.n2704 5.761
R55203 vp_n.n4358 vp_n.n4357 5.761
R55204 vp_n.n1154 vp_n.n1153 5.761
R55205 vp_n.n2715 vp_n.n2714 5.761
R55206 vp_n.n4368 vp_n.n4367 5.761
R55207 vp_n.n1164 vp_n.n1163 5.761
R55208 vp_n.n2725 vp_n.n2724 5.761
R55209 vp_n.n4378 vp_n.n4377 5.761
R55210 vp_n.n1174 vp_n.n1173 5.761
R55211 vp_n.n2735 vp_n.n2734 5.761
R55212 vp_n.n4388 vp_n.n4387 5.761
R55213 vp_n.n1184 vp_n.n1183 5.761
R55214 vp_n.n2745 vp_n.n2744 5.761
R55215 vp_n.n4398 vp_n.n4397 5.761
R55216 vp_n.n1194 vp_n.n1193 5.761
R55217 vp_n.n2755 vp_n.n2754 5.761
R55218 vp_n.n4408 vp_n.n4407 5.761
R55219 vp_n.n1204 vp_n.n1203 5.761
R55220 vp_n.n2765 vp_n.n2764 5.761
R55221 vp_n.n4418 vp_n.n4417 5.761
R55222 vp_n.n1214 vp_n.n1213 5.761
R55223 vp_n.n2775 vp_n.n2774 5.761
R55224 vp_n.n4428 vp_n.n4427 5.761
R55225 vp_n.n1224 vp_n.n1223 5.761
R55226 vp_n.n2785 vp_n.n2784 5.761
R55227 vp_n.n4438 vp_n.n4437 5.761
R55228 vp_n.n1234 vp_n.n1233 5.761
R55229 vp_n.n2795 vp_n.n2794 5.761
R55230 vp_n.n4448 vp_n.n4447 5.761
R55231 vp_n.n1244 vp_n.n1243 5.761
R55232 vp_n.n2805 vp_n.n2804 5.761
R55233 vp_n.n4458 vp_n.n4457 5.761
R55234 vp_n.n1254 vp_n.n1253 5.761
R55235 vp_n.n2815 vp_n.n2814 5.761
R55236 vp_n.n4468 vp_n.n4467 5.761
R55237 vp_n.n1264 vp_n.n1263 5.761
R55238 vp_n.n2825 vp_n.n2824 5.761
R55239 vp_n.n4478 vp_n.n4477 5.761
R55240 vp_n.n1274 vp_n.n1273 5.761
R55241 vp_n.n2835 vp_n.n2834 5.761
R55242 vp_n.n4488 vp_n.n4487 5.761
R55243 vp_n.n1284 vp_n.n1283 5.761
R55244 vp_n.n2845 vp_n.n2844 5.761
R55245 vp_n.n4498 vp_n.n4497 5.761
R55246 vp_n.n1294 vp_n.n1293 5.761
R55247 vp_n.n2855 vp_n.n2854 5.761
R55248 vp_n.n4508 vp_n.n4507 5.761
R55249 vp_n.n1304 vp_n.n1303 5.761
R55250 vp_n.n2865 vp_n.n2864 5.761
R55251 vp_n.n4518 vp_n.n4517 5.761
R55252 vp_n.n1314 vp_n.n1313 5.761
R55253 vp_n.n2875 vp_n.n2874 5.761
R55254 vp_n.n4528 vp_n.n4527 5.761
R55255 vp_n.n1324 vp_n.n1323 5.761
R55256 vp_n.n2885 vp_n.n2884 5.761
R55257 vp_n.n4538 vp_n.n4537 5.761
R55258 vp_n.n1334 vp_n.n1333 5.761
R55259 vp_n.n2895 vp_n.n2894 5.761
R55260 vp_n.n4548 vp_n.n4547 5.761
R55261 vp_n.n1344 vp_n.n1343 5.761
R55262 vp_n.n2905 vp_n.n2904 5.761
R55263 vp_n.n4558 vp_n.n4557 5.761
R55264 vp_n.n1354 vp_n.n1353 5.761
R55265 vp_n.n2915 vp_n.n2914 5.761
R55266 vp_n.n4568 vp_n.n4567 5.761
R55267 vp_n.n1364 vp_n.n1363 5.761
R55268 vp_n.n2925 vp_n.n2924 5.761
R55269 vp_n.n4578 vp_n.n4577 5.761
R55270 vp_n.n1374 vp_n.n1373 5.761
R55271 vp_n.n2935 vp_n.n2934 5.761
R55272 vp_n.n4588 vp_n.n4587 5.761
R55273 vp_n.n1384 vp_n.n1383 5.761
R55274 vp_n.n2945 vp_n.n2944 5.761
R55275 vp_n.n4598 vp_n.n4597 5.761
R55276 vp_n.n1394 vp_n.n1393 5.761
R55277 vp_n.n2955 vp_n.n2954 5.761
R55278 vp_n.n4608 vp_n.n4607 5.761
R55279 vp_n.n1404 vp_n.n1403 5.761
R55280 vp_n.n2965 vp_n.n2964 5.761
R55281 vp_n.n4618 vp_n.n4617 5.761
R55282 vp_n.n1414 vp_n.n1413 5.761
R55283 vp_n.n2975 vp_n.n2974 5.761
R55284 vp_n.n4628 vp_n.n4627 5.761
R55285 vp_n.n1424 vp_n.n1423 5.761
R55286 vp_n.n2985 vp_n.n2984 5.761
R55287 vp_n.n4638 vp_n.n4637 5.761
R55288 vp_n.n1434 vp_n.n1433 5.761
R55289 vp_n.n2995 vp_n.n2994 5.761
R55290 vp_n.n4648 vp_n.n4647 5.761
R55291 vp_n.n1444 vp_n.n1443 5.761
R55292 vp_n.n3005 vp_n.n3004 5.761
R55293 vp_n.n4658 vp_n.n4657 5.761
R55294 vp_n.n1454 vp_n.n1453 5.761
R55295 vp_n.n3015 vp_n.n3014 5.761
R55296 vp_n.n4668 vp_n.n4667 5.761
R55297 vp_n.n1464 vp_n.n1463 5.761
R55298 vp_n.n3025 vp_n.n3024 5.761
R55299 vp_n.n4678 vp_n.n4677 5.761
R55300 vp_n.n1474 vp_n.n1473 5.761
R55301 vp_n.n3035 vp_n.n3034 5.761
R55302 vp_n.n4688 vp_n.n4687 5.761
R55303 vp_n.n1484 vp_n.n1483 5.761
R55304 vp_n.n1494 vp_n.n1493 5.761
R55305 vp_n.n4698 vp_n.n4697 5.761
R55306 vp_n.n3045 vp_n.n3044 5.761
R55307 vp_n.n1565 vp_n.n1564 5.761
R55308 vp_n.n3218 vp_n.n3217 5.761
R55309 vp_n.n3208 vp_n.n3207 5.761
R55310 vp_n.n1558 vp_n.n1557 5.422
R55311 vp_n.n7 vp_n.n6 5.422
R55312 vp_n.n17 vp_n.n16 5.422
R55313 vp_n.n1578 vp_n.n1577 5.422
R55314 vp_n.n3231 vp_n.n3230 5.422
R55315 vp_n.n27 vp_n.n26 5.422
R55316 vp_n.n1588 vp_n.n1587 5.422
R55317 vp_n.n3241 vp_n.n3240 5.422
R55318 vp_n.n37 vp_n.n36 5.422
R55319 vp_n.n1598 vp_n.n1597 5.422
R55320 vp_n.n3251 vp_n.n3250 5.422
R55321 vp_n.n47 vp_n.n46 5.422
R55322 vp_n.n1608 vp_n.n1607 5.422
R55323 vp_n.n3261 vp_n.n3260 5.422
R55324 vp_n.n57 vp_n.n56 5.422
R55325 vp_n.n1618 vp_n.n1617 5.422
R55326 vp_n.n3271 vp_n.n3270 5.422
R55327 vp_n.n67 vp_n.n66 5.422
R55328 vp_n.n1628 vp_n.n1627 5.422
R55329 vp_n.n3281 vp_n.n3280 5.422
R55330 vp_n.n77 vp_n.n76 5.422
R55331 vp_n.n1638 vp_n.n1637 5.422
R55332 vp_n.n3291 vp_n.n3290 5.422
R55333 vp_n.n87 vp_n.n86 5.422
R55334 vp_n.n1648 vp_n.n1647 5.422
R55335 vp_n.n3301 vp_n.n3300 5.422
R55336 vp_n.n97 vp_n.n96 5.422
R55337 vp_n.n1658 vp_n.n1657 5.422
R55338 vp_n.n3311 vp_n.n3310 5.422
R55339 vp_n.n107 vp_n.n106 5.422
R55340 vp_n.n1668 vp_n.n1667 5.422
R55341 vp_n.n3321 vp_n.n3320 5.422
R55342 vp_n.n117 vp_n.n116 5.422
R55343 vp_n.n1678 vp_n.n1677 5.422
R55344 vp_n.n3331 vp_n.n3330 5.422
R55345 vp_n.n127 vp_n.n126 5.422
R55346 vp_n.n1688 vp_n.n1687 5.422
R55347 vp_n.n3341 vp_n.n3340 5.422
R55348 vp_n.n137 vp_n.n136 5.422
R55349 vp_n.n1698 vp_n.n1697 5.422
R55350 vp_n.n3351 vp_n.n3350 5.422
R55351 vp_n.n147 vp_n.n146 5.422
R55352 vp_n.n1708 vp_n.n1707 5.422
R55353 vp_n.n3361 vp_n.n3360 5.422
R55354 vp_n.n157 vp_n.n156 5.422
R55355 vp_n.n1718 vp_n.n1717 5.422
R55356 vp_n.n3371 vp_n.n3370 5.422
R55357 vp_n.n167 vp_n.n166 5.422
R55358 vp_n.n1728 vp_n.n1727 5.422
R55359 vp_n.n3381 vp_n.n3380 5.422
R55360 vp_n.n177 vp_n.n176 5.422
R55361 vp_n.n1738 vp_n.n1737 5.422
R55362 vp_n.n3391 vp_n.n3390 5.422
R55363 vp_n.n187 vp_n.n186 5.422
R55364 vp_n.n1748 vp_n.n1747 5.422
R55365 vp_n.n3401 vp_n.n3400 5.422
R55366 vp_n.n197 vp_n.n196 5.422
R55367 vp_n.n1758 vp_n.n1757 5.422
R55368 vp_n.n3411 vp_n.n3410 5.422
R55369 vp_n.n207 vp_n.n206 5.422
R55370 vp_n.n1768 vp_n.n1767 5.422
R55371 vp_n.n3421 vp_n.n3420 5.422
R55372 vp_n.n217 vp_n.n216 5.422
R55373 vp_n.n1778 vp_n.n1777 5.422
R55374 vp_n.n3431 vp_n.n3430 5.422
R55375 vp_n.n227 vp_n.n226 5.422
R55376 vp_n.n1788 vp_n.n1787 5.422
R55377 vp_n.n3441 vp_n.n3440 5.422
R55378 vp_n.n237 vp_n.n236 5.422
R55379 vp_n.n1798 vp_n.n1797 5.422
R55380 vp_n.n3451 vp_n.n3450 5.422
R55381 vp_n.n247 vp_n.n246 5.422
R55382 vp_n.n1808 vp_n.n1807 5.422
R55383 vp_n.n3461 vp_n.n3460 5.422
R55384 vp_n.n257 vp_n.n256 5.422
R55385 vp_n.n1818 vp_n.n1817 5.422
R55386 vp_n.n3471 vp_n.n3470 5.422
R55387 vp_n.n267 vp_n.n266 5.422
R55388 vp_n.n1828 vp_n.n1827 5.422
R55389 vp_n.n3481 vp_n.n3480 5.422
R55390 vp_n.n277 vp_n.n276 5.422
R55391 vp_n.n1838 vp_n.n1837 5.422
R55392 vp_n.n3491 vp_n.n3490 5.422
R55393 vp_n.n287 vp_n.n286 5.422
R55394 vp_n.n1848 vp_n.n1847 5.422
R55395 vp_n.n3501 vp_n.n3500 5.422
R55396 vp_n.n297 vp_n.n296 5.422
R55397 vp_n.n1858 vp_n.n1857 5.422
R55398 vp_n.n3511 vp_n.n3510 5.422
R55399 vp_n.n307 vp_n.n306 5.422
R55400 vp_n.n1868 vp_n.n1867 5.422
R55401 vp_n.n3521 vp_n.n3520 5.422
R55402 vp_n.n317 vp_n.n316 5.422
R55403 vp_n.n1878 vp_n.n1877 5.422
R55404 vp_n.n3531 vp_n.n3530 5.422
R55405 vp_n.n327 vp_n.n326 5.422
R55406 vp_n.n1888 vp_n.n1887 5.422
R55407 vp_n.n3541 vp_n.n3540 5.422
R55408 vp_n.n337 vp_n.n336 5.422
R55409 vp_n.n1898 vp_n.n1897 5.422
R55410 vp_n.n3551 vp_n.n3550 5.422
R55411 vp_n.n347 vp_n.n346 5.422
R55412 vp_n.n1908 vp_n.n1907 5.422
R55413 vp_n.n3561 vp_n.n3560 5.422
R55414 vp_n.n357 vp_n.n356 5.422
R55415 vp_n.n1918 vp_n.n1917 5.422
R55416 vp_n.n3571 vp_n.n3570 5.422
R55417 vp_n.n367 vp_n.n366 5.422
R55418 vp_n.n1928 vp_n.n1927 5.422
R55419 vp_n.n3581 vp_n.n3580 5.422
R55420 vp_n.n377 vp_n.n376 5.422
R55421 vp_n.n1938 vp_n.n1937 5.422
R55422 vp_n.n3591 vp_n.n3590 5.422
R55423 vp_n.n387 vp_n.n386 5.422
R55424 vp_n.n1948 vp_n.n1947 5.422
R55425 vp_n.n3601 vp_n.n3600 5.422
R55426 vp_n.n397 vp_n.n396 5.422
R55427 vp_n.n1958 vp_n.n1957 5.422
R55428 vp_n.n3611 vp_n.n3610 5.422
R55429 vp_n.n407 vp_n.n406 5.422
R55430 vp_n.n1968 vp_n.n1967 5.422
R55431 vp_n.n3621 vp_n.n3620 5.422
R55432 vp_n.n417 vp_n.n416 5.422
R55433 vp_n.n1978 vp_n.n1977 5.422
R55434 vp_n.n3631 vp_n.n3630 5.422
R55435 vp_n.n427 vp_n.n426 5.422
R55436 vp_n.n1988 vp_n.n1987 5.422
R55437 vp_n.n3641 vp_n.n3640 5.422
R55438 vp_n.n437 vp_n.n436 5.422
R55439 vp_n.n1998 vp_n.n1997 5.422
R55440 vp_n.n3651 vp_n.n3650 5.422
R55441 vp_n.n447 vp_n.n446 5.422
R55442 vp_n.n2008 vp_n.n2007 5.422
R55443 vp_n.n3661 vp_n.n3660 5.422
R55444 vp_n.n457 vp_n.n456 5.422
R55445 vp_n.n2018 vp_n.n2017 5.422
R55446 vp_n.n3671 vp_n.n3670 5.422
R55447 vp_n.n467 vp_n.n466 5.422
R55448 vp_n.n2028 vp_n.n2027 5.422
R55449 vp_n.n3681 vp_n.n3680 5.422
R55450 vp_n.n477 vp_n.n476 5.422
R55451 vp_n.n2038 vp_n.n2037 5.422
R55452 vp_n.n3691 vp_n.n3690 5.422
R55453 vp_n.n487 vp_n.n486 5.422
R55454 vp_n.n2048 vp_n.n2047 5.422
R55455 vp_n.n3701 vp_n.n3700 5.422
R55456 vp_n.n497 vp_n.n496 5.422
R55457 vp_n.n2058 vp_n.n2057 5.422
R55458 vp_n.n3711 vp_n.n3710 5.422
R55459 vp_n.n507 vp_n.n506 5.422
R55460 vp_n.n2068 vp_n.n2067 5.422
R55461 vp_n.n3721 vp_n.n3720 5.422
R55462 vp_n.n517 vp_n.n516 5.422
R55463 vp_n.n2078 vp_n.n2077 5.422
R55464 vp_n.n3731 vp_n.n3730 5.422
R55465 vp_n.n527 vp_n.n526 5.422
R55466 vp_n.n2088 vp_n.n2087 5.422
R55467 vp_n.n3741 vp_n.n3740 5.422
R55468 vp_n.n537 vp_n.n536 5.422
R55469 vp_n.n2098 vp_n.n2097 5.422
R55470 vp_n.n3751 vp_n.n3750 5.422
R55471 vp_n.n547 vp_n.n546 5.422
R55472 vp_n.n2108 vp_n.n2107 5.422
R55473 vp_n.n3761 vp_n.n3760 5.422
R55474 vp_n.n557 vp_n.n556 5.422
R55475 vp_n.n2118 vp_n.n2117 5.422
R55476 vp_n.n3771 vp_n.n3770 5.422
R55477 vp_n.n567 vp_n.n566 5.422
R55478 vp_n.n2128 vp_n.n2127 5.422
R55479 vp_n.n3781 vp_n.n3780 5.422
R55480 vp_n.n577 vp_n.n576 5.422
R55481 vp_n.n2138 vp_n.n2137 5.422
R55482 vp_n.n3791 vp_n.n3790 5.422
R55483 vp_n.n587 vp_n.n586 5.422
R55484 vp_n.n2148 vp_n.n2147 5.422
R55485 vp_n.n3801 vp_n.n3800 5.422
R55486 vp_n.n597 vp_n.n596 5.422
R55487 vp_n.n2158 vp_n.n2157 5.422
R55488 vp_n.n3811 vp_n.n3810 5.422
R55489 vp_n.n607 vp_n.n606 5.422
R55490 vp_n.n2168 vp_n.n2167 5.422
R55491 vp_n.n3821 vp_n.n3820 5.422
R55492 vp_n.n617 vp_n.n616 5.422
R55493 vp_n.n2178 vp_n.n2177 5.422
R55494 vp_n.n3831 vp_n.n3830 5.422
R55495 vp_n.n627 vp_n.n626 5.422
R55496 vp_n.n2188 vp_n.n2187 5.422
R55497 vp_n.n3841 vp_n.n3840 5.422
R55498 vp_n.n637 vp_n.n636 5.422
R55499 vp_n.n2198 vp_n.n2197 5.422
R55500 vp_n.n3851 vp_n.n3850 5.422
R55501 vp_n.n647 vp_n.n646 5.422
R55502 vp_n.n2208 vp_n.n2207 5.422
R55503 vp_n.n3861 vp_n.n3860 5.422
R55504 vp_n.n657 vp_n.n656 5.422
R55505 vp_n.n2218 vp_n.n2217 5.422
R55506 vp_n.n3871 vp_n.n3870 5.422
R55507 vp_n.n667 vp_n.n666 5.422
R55508 vp_n.n2228 vp_n.n2227 5.422
R55509 vp_n.n3881 vp_n.n3880 5.422
R55510 vp_n.n677 vp_n.n676 5.422
R55511 vp_n.n2238 vp_n.n2237 5.422
R55512 vp_n.n3891 vp_n.n3890 5.422
R55513 vp_n.n687 vp_n.n686 5.422
R55514 vp_n.n2248 vp_n.n2247 5.422
R55515 vp_n.n3901 vp_n.n3900 5.422
R55516 vp_n.n697 vp_n.n696 5.422
R55517 vp_n.n2258 vp_n.n2257 5.422
R55518 vp_n.n3911 vp_n.n3910 5.422
R55519 vp_n.n707 vp_n.n706 5.422
R55520 vp_n.n2268 vp_n.n2267 5.422
R55521 vp_n.n3921 vp_n.n3920 5.422
R55522 vp_n.n717 vp_n.n716 5.422
R55523 vp_n.n2278 vp_n.n2277 5.422
R55524 vp_n.n3931 vp_n.n3930 5.422
R55525 vp_n.n727 vp_n.n726 5.422
R55526 vp_n.n2288 vp_n.n2287 5.422
R55527 vp_n.n3941 vp_n.n3940 5.422
R55528 vp_n.n737 vp_n.n736 5.422
R55529 vp_n.n2298 vp_n.n2297 5.422
R55530 vp_n.n3951 vp_n.n3950 5.422
R55531 vp_n.n747 vp_n.n746 5.422
R55532 vp_n.n2308 vp_n.n2307 5.422
R55533 vp_n.n3961 vp_n.n3960 5.422
R55534 vp_n.n757 vp_n.n756 5.422
R55535 vp_n.n2318 vp_n.n2317 5.422
R55536 vp_n.n3971 vp_n.n3970 5.422
R55537 vp_n.n767 vp_n.n766 5.422
R55538 vp_n.n2328 vp_n.n2327 5.422
R55539 vp_n.n3981 vp_n.n3980 5.422
R55540 vp_n.n777 vp_n.n776 5.422
R55541 vp_n.n2338 vp_n.n2337 5.422
R55542 vp_n.n3991 vp_n.n3990 5.422
R55543 vp_n.n787 vp_n.n786 5.422
R55544 vp_n.n2348 vp_n.n2347 5.422
R55545 vp_n.n4001 vp_n.n4000 5.422
R55546 vp_n.n797 vp_n.n796 5.422
R55547 vp_n.n2358 vp_n.n2357 5.422
R55548 vp_n.n4011 vp_n.n4010 5.422
R55549 vp_n.n807 vp_n.n806 5.422
R55550 vp_n.n2368 vp_n.n2367 5.422
R55551 vp_n.n4021 vp_n.n4020 5.422
R55552 vp_n.n817 vp_n.n816 5.422
R55553 vp_n.n2378 vp_n.n2377 5.422
R55554 vp_n.n4031 vp_n.n4030 5.422
R55555 vp_n.n827 vp_n.n826 5.422
R55556 vp_n.n2388 vp_n.n2387 5.422
R55557 vp_n.n4041 vp_n.n4040 5.422
R55558 vp_n.n837 vp_n.n836 5.422
R55559 vp_n.n2398 vp_n.n2397 5.422
R55560 vp_n.n4051 vp_n.n4050 5.422
R55561 vp_n.n847 vp_n.n846 5.422
R55562 vp_n.n2408 vp_n.n2407 5.422
R55563 vp_n.n4061 vp_n.n4060 5.422
R55564 vp_n.n857 vp_n.n856 5.422
R55565 vp_n.n2418 vp_n.n2417 5.422
R55566 vp_n.n4071 vp_n.n4070 5.422
R55567 vp_n.n867 vp_n.n866 5.422
R55568 vp_n.n2428 vp_n.n2427 5.422
R55569 vp_n.n4081 vp_n.n4080 5.422
R55570 vp_n.n877 vp_n.n876 5.422
R55571 vp_n.n2438 vp_n.n2437 5.422
R55572 vp_n.n4091 vp_n.n4090 5.422
R55573 vp_n.n887 vp_n.n886 5.422
R55574 vp_n.n2448 vp_n.n2447 5.422
R55575 vp_n.n4101 vp_n.n4100 5.422
R55576 vp_n.n897 vp_n.n896 5.422
R55577 vp_n.n2458 vp_n.n2457 5.422
R55578 vp_n.n4111 vp_n.n4110 5.422
R55579 vp_n.n907 vp_n.n906 5.422
R55580 vp_n.n2468 vp_n.n2467 5.422
R55581 vp_n.n4121 vp_n.n4120 5.422
R55582 vp_n.n917 vp_n.n916 5.422
R55583 vp_n.n2478 vp_n.n2477 5.422
R55584 vp_n.n4131 vp_n.n4130 5.422
R55585 vp_n.n927 vp_n.n926 5.422
R55586 vp_n.n2488 vp_n.n2487 5.422
R55587 vp_n.n4141 vp_n.n4140 5.422
R55588 vp_n.n937 vp_n.n936 5.422
R55589 vp_n.n2498 vp_n.n2497 5.422
R55590 vp_n.n4151 vp_n.n4150 5.422
R55591 vp_n.n947 vp_n.n946 5.422
R55592 vp_n.n2508 vp_n.n2507 5.422
R55593 vp_n.n4161 vp_n.n4160 5.422
R55594 vp_n.n957 vp_n.n956 5.422
R55595 vp_n.n2518 vp_n.n2517 5.422
R55596 vp_n.n4171 vp_n.n4170 5.422
R55597 vp_n.n967 vp_n.n966 5.422
R55598 vp_n.n2528 vp_n.n2527 5.422
R55599 vp_n.n4181 vp_n.n4180 5.422
R55600 vp_n.n977 vp_n.n976 5.422
R55601 vp_n.n2538 vp_n.n2537 5.422
R55602 vp_n.n4191 vp_n.n4190 5.422
R55603 vp_n.n987 vp_n.n986 5.422
R55604 vp_n.n2548 vp_n.n2547 5.422
R55605 vp_n.n4201 vp_n.n4200 5.422
R55606 vp_n.n997 vp_n.n996 5.422
R55607 vp_n.n2558 vp_n.n2557 5.422
R55608 vp_n.n4211 vp_n.n4210 5.422
R55609 vp_n.n1007 vp_n.n1006 5.422
R55610 vp_n.n2568 vp_n.n2567 5.422
R55611 vp_n.n4221 vp_n.n4220 5.422
R55612 vp_n.n1017 vp_n.n1016 5.422
R55613 vp_n.n2578 vp_n.n2577 5.422
R55614 vp_n.n4231 vp_n.n4230 5.422
R55615 vp_n.n1027 vp_n.n1026 5.422
R55616 vp_n.n2588 vp_n.n2587 5.422
R55617 vp_n.n4241 vp_n.n4240 5.422
R55618 vp_n.n1037 vp_n.n1036 5.422
R55619 vp_n.n2598 vp_n.n2597 5.422
R55620 vp_n.n4251 vp_n.n4250 5.422
R55621 vp_n.n1047 vp_n.n1046 5.422
R55622 vp_n.n2608 vp_n.n2607 5.422
R55623 vp_n.n4261 vp_n.n4260 5.422
R55624 vp_n.n1057 vp_n.n1056 5.422
R55625 vp_n.n2618 vp_n.n2617 5.422
R55626 vp_n.n4271 vp_n.n4270 5.422
R55627 vp_n.n1067 vp_n.n1066 5.422
R55628 vp_n.n2628 vp_n.n2627 5.422
R55629 vp_n.n4281 vp_n.n4280 5.422
R55630 vp_n.n1077 vp_n.n1076 5.422
R55631 vp_n.n2638 vp_n.n2637 5.422
R55632 vp_n.n4291 vp_n.n4290 5.422
R55633 vp_n.n1087 vp_n.n1086 5.422
R55634 vp_n.n2648 vp_n.n2647 5.422
R55635 vp_n.n4301 vp_n.n4300 5.422
R55636 vp_n.n1097 vp_n.n1096 5.422
R55637 vp_n.n2658 vp_n.n2657 5.422
R55638 vp_n.n4311 vp_n.n4310 5.422
R55639 vp_n.n1107 vp_n.n1106 5.422
R55640 vp_n.n2668 vp_n.n2667 5.422
R55641 vp_n.n4321 vp_n.n4320 5.422
R55642 vp_n.n1117 vp_n.n1116 5.422
R55643 vp_n.n2678 vp_n.n2677 5.422
R55644 vp_n.n4331 vp_n.n4330 5.422
R55645 vp_n.n1127 vp_n.n1126 5.422
R55646 vp_n.n2688 vp_n.n2687 5.422
R55647 vp_n.n4341 vp_n.n4340 5.422
R55648 vp_n.n1137 vp_n.n1136 5.422
R55649 vp_n.n2698 vp_n.n2697 5.422
R55650 vp_n.n4351 vp_n.n4350 5.422
R55651 vp_n.n1147 vp_n.n1146 5.422
R55652 vp_n.n2708 vp_n.n2707 5.422
R55653 vp_n.n4361 vp_n.n4360 5.422
R55654 vp_n.n1157 vp_n.n1156 5.422
R55655 vp_n.n2718 vp_n.n2717 5.422
R55656 vp_n.n4371 vp_n.n4370 5.422
R55657 vp_n.n1167 vp_n.n1166 5.422
R55658 vp_n.n2728 vp_n.n2727 5.422
R55659 vp_n.n4381 vp_n.n4380 5.422
R55660 vp_n.n1177 vp_n.n1176 5.422
R55661 vp_n.n2738 vp_n.n2737 5.422
R55662 vp_n.n4391 vp_n.n4390 5.422
R55663 vp_n.n1187 vp_n.n1186 5.422
R55664 vp_n.n2748 vp_n.n2747 5.422
R55665 vp_n.n4401 vp_n.n4400 5.422
R55666 vp_n.n1197 vp_n.n1196 5.422
R55667 vp_n.n2758 vp_n.n2757 5.422
R55668 vp_n.n4411 vp_n.n4410 5.422
R55669 vp_n.n1207 vp_n.n1206 5.422
R55670 vp_n.n2768 vp_n.n2767 5.422
R55671 vp_n.n4421 vp_n.n4420 5.422
R55672 vp_n.n1217 vp_n.n1216 5.422
R55673 vp_n.n2778 vp_n.n2777 5.422
R55674 vp_n.n4431 vp_n.n4430 5.422
R55675 vp_n.n1227 vp_n.n1226 5.422
R55676 vp_n.n2788 vp_n.n2787 5.422
R55677 vp_n.n4441 vp_n.n4440 5.422
R55678 vp_n.n1237 vp_n.n1236 5.422
R55679 vp_n.n2798 vp_n.n2797 5.422
R55680 vp_n.n4451 vp_n.n4450 5.422
R55681 vp_n.n1247 vp_n.n1246 5.422
R55682 vp_n.n2808 vp_n.n2807 5.422
R55683 vp_n.n4461 vp_n.n4460 5.422
R55684 vp_n.n1257 vp_n.n1256 5.422
R55685 vp_n.n2818 vp_n.n2817 5.422
R55686 vp_n.n4471 vp_n.n4470 5.422
R55687 vp_n.n1267 vp_n.n1266 5.422
R55688 vp_n.n2828 vp_n.n2827 5.422
R55689 vp_n.n4481 vp_n.n4480 5.422
R55690 vp_n.n1277 vp_n.n1276 5.422
R55691 vp_n.n2838 vp_n.n2837 5.422
R55692 vp_n.n4491 vp_n.n4490 5.422
R55693 vp_n.n1287 vp_n.n1286 5.422
R55694 vp_n.n2848 vp_n.n2847 5.422
R55695 vp_n.n4501 vp_n.n4500 5.422
R55696 vp_n.n1297 vp_n.n1296 5.422
R55697 vp_n.n2858 vp_n.n2857 5.422
R55698 vp_n.n4511 vp_n.n4510 5.422
R55699 vp_n.n1307 vp_n.n1306 5.422
R55700 vp_n.n2868 vp_n.n2867 5.422
R55701 vp_n.n4521 vp_n.n4520 5.422
R55702 vp_n.n1317 vp_n.n1316 5.422
R55703 vp_n.n2878 vp_n.n2877 5.422
R55704 vp_n.n4531 vp_n.n4530 5.422
R55705 vp_n.n1327 vp_n.n1326 5.422
R55706 vp_n.n2888 vp_n.n2887 5.422
R55707 vp_n.n4541 vp_n.n4540 5.422
R55708 vp_n.n1337 vp_n.n1336 5.422
R55709 vp_n.n2898 vp_n.n2897 5.422
R55710 vp_n.n4551 vp_n.n4550 5.422
R55711 vp_n.n1347 vp_n.n1346 5.422
R55712 vp_n.n2908 vp_n.n2907 5.422
R55713 vp_n.n4561 vp_n.n4560 5.422
R55714 vp_n.n1357 vp_n.n1356 5.422
R55715 vp_n.n2918 vp_n.n2917 5.422
R55716 vp_n.n4571 vp_n.n4570 5.422
R55717 vp_n.n1367 vp_n.n1366 5.422
R55718 vp_n.n2928 vp_n.n2927 5.422
R55719 vp_n.n4581 vp_n.n4580 5.422
R55720 vp_n.n1377 vp_n.n1376 5.422
R55721 vp_n.n2938 vp_n.n2937 5.422
R55722 vp_n.n4591 vp_n.n4590 5.422
R55723 vp_n.n1387 vp_n.n1386 5.422
R55724 vp_n.n2948 vp_n.n2947 5.422
R55725 vp_n.n4601 vp_n.n4600 5.422
R55726 vp_n.n1397 vp_n.n1396 5.422
R55727 vp_n.n2958 vp_n.n2957 5.422
R55728 vp_n.n4611 vp_n.n4610 5.422
R55729 vp_n.n1407 vp_n.n1406 5.422
R55730 vp_n.n2968 vp_n.n2967 5.422
R55731 vp_n.n4621 vp_n.n4620 5.422
R55732 vp_n.n1417 vp_n.n1416 5.422
R55733 vp_n.n2978 vp_n.n2977 5.422
R55734 vp_n.n4631 vp_n.n4630 5.422
R55735 vp_n.n1427 vp_n.n1426 5.422
R55736 vp_n.n2988 vp_n.n2987 5.422
R55737 vp_n.n4641 vp_n.n4640 5.422
R55738 vp_n.n1437 vp_n.n1436 5.422
R55739 vp_n.n2998 vp_n.n2997 5.422
R55740 vp_n.n4651 vp_n.n4650 5.422
R55741 vp_n.n1447 vp_n.n1446 5.422
R55742 vp_n.n3008 vp_n.n3007 5.422
R55743 vp_n.n4661 vp_n.n4660 5.422
R55744 vp_n.n1457 vp_n.n1456 5.422
R55745 vp_n.n3018 vp_n.n3017 5.422
R55746 vp_n.n4671 vp_n.n4670 5.422
R55747 vp_n.n1467 vp_n.n1466 5.422
R55748 vp_n.n3028 vp_n.n3027 5.422
R55749 vp_n.n4681 vp_n.n4680 5.422
R55750 vp_n.n1477 vp_n.n1476 5.422
R55751 vp_n.n3038 vp_n.n3037 5.422
R55752 vp_n.n4691 vp_n.n4690 5.422
R55753 vp_n.n1487 vp_n.n1486 5.422
R55754 vp_n.n1497 vp_n.n1496 5.422
R55755 vp_n.n4701 vp_n.n4700 5.422
R55756 vp_n.n3048 vp_n.n3047 5.422
R55757 vp_n.n1568 vp_n.n1567 5.422
R55758 vp_n.n3221 vp_n.n3220 5.422
R55759 vp_n.n3211 vp_n.n3210 5.422
R55760 vp_n.n1551 vp_n.n1550 1.238
R55761 vp_n.n3204 vp_n.n3203 1.238
R55762 vp_n.n3152 vp_n.n3151 1.208
R55763 vp_n.n4805 vp_n.n4804 1.208
R55764 vp_n.n1550 vp_n.n1549 1.043
R55765 vp_n.n1549 vp_n.n1548 1.043
R55766 vp_n.n1548 vp_n.n1547 1.043
R55767 vp_n.n1547 vp_n.n1546 1.043
R55768 vp_n.n1546 vp_n.n1545 1.043
R55769 vp_n.n1545 vp_n.n1544 1.043
R55770 vp_n.n1544 vp_n.n1543 1.043
R55771 vp_n.n1543 vp_n.n1542 1.043
R55772 vp_n.n1542 vp_n.n1541 1.043
R55773 vp_n.n1541 vp_n.n1540 1.043
R55774 vp_n.n1540 vp_n.n1539 1.043
R55775 vp_n.n1539 vp_n.n1538 1.043
R55776 vp_n.n1538 vp_n.n1537 1.043
R55777 vp_n.n1537 vp_n.n1536 1.043
R55778 vp_n.n1536 vp_n.n1535 1.043
R55779 vp_n.n1535 vp_n.n1534 1.043
R55780 vp_n.n1534 vp_n.n1533 1.043
R55781 vp_n.n1533 vp_n.n1532 1.043
R55782 vp_n.n1532 vp_n.n1531 1.043
R55783 vp_n.n1531 vp_n.n1530 1.043
R55784 vp_n.n1530 vp_n.n1529 1.043
R55785 vp_n.n1529 vp_n.n1528 1.043
R55786 vp_n.n1528 vp_n.n1527 1.043
R55787 vp_n.n1527 vp_n.n1526 1.043
R55788 vp_n.n1526 vp_n.n1525 1.043
R55789 vp_n.n1525 vp_n.n1524 1.043
R55790 vp_n.n1524 vp_n.n1523 1.043
R55791 vp_n.n1523 vp_n.n1522 1.043
R55792 vp_n.n1522 vp_n.n1521 1.043
R55793 vp_n.n1521 vp_n.n1520 1.043
R55794 vp_n.n1520 vp_n.n1519 1.043
R55795 vp_n.n1519 vp_n.n1518 1.043
R55796 vp_n.n1518 vp_n.n1517 1.043
R55797 vp_n.n1517 vp_n.n1516 1.043
R55798 vp_n.n1516 vp_n.n1515 1.043
R55799 vp_n.n1515 vp_n.n1514 1.043
R55800 vp_n.n1514 vp_n.n1513 1.043
R55801 vp_n.n1513 vp_n.n1512 1.043
R55802 vp_n.n1512 vp_n.n1511 1.043
R55803 vp_n.n1511 vp_n.n1510 1.043
R55804 vp_n.n1510 vp_n.n1509 1.043
R55805 vp_n.n1509 vp_n.n1508 1.043
R55806 vp_n.n1508 vp_n.n1507 1.043
R55807 vp_n.n1507 vp_n.n1506 1.043
R55808 vp_n.n1506 vp_n.n1505 1.043
R55809 vp_n.n1505 vp_n.n1504 1.043
R55810 vp_n.n1504 vp_n.n1503 1.043
R55811 vp_n.n1503 vp_n.n1502 1.043
R55812 vp_n.n1502 vp_n.n1501 1.043
R55813 vp_n.n3053 vp_n.n3052 1.043
R55814 vp_n.n3054 vp_n.n3053 1.043
R55815 vp_n.n3055 vp_n.n3054 1.043
R55816 vp_n.n3056 vp_n.n3055 1.043
R55817 vp_n.n3057 vp_n.n3056 1.043
R55818 vp_n.n3058 vp_n.n3057 1.043
R55819 vp_n.n3059 vp_n.n3058 1.043
R55820 vp_n.n3060 vp_n.n3059 1.043
R55821 vp_n.n3061 vp_n.n3060 1.043
R55822 vp_n.n3062 vp_n.n3061 1.043
R55823 vp_n.n3063 vp_n.n3062 1.043
R55824 vp_n.n3064 vp_n.n3063 1.043
R55825 vp_n.n3065 vp_n.n3064 1.043
R55826 vp_n.n3066 vp_n.n3065 1.043
R55827 vp_n.n3067 vp_n.n3066 1.043
R55828 vp_n.n3068 vp_n.n3067 1.043
R55829 vp_n.n3069 vp_n.n3068 1.043
R55830 vp_n.n3070 vp_n.n3069 1.043
R55831 vp_n.n3071 vp_n.n3070 1.043
R55832 vp_n.n3072 vp_n.n3071 1.043
R55833 vp_n.n3073 vp_n.n3072 1.043
R55834 vp_n.n3074 vp_n.n3073 1.043
R55835 vp_n.n3075 vp_n.n3074 1.043
R55836 vp_n.n3076 vp_n.n3075 1.043
R55837 vp_n.n3077 vp_n.n3076 1.043
R55838 vp_n.n3078 vp_n.n3077 1.043
R55839 vp_n.n3079 vp_n.n3078 1.043
R55840 vp_n.n3080 vp_n.n3079 1.043
R55841 vp_n.n3081 vp_n.n3080 1.043
R55842 vp_n.n3082 vp_n.n3081 1.043
R55843 vp_n.n3083 vp_n.n3082 1.043
R55844 vp_n.n3084 vp_n.n3083 1.043
R55845 vp_n.n3085 vp_n.n3084 1.043
R55846 vp_n.n3086 vp_n.n3085 1.043
R55847 vp_n.n3087 vp_n.n3086 1.043
R55848 vp_n.n3088 vp_n.n3087 1.043
R55849 vp_n.n3089 vp_n.n3088 1.043
R55850 vp_n.n3090 vp_n.n3089 1.043
R55851 vp_n.n3091 vp_n.n3090 1.043
R55852 vp_n.n3092 vp_n.n3091 1.043
R55853 vp_n.n3093 vp_n.n3092 1.043
R55854 vp_n.n3094 vp_n.n3093 1.043
R55855 vp_n.n3095 vp_n.n3094 1.043
R55856 vp_n.n3096 vp_n.n3095 1.043
R55857 vp_n.n3097 vp_n.n3096 1.043
R55858 vp_n.n3098 vp_n.n3097 1.043
R55859 vp_n.n3099 vp_n.n3098 1.043
R55860 vp_n.n3100 vp_n.n3099 1.043
R55861 vp_n.n3101 vp_n.n3100 1.043
R55862 vp_n.n3102 vp_n.n3101 1.043
R55863 vp_n.n3103 vp_n.n3102 1.043
R55864 vp_n.n3104 vp_n.n3103 1.043
R55865 vp_n.n3105 vp_n.n3104 1.043
R55866 vp_n.n3106 vp_n.n3105 1.043
R55867 vp_n.n3107 vp_n.n3106 1.043
R55868 vp_n.n3108 vp_n.n3107 1.043
R55869 vp_n.n3109 vp_n.n3108 1.043
R55870 vp_n.n3110 vp_n.n3109 1.043
R55871 vp_n.n3111 vp_n.n3110 1.043
R55872 vp_n.n3112 vp_n.n3111 1.043
R55873 vp_n.n3113 vp_n.n3112 1.043
R55874 vp_n.n3114 vp_n.n3113 1.043
R55875 vp_n.n3115 vp_n.n3114 1.043
R55876 vp_n.n3116 vp_n.n3115 1.043
R55877 vp_n.n3117 vp_n.n3116 1.043
R55878 vp_n.n3118 vp_n.n3117 1.043
R55879 vp_n.n3119 vp_n.n3118 1.043
R55880 vp_n.n3120 vp_n.n3119 1.043
R55881 vp_n.n3121 vp_n.n3120 1.043
R55882 vp_n.n3122 vp_n.n3121 1.043
R55883 vp_n.n3123 vp_n.n3122 1.043
R55884 vp_n.n3124 vp_n.n3123 1.043
R55885 vp_n.n3125 vp_n.n3124 1.043
R55886 vp_n.n3126 vp_n.n3125 1.043
R55887 vp_n.n3127 vp_n.n3126 1.043
R55888 vp_n.n3128 vp_n.n3127 1.043
R55889 vp_n.n3129 vp_n.n3128 1.043
R55890 vp_n.n3130 vp_n.n3129 1.043
R55891 vp_n.n3131 vp_n.n3130 1.043
R55892 vp_n.n3132 vp_n.n3131 1.043
R55893 vp_n.n3133 vp_n.n3132 1.043
R55894 vp_n.n3134 vp_n.n3133 1.043
R55895 vp_n.n3135 vp_n.n3134 1.043
R55896 vp_n.n3136 vp_n.n3135 1.043
R55897 vp_n.n3137 vp_n.n3136 1.043
R55898 vp_n.n3138 vp_n.n3137 1.043
R55899 vp_n.n3139 vp_n.n3138 1.043
R55900 vp_n.n3140 vp_n.n3139 1.043
R55901 vp_n.n3141 vp_n.n3140 1.043
R55902 vp_n.n3142 vp_n.n3141 1.043
R55903 vp_n.n3143 vp_n.n3142 1.043
R55904 vp_n.n3144 vp_n.n3143 1.043
R55905 vp_n.n3145 vp_n.n3144 1.043
R55906 vp_n.n3146 vp_n.n3145 1.043
R55907 vp_n.n3147 vp_n.n3146 1.043
R55908 vp_n.n3148 vp_n.n3147 1.043
R55909 vp_n.n3149 vp_n.n3148 1.043
R55910 vp_n.n3150 vp_n.n3149 1.043
R55911 vp_n.n3151 vp_n.n3150 1.043
R55912 vp_n.n3203 vp_n.n3202 1.043
R55913 vp_n.n3202 vp_n.n3201 1.043
R55914 vp_n.n3201 vp_n.n3200 1.043
R55915 vp_n.n3200 vp_n.n3199 1.043
R55916 vp_n.n3199 vp_n.n3198 1.043
R55917 vp_n.n3198 vp_n.n3197 1.043
R55918 vp_n.n3197 vp_n.n3196 1.043
R55919 vp_n.n3196 vp_n.n3195 1.043
R55920 vp_n.n3195 vp_n.n3194 1.043
R55921 vp_n.n3194 vp_n.n3193 1.043
R55922 vp_n.n3193 vp_n.n3192 1.043
R55923 vp_n.n3192 vp_n.n3191 1.043
R55924 vp_n.n3191 vp_n.n3190 1.043
R55925 vp_n.n3190 vp_n.n3189 1.043
R55926 vp_n.n3189 vp_n.n3188 1.043
R55927 vp_n.n3188 vp_n.n3187 1.043
R55928 vp_n.n3187 vp_n.n3186 1.043
R55929 vp_n.n3186 vp_n.n3185 1.043
R55930 vp_n.n3185 vp_n.n3184 1.043
R55931 vp_n.n3184 vp_n.n3183 1.043
R55932 vp_n.n3183 vp_n.n3182 1.043
R55933 vp_n.n3182 vp_n.n3181 1.043
R55934 vp_n.n3181 vp_n.n3180 1.043
R55935 vp_n.n3180 vp_n.n3179 1.043
R55936 vp_n.n3179 vp_n.n3178 1.043
R55937 vp_n.n3178 vp_n.n3177 1.043
R55938 vp_n.n3177 vp_n.n3176 1.043
R55939 vp_n.n3176 vp_n.n3175 1.043
R55940 vp_n.n3175 vp_n.n3174 1.043
R55941 vp_n.n3174 vp_n.n3173 1.043
R55942 vp_n.n3173 vp_n.n3172 1.043
R55943 vp_n.n3172 vp_n.n3171 1.043
R55944 vp_n.n3171 vp_n.n3170 1.043
R55945 vp_n.n3170 vp_n.n3169 1.043
R55946 vp_n.n3169 vp_n.n3168 1.043
R55947 vp_n.n3168 vp_n.n3167 1.043
R55948 vp_n.n3167 vp_n.n3166 1.043
R55949 vp_n.n3166 vp_n.n3165 1.043
R55950 vp_n.n3165 vp_n.n3164 1.043
R55951 vp_n.n3164 vp_n.n3163 1.043
R55952 vp_n.n3163 vp_n.n3162 1.043
R55953 vp_n.n3162 vp_n.n3161 1.043
R55954 vp_n.n3161 vp_n.n3160 1.043
R55955 vp_n.n3160 vp_n.n3159 1.043
R55956 vp_n.n3159 vp_n.n3158 1.043
R55957 vp_n.n3158 vp_n.n3157 1.043
R55958 vp_n.n3157 vp_n.n3156 1.043
R55959 vp_n.n3156 vp_n.n3155 1.043
R55960 vp_n.n3155 vp_n.n3154 1.043
R55961 vp_n.n4706 vp_n.n4705 1.043
R55962 vp_n.n4707 vp_n.n4706 1.043
R55963 vp_n.n4708 vp_n.n4707 1.043
R55964 vp_n.n4709 vp_n.n4708 1.043
R55965 vp_n.n4710 vp_n.n4709 1.043
R55966 vp_n.n4711 vp_n.n4710 1.043
R55967 vp_n.n4712 vp_n.n4711 1.043
R55968 vp_n.n4713 vp_n.n4712 1.043
R55969 vp_n.n4714 vp_n.n4713 1.043
R55970 vp_n.n4715 vp_n.n4714 1.043
R55971 vp_n.n4716 vp_n.n4715 1.043
R55972 vp_n.n4717 vp_n.n4716 1.043
R55973 vp_n.n4718 vp_n.n4717 1.043
R55974 vp_n.n4719 vp_n.n4718 1.043
R55975 vp_n.n4720 vp_n.n4719 1.043
R55976 vp_n.n4721 vp_n.n4720 1.043
R55977 vp_n.n4722 vp_n.n4721 1.043
R55978 vp_n.n4723 vp_n.n4722 1.043
R55979 vp_n.n4724 vp_n.n4723 1.043
R55980 vp_n.n4725 vp_n.n4724 1.043
R55981 vp_n.n4726 vp_n.n4725 1.043
R55982 vp_n.n4727 vp_n.n4726 1.043
R55983 vp_n.n4728 vp_n.n4727 1.043
R55984 vp_n.n4729 vp_n.n4728 1.043
R55985 vp_n.n4730 vp_n.n4729 1.043
R55986 vp_n.n4731 vp_n.n4730 1.043
R55987 vp_n.n4732 vp_n.n4731 1.043
R55988 vp_n.n4733 vp_n.n4732 1.043
R55989 vp_n.n4734 vp_n.n4733 1.043
R55990 vp_n.n4735 vp_n.n4734 1.043
R55991 vp_n.n4736 vp_n.n4735 1.043
R55992 vp_n.n4737 vp_n.n4736 1.043
R55993 vp_n.n4738 vp_n.n4737 1.043
R55994 vp_n.n4739 vp_n.n4738 1.043
R55995 vp_n.n4740 vp_n.n4739 1.043
R55996 vp_n.n4741 vp_n.n4740 1.043
R55997 vp_n.n4742 vp_n.n4741 1.043
R55998 vp_n.n4743 vp_n.n4742 1.043
R55999 vp_n.n4744 vp_n.n4743 1.043
R56000 vp_n.n4745 vp_n.n4744 1.043
R56001 vp_n.n4746 vp_n.n4745 1.043
R56002 vp_n.n4747 vp_n.n4746 1.043
R56003 vp_n.n4748 vp_n.n4747 1.043
R56004 vp_n.n4749 vp_n.n4748 1.043
R56005 vp_n.n4750 vp_n.n4749 1.043
R56006 vp_n.n4751 vp_n.n4750 1.043
R56007 vp_n.n4752 vp_n.n4751 1.043
R56008 vp_n.n4753 vp_n.n4752 1.043
R56009 vp_n.n4754 vp_n.n4753 1.043
R56010 vp_n.n4755 vp_n.n4754 1.043
R56011 vp_n.n4756 vp_n.n4755 1.043
R56012 vp_n.n4757 vp_n.n4756 1.043
R56013 vp_n.n4758 vp_n.n4757 1.043
R56014 vp_n.n4759 vp_n.n4758 1.043
R56015 vp_n.n4760 vp_n.n4759 1.043
R56016 vp_n.n4761 vp_n.n4760 1.043
R56017 vp_n.n4762 vp_n.n4761 1.043
R56018 vp_n.n4763 vp_n.n4762 1.043
R56019 vp_n.n4764 vp_n.n4763 1.043
R56020 vp_n.n4765 vp_n.n4764 1.043
R56021 vp_n.n4766 vp_n.n4765 1.043
R56022 vp_n.n4767 vp_n.n4766 1.043
R56023 vp_n.n4768 vp_n.n4767 1.043
R56024 vp_n.n4769 vp_n.n4768 1.043
R56025 vp_n.n4770 vp_n.n4769 1.043
R56026 vp_n.n4771 vp_n.n4770 1.043
R56027 vp_n.n4772 vp_n.n4771 1.043
R56028 vp_n.n4773 vp_n.n4772 1.043
R56029 vp_n.n4774 vp_n.n4773 1.043
R56030 vp_n.n4775 vp_n.n4774 1.043
R56031 vp_n.n4776 vp_n.n4775 1.043
R56032 vp_n.n4777 vp_n.n4776 1.043
R56033 vp_n.n4778 vp_n.n4777 1.043
R56034 vp_n.n4779 vp_n.n4778 1.043
R56035 vp_n.n4780 vp_n.n4779 1.043
R56036 vp_n.n4781 vp_n.n4780 1.043
R56037 vp_n.n4782 vp_n.n4781 1.043
R56038 vp_n.n4783 vp_n.n4782 1.043
R56039 vp_n.n4784 vp_n.n4783 1.043
R56040 vp_n.n4785 vp_n.n4784 1.043
R56041 vp_n.n4786 vp_n.n4785 1.043
R56042 vp_n.n4787 vp_n.n4786 1.043
R56043 vp_n.n4788 vp_n.n4787 1.043
R56044 vp_n.n4789 vp_n.n4788 1.043
R56045 vp_n.n4790 vp_n.n4789 1.043
R56046 vp_n.n4791 vp_n.n4790 1.043
R56047 vp_n.n4792 vp_n.n4791 1.043
R56048 vp_n.n4793 vp_n.n4792 1.043
R56049 vp_n.n4794 vp_n.n4793 1.043
R56050 vp_n.n4795 vp_n.n4794 1.043
R56051 vp_n.n4796 vp_n.n4795 1.043
R56052 vp_n.n4797 vp_n.n4796 1.043
R56053 vp_n.n4798 vp_n.n4797 1.043
R56054 vp_n.n4799 vp_n.n4798 1.043
R56055 vp_n.n4800 vp_n.n4799 1.043
R56056 vp_n.n4801 vp_n.n4800 1.043
R56057 vp_n.n4802 vp_n.n4801 1.043
R56058 vp_n.n4803 vp_n.n4802 1.043
R56059 vp_n.n4804 vp_n.n4803 1.043
R56060 vp_n.n1 vp_n.n0 0.332
R56061 vp_n.n1552 vp_n.n1551 0.332
R56062 vp_n.n3205 vp_n.n3204 0.332
R56063 vp_n.n3153 vp_n.n1500 0.331
R56064 vp_n.n3152 vp_n.n3051 0.331
R56065 vp_n.n4805 vp_n.n4704 0.331
R56066 vp_n.n11 vp_n.n10 0.319
R56067 vp_n.n21 vp_n.n20 0.319
R56068 vp_n.n31 vp_n.n30 0.319
R56069 vp_n.n41 vp_n.n40 0.319
R56070 vp_n.n51 vp_n.n50 0.319
R56071 vp_n.n61 vp_n.n60 0.319
R56072 vp_n.n71 vp_n.n70 0.319
R56073 vp_n.n81 vp_n.n80 0.319
R56074 vp_n.n91 vp_n.n90 0.319
R56075 vp_n.n101 vp_n.n100 0.319
R56076 vp_n.n111 vp_n.n110 0.319
R56077 vp_n.n121 vp_n.n120 0.319
R56078 vp_n.n131 vp_n.n130 0.319
R56079 vp_n.n141 vp_n.n140 0.319
R56080 vp_n.n151 vp_n.n150 0.319
R56081 vp_n.n161 vp_n.n160 0.319
R56082 vp_n.n171 vp_n.n170 0.319
R56083 vp_n.n181 vp_n.n180 0.319
R56084 vp_n.n191 vp_n.n190 0.319
R56085 vp_n.n201 vp_n.n200 0.319
R56086 vp_n.n211 vp_n.n210 0.319
R56087 vp_n.n221 vp_n.n220 0.319
R56088 vp_n.n231 vp_n.n230 0.319
R56089 vp_n.n241 vp_n.n240 0.319
R56090 vp_n.n251 vp_n.n250 0.319
R56091 vp_n.n261 vp_n.n260 0.319
R56092 vp_n.n271 vp_n.n270 0.319
R56093 vp_n.n281 vp_n.n280 0.319
R56094 vp_n.n291 vp_n.n290 0.319
R56095 vp_n.n301 vp_n.n300 0.319
R56096 vp_n.n311 vp_n.n310 0.319
R56097 vp_n.n321 vp_n.n320 0.319
R56098 vp_n.n331 vp_n.n330 0.319
R56099 vp_n.n341 vp_n.n340 0.319
R56100 vp_n.n351 vp_n.n350 0.319
R56101 vp_n.n361 vp_n.n360 0.319
R56102 vp_n.n371 vp_n.n370 0.319
R56103 vp_n.n381 vp_n.n380 0.319
R56104 vp_n.n391 vp_n.n390 0.319
R56105 vp_n.n401 vp_n.n400 0.319
R56106 vp_n.n411 vp_n.n410 0.319
R56107 vp_n.n421 vp_n.n420 0.319
R56108 vp_n.n431 vp_n.n430 0.319
R56109 vp_n.n441 vp_n.n440 0.319
R56110 vp_n.n451 vp_n.n450 0.319
R56111 vp_n.n461 vp_n.n460 0.319
R56112 vp_n.n471 vp_n.n470 0.319
R56113 vp_n.n481 vp_n.n480 0.319
R56114 vp_n.n491 vp_n.n490 0.319
R56115 vp_n.n501 vp_n.n500 0.319
R56116 vp_n.n511 vp_n.n510 0.319
R56117 vp_n.n521 vp_n.n520 0.319
R56118 vp_n.n531 vp_n.n530 0.319
R56119 vp_n.n541 vp_n.n540 0.319
R56120 vp_n.n551 vp_n.n550 0.319
R56121 vp_n.n561 vp_n.n560 0.319
R56122 vp_n.n571 vp_n.n570 0.319
R56123 vp_n.n581 vp_n.n580 0.319
R56124 vp_n.n591 vp_n.n590 0.319
R56125 vp_n.n601 vp_n.n600 0.319
R56126 vp_n.n611 vp_n.n610 0.319
R56127 vp_n.n621 vp_n.n620 0.319
R56128 vp_n.n631 vp_n.n630 0.319
R56129 vp_n.n641 vp_n.n640 0.319
R56130 vp_n.n651 vp_n.n650 0.319
R56131 vp_n.n661 vp_n.n660 0.319
R56132 vp_n.n671 vp_n.n670 0.319
R56133 vp_n.n681 vp_n.n680 0.319
R56134 vp_n.n691 vp_n.n690 0.319
R56135 vp_n.n701 vp_n.n700 0.319
R56136 vp_n.n711 vp_n.n710 0.319
R56137 vp_n.n721 vp_n.n720 0.319
R56138 vp_n.n731 vp_n.n730 0.319
R56139 vp_n.n741 vp_n.n740 0.319
R56140 vp_n.n751 vp_n.n750 0.319
R56141 vp_n.n761 vp_n.n760 0.319
R56142 vp_n.n771 vp_n.n770 0.319
R56143 vp_n.n781 vp_n.n780 0.319
R56144 vp_n.n791 vp_n.n790 0.319
R56145 vp_n.n801 vp_n.n800 0.319
R56146 vp_n.n811 vp_n.n810 0.319
R56147 vp_n.n821 vp_n.n820 0.319
R56148 vp_n.n831 vp_n.n830 0.319
R56149 vp_n.n841 vp_n.n840 0.319
R56150 vp_n.n851 vp_n.n850 0.319
R56151 vp_n.n861 vp_n.n860 0.319
R56152 vp_n.n871 vp_n.n870 0.319
R56153 vp_n.n881 vp_n.n880 0.319
R56154 vp_n.n891 vp_n.n890 0.319
R56155 vp_n.n901 vp_n.n900 0.319
R56156 vp_n.n911 vp_n.n910 0.319
R56157 vp_n.n921 vp_n.n920 0.319
R56158 vp_n.n931 vp_n.n930 0.319
R56159 vp_n.n941 vp_n.n940 0.319
R56160 vp_n.n951 vp_n.n950 0.319
R56161 vp_n.n961 vp_n.n960 0.319
R56162 vp_n.n971 vp_n.n970 0.319
R56163 vp_n.n981 vp_n.n980 0.319
R56164 vp_n.n991 vp_n.n990 0.319
R56165 vp_n.n1001 vp_n.n1000 0.319
R56166 vp_n.n1011 vp_n.n1010 0.319
R56167 vp_n.n1021 vp_n.n1020 0.319
R56168 vp_n.n1031 vp_n.n1030 0.319
R56169 vp_n.n1041 vp_n.n1040 0.319
R56170 vp_n.n1051 vp_n.n1050 0.319
R56171 vp_n.n1061 vp_n.n1060 0.319
R56172 vp_n.n1071 vp_n.n1070 0.319
R56173 vp_n.n1081 vp_n.n1080 0.319
R56174 vp_n.n1091 vp_n.n1090 0.319
R56175 vp_n.n1101 vp_n.n1100 0.319
R56176 vp_n.n1111 vp_n.n1110 0.319
R56177 vp_n.n1121 vp_n.n1120 0.319
R56178 vp_n.n1131 vp_n.n1130 0.319
R56179 vp_n.n1141 vp_n.n1140 0.319
R56180 vp_n.n1151 vp_n.n1150 0.319
R56181 vp_n.n1161 vp_n.n1160 0.319
R56182 vp_n.n1171 vp_n.n1170 0.319
R56183 vp_n.n1181 vp_n.n1180 0.319
R56184 vp_n.n1191 vp_n.n1190 0.319
R56185 vp_n.n1201 vp_n.n1200 0.319
R56186 vp_n.n1211 vp_n.n1210 0.319
R56187 vp_n.n1221 vp_n.n1220 0.319
R56188 vp_n.n1231 vp_n.n1230 0.319
R56189 vp_n.n1241 vp_n.n1240 0.319
R56190 vp_n.n1251 vp_n.n1250 0.319
R56191 vp_n.n1261 vp_n.n1260 0.319
R56192 vp_n.n1271 vp_n.n1270 0.319
R56193 vp_n.n1281 vp_n.n1280 0.319
R56194 vp_n.n1291 vp_n.n1290 0.319
R56195 vp_n.n1301 vp_n.n1300 0.319
R56196 vp_n.n1311 vp_n.n1310 0.319
R56197 vp_n.n1321 vp_n.n1320 0.319
R56198 vp_n.n1331 vp_n.n1330 0.319
R56199 vp_n.n1341 vp_n.n1340 0.319
R56200 vp_n.n1351 vp_n.n1350 0.319
R56201 vp_n.n1361 vp_n.n1360 0.319
R56202 vp_n.n1371 vp_n.n1370 0.319
R56203 vp_n.n1381 vp_n.n1380 0.319
R56204 vp_n.n1391 vp_n.n1390 0.319
R56205 vp_n.n1401 vp_n.n1400 0.319
R56206 vp_n.n1411 vp_n.n1410 0.319
R56207 vp_n.n1421 vp_n.n1420 0.319
R56208 vp_n.n1431 vp_n.n1430 0.319
R56209 vp_n.n1441 vp_n.n1440 0.319
R56210 vp_n.n1451 vp_n.n1450 0.319
R56211 vp_n.n1461 vp_n.n1460 0.319
R56212 vp_n.n1471 vp_n.n1470 0.319
R56213 vp_n.n1481 vp_n.n1480 0.319
R56214 vp_n.n1491 vp_n.n1490 0.319
R56215 vp_n.n1562 vp_n.n1561 0.319
R56216 vp_n.n1572 vp_n.n1571 0.319
R56217 vp_n.n1582 vp_n.n1581 0.319
R56218 vp_n.n1592 vp_n.n1591 0.319
R56219 vp_n.n1602 vp_n.n1601 0.319
R56220 vp_n.n1612 vp_n.n1611 0.319
R56221 vp_n.n1622 vp_n.n1621 0.319
R56222 vp_n.n1632 vp_n.n1631 0.319
R56223 vp_n.n1642 vp_n.n1641 0.319
R56224 vp_n.n1652 vp_n.n1651 0.319
R56225 vp_n.n1662 vp_n.n1661 0.319
R56226 vp_n.n1672 vp_n.n1671 0.319
R56227 vp_n.n1682 vp_n.n1681 0.319
R56228 vp_n.n1692 vp_n.n1691 0.319
R56229 vp_n.n1702 vp_n.n1701 0.319
R56230 vp_n.n1712 vp_n.n1711 0.319
R56231 vp_n.n1722 vp_n.n1721 0.319
R56232 vp_n.n1732 vp_n.n1731 0.319
R56233 vp_n.n1742 vp_n.n1741 0.319
R56234 vp_n.n1752 vp_n.n1751 0.319
R56235 vp_n.n1762 vp_n.n1761 0.319
R56236 vp_n.n1772 vp_n.n1771 0.319
R56237 vp_n.n1782 vp_n.n1781 0.319
R56238 vp_n.n1792 vp_n.n1791 0.319
R56239 vp_n.n1802 vp_n.n1801 0.319
R56240 vp_n.n1812 vp_n.n1811 0.319
R56241 vp_n.n1822 vp_n.n1821 0.319
R56242 vp_n.n1832 vp_n.n1831 0.319
R56243 vp_n.n1842 vp_n.n1841 0.319
R56244 vp_n.n1852 vp_n.n1851 0.319
R56245 vp_n.n1862 vp_n.n1861 0.319
R56246 vp_n.n1872 vp_n.n1871 0.319
R56247 vp_n.n1882 vp_n.n1881 0.319
R56248 vp_n.n1892 vp_n.n1891 0.319
R56249 vp_n.n1902 vp_n.n1901 0.319
R56250 vp_n.n1912 vp_n.n1911 0.319
R56251 vp_n.n1922 vp_n.n1921 0.319
R56252 vp_n.n1932 vp_n.n1931 0.319
R56253 vp_n.n1942 vp_n.n1941 0.319
R56254 vp_n.n1952 vp_n.n1951 0.319
R56255 vp_n.n1962 vp_n.n1961 0.319
R56256 vp_n.n1972 vp_n.n1971 0.319
R56257 vp_n.n1982 vp_n.n1981 0.319
R56258 vp_n.n1992 vp_n.n1991 0.319
R56259 vp_n.n2002 vp_n.n2001 0.319
R56260 vp_n.n2012 vp_n.n2011 0.319
R56261 vp_n.n2022 vp_n.n2021 0.319
R56262 vp_n.n2032 vp_n.n2031 0.319
R56263 vp_n.n2042 vp_n.n2041 0.319
R56264 vp_n.n2052 vp_n.n2051 0.319
R56265 vp_n.n2062 vp_n.n2061 0.319
R56266 vp_n.n2072 vp_n.n2071 0.319
R56267 vp_n.n2082 vp_n.n2081 0.319
R56268 vp_n.n2092 vp_n.n2091 0.319
R56269 vp_n.n2102 vp_n.n2101 0.319
R56270 vp_n.n2112 vp_n.n2111 0.319
R56271 vp_n.n2122 vp_n.n2121 0.319
R56272 vp_n.n2132 vp_n.n2131 0.319
R56273 vp_n.n2142 vp_n.n2141 0.319
R56274 vp_n.n2152 vp_n.n2151 0.319
R56275 vp_n.n2162 vp_n.n2161 0.319
R56276 vp_n.n2172 vp_n.n2171 0.319
R56277 vp_n.n2182 vp_n.n2181 0.319
R56278 vp_n.n2192 vp_n.n2191 0.319
R56279 vp_n.n2202 vp_n.n2201 0.319
R56280 vp_n.n2212 vp_n.n2211 0.319
R56281 vp_n.n2222 vp_n.n2221 0.319
R56282 vp_n.n2232 vp_n.n2231 0.319
R56283 vp_n.n2242 vp_n.n2241 0.319
R56284 vp_n.n2252 vp_n.n2251 0.319
R56285 vp_n.n2262 vp_n.n2261 0.319
R56286 vp_n.n2272 vp_n.n2271 0.319
R56287 vp_n.n2282 vp_n.n2281 0.319
R56288 vp_n.n2292 vp_n.n2291 0.319
R56289 vp_n.n2302 vp_n.n2301 0.319
R56290 vp_n.n2312 vp_n.n2311 0.319
R56291 vp_n.n2322 vp_n.n2321 0.319
R56292 vp_n.n2332 vp_n.n2331 0.319
R56293 vp_n.n2342 vp_n.n2341 0.319
R56294 vp_n.n2352 vp_n.n2351 0.319
R56295 vp_n.n2362 vp_n.n2361 0.319
R56296 vp_n.n2372 vp_n.n2371 0.319
R56297 vp_n.n2382 vp_n.n2381 0.319
R56298 vp_n.n2392 vp_n.n2391 0.319
R56299 vp_n.n2402 vp_n.n2401 0.319
R56300 vp_n.n2412 vp_n.n2411 0.319
R56301 vp_n.n2422 vp_n.n2421 0.319
R56302 vp_n.n2432 vp_n.n2431 0.319
R56303 vp_n.n2442 vp_n.n2441 0.319
R56304 vp_n.n2452 vp_n.n2451 0.319
R56305 vp_n.n2462 vp_n.n2461 0.319
R56306 vp_n.n2472 vp_n.n2471 0.319
R56307 vp_n.n2482 vp_n.n2481 0.319
R56308 vp_n.n2492 vp_n.n2491 0.319
R56309 vp_n.n2502 vp_n.n2501 0.319
R56310 vp_n.n2512 vp_n.n2511 0.319
R56311 vp_n.n2522 vp_n.n2521 0.319
R56312 vp_n.n2532 vp_n.n2531 0.319
R56313 vp_n.n2542 vp_n.n2541 0.319
R56314 vp_n.n2552 vp_n.n2551 0.319
R56315 vp_n.n2562 vp_n.n2561 0.319
R56316 vp_n.n2572 vp_n.n2571 0.319
R56317 vp_n.n2582 vp_n.n2581 0.319
R56318 vp_n.n2592 vp_n.n2591 0.319
R56319 vp_n.n2602 vp_n.n2601 0.319
R56320 vp_n.n2612 vp_n.n2611 0.319
R56321 vp_n.n2622 vp_n.n2621 0.319
R56322 vp_n.n2632 vp_n.n2631 0.319
R56323 vp_n.n2642 vp_n.n2641 0.319
R56324 vp_n.n2652 vp_n.n2651 0.319
R56325 vp_n.n2662 vp_n.n2661 0.319
R56326 vp_n.n2672 vp_n.n2671 0.319
R56327 vp_n.n2682 vp_n.n2681 0.319
R56328 vp_n.n2692 vp_n.n2691 0.319
R56329 vp_n.n2702 vp_n.n2701 0.319
R56330 vp_n.n2712 vp_n.n2711 0.319
R56331 vp_n.n2722 vp_n.n2721 0.319
R56332 vp_n.n2732 vp_n.n2731 0.319
R56333 vp_n.n2742 vp_n.n2741 0.319
R56334 vp_n.n2752 vp_n.n2751 0.319
R56335 vp_n.n2762 vp_n.n2761 0.319
R56336 vp_n.n2772 vp_n.n2771 0.319
R56337 vp_n.n2782 vp_n.n2781 0.319
R56338 vp_n.n2792 vp_n.n2791 0.319
R56339 vp_n.n2802 vp_n.n2801 0.319
R56340 vp_n.n2812 vp_n.n2811 0.319
R56341 vp_n.n2822 vp_n.n2821 0.319
R56342 vp_n.n2832 vp_n.n2831 0.319
R56343 vp_n.n2842 vp_n.n2841 0.319
R56344 vp_n.n2852 vp_n.n2851 0.319
R56345 vp_n.n2862 vp_n.n2861 0.319
R56346 vp_n.n2872 vp_n.n2871 0.319
R56347 vp_n.n2882 vp_n.n2881 0.319
R56348 vp_n.n2892 vp_n.n2891 0.319
R56349 vp_n.n2902 vp_n.n2901 0.319
R56350 vp_n.n2912 vp_n.n2911 0.319
R56351 vp_n.n2922 vp_n.n2921 0.319
R56352 vp_n.n2932 vp_n.n2931 0.319
R56353 vp_n.n2942 vp_n.n2941 0.319
R56354 vp_n.n2952 vp_n.n2951 0.319
R56355 vp_n.n2962 vp_n.n2961 0.319
R56356 vp_n.n2972 vp_n.n2971 0.319
R56357 vp_n.n2982 vp_n.n2981 0.319
R56358 vp_n.n2992 vp_n.n2991 0.319
R56359 vp_n.n3002 vp_n.n3001 0.319
R56360 vp_n.n3012 vp_n.n3011 0.319
R56361 vp_n.n3022 vp_n.n3021 0.319
R56362 vp_n.n3032 vp_n.n3031 0.319
R56363 vp_n.n3042 vp_n.n3041 0.319
R56364 vp_n.n3215 vp_n.n3214 0.319
R56365 vp_n.n3225 vp_n.n3224 0.319
R56366 vp_n.n3235 vp_n.n3234 0.319
R56367 vp_n.n3245 vp_n.n3244 0.319
R56368 vp_n.n3255 vp_n.n3254 0.319
R56369 vp_n.n3265 vp_n.n3264 0.319
R56370 vp_n.n3275 vp_n.n3274 0.319
R56371 vp_n.n3285 vp_n.n3284 0.319
R56372 vp_n.n3295 vp_n.n3294 0.319
R56373 vp_n.n3305 vp_n.n3304 0.319
R56374 vp_n.n3315 vp_n.n3314 0.319
R56375 vp_n.n3325 vp_n.n3324 0.319
R56376 vp_n.n3335 vp_n.n3334 0.319
R56377 vp_n.n3345 vp_n.n3344 0.319
R56378 vp_n.n3355 vp_n.n3354 0.319
R56379 vp_n.n3365 vp_n.n3364 0.319
R56380 vp_n.n3375 vp_n.n3374 0.319
R56381 vp_n.n3385 vp_n.n3384 0.319
R56382 vp_n.n3395 vp_n.n3394 0.319
R56383 vp_n.n3405 vp_n.n3404 0.319
R56384 vp_n.n3415 vp_n.n3414 0.319
R56385 vp_n.n3425 vp_n.n3424 0.319
R56386 vp_n.n3435 vp_n.n3434 0.319
R56387 vp_n.n3445 vp_n.n3444 0.319
R56388 vp_n.n3455 vp_n.n3454 0.319
R56389 vp_n.n3465 vp_n.n3464 0.319
R56390 vp_n.n3475 vp_n.n3474 0.319
R56391 vp_n.n3485 vp_n.n3484 0.319
R56392 vp_n.n3495 vp_n.n3494 0.319
R56393 vp_n.n3505 vp_n.n3504 0.319
R56394 vp_n.n3515 vp_n.n3514 0.319
R56395 vp_n.n3525 vp_n.n3524 0.319
R56396 vp_n.n3535 vp_n.n3534 0.319
R56397 vp_n.n3545 vp_n.n3544 0.319
R56398 vp_n.n3555 vp_n.n3554 0.319
R56399 vp_n.n3565 vp_n.n3564 0.319
R56400 vp_n.n3575 vp_n.n3574 0.319
R56401 vp_n.n3585 vp_n.n3584 0.319
R56402 vp_n.n3595 vp_n.n3594 0.319
R56403 vp_n.n3605 vp_n.n3604 0.319
R56404 vp_n.n3615 vp_n.n3614 0.319
R56405 vp_n.n3625 vp_n.n3624 0.319
R56406 vp_n.n3635 vp_n.n3634 0.319
R56407 vp_n.n3645 vp_n.n3644 0.319
R56408 vp_n.n3655 vp_n.n3654 0.319
R56409 vp_n.n3665 vp_n.n3664 0.319
R56410 vp_n.n3675 vp_n.n3674 0.319
R56411 vp_n.n3685 vp_n.n3684 0.319
R56412 vp_n.n3695 vp_n.n3694 0.319
R56413 vp_n.n3705 vp_n.n3704 0.319
R56414 vp_n.n3715 vp_n.n3714 0.319
R56415 vp_n.n3725 vp_n.n3724 0.319
R56416 vp_n.n3735 vp_n.n3734 0.319
R56417 vp_n.n3745 vp_n.n3744 0.319
R56418 vp_n.n3755 vp_n.n3754 0.319
R56419 vp_n.n3765 vp_n.n3764 0.319
R56420 vp_n.n3775 vp_n.n3774 0.319
R56421 vp_n.n3785 vp_n.n3784 0.319
R56422 vp_n.n3795 vp_n.n3794 0.319
R56423 vp_n.n3805 vp_n.n3804 0.319
R56424 vp_n.n3815 vp_n.n3814 0.319
R56425 vp_n.n3825 vp_n.n3824 0.319
R56426 vp_n.n3835 vp_n.n3834 0.319
R56427 vp_n.n3845 vp_n.n3844 0.319
R56428 vp_n.n3855 vp_n.n3854 0.319
R56429 vp_n.n3865 vp_n.n3864 0.319
R56430 vp_n.n3875 vp_n.n3874 0.319
R56431 vp_n.n3885 vp_n.n3884 0.319
R56432 vp_n.n3895 vp_n.n3894 0.319
R56433 vp_n.n3905 vp_n.n3904 0.319
R56434 vp_n.n3915 vp_n.n3914 0.319
R56435 vp_n.n3925 vp_n.n3924 0.319
R56436 vp_n.n3935 vp_n.n3934 0.319
R56437 vp_n.n3945 vp_n.n3944 0.319
R56438 vp_n.n3955 vp_n.n3954 0.319
R56439 vp_n.n3965 vp_n.n3964 0.319
R56440 vp_n.n3975 vp_n.n3974 0.319
R56441 vp_n.n3985 vp_n.n3984 0.319
R56442 vp_n.n3995 vp_n.n3994 0.319
R56443 vp_n.n4005 vp_n.n4004 0.319
R56444 vp_n.n4015 vp_n.n4014 0.319
R56445 vp_n.n4025 vp_n.n4024 0.319
R56446 vp_n.n4035 vp_n.n4034 0.319
R56447 vp_n.n4045 vp_n.n4044 0.319
R56448 vp_n.n4055 vp_n.n4054 0.319
R56449 vp_n.n4065 vp_n.n4064 0.319
R56450 vp_n.n4075 vp_n.n4074 0.319
R56451 vp_n.n4085 vp_n.n4084 0.319
R56452 vp_n.n4095 vp_n.n4094 0.319
R56453 vp_n.n4105 vp_n.n4104 0.319
R56454 vp_n.n4115 vp_n.n4114 0.319
R56455 vp_n.n4125 vp_n.n4124 0.319
R56456 vp_n.n4135 vp_n.n4134 0.319
R56457 vp_n.n4145 vp_n.n4144 0.319
R56458 vp_n.n4155 vp_n.n4154 0.319
R56459 vp_n.n4165 vp_n.n4164 0.319
R56460 vp_n.n4175 vp_n.n4174 0.319
R56461 vp_n.n4185 vp_n.n4184 0.319
R56462 vp_n.n4195 vp_n.n4194 0.319
R56463 vp_n.n4205 vp_n.n4204 0.319
R56464 vp_n.n4215 vp_n.n4214 0.319
R56465 vp_n.n4225 vp_n.n4224 0.319
R56466 vp_n.n4235 vp_n.n4234 0.319
R56467 vp_n.n4245 vp_n.n4244 0.319
R56468 vp_n.n4255 vp_n.n4254 0.319
R56469 vp_n.n4265 vp_n.n4264 0.319
R56470 vp_n.n4275 vp_n.n4274 0.319
R56471 vp_n.n4285 vp_n.n4284 0.319
R56472 vp_n.n4295 vp_n.n4294 0.319
R56473 vp_n.n4305 vp_n.n4304 0.319
R56474 vp_n.n4315 vp_n.n4314 0.319
R56475 vp_n.n4325 vp_n.n4324 0.319
R56476 vp_n.n4335 vp_n.n4334 0.319
R56477 vp_n.n4345 vp_n.n4344 0.319
R56478 vp_n.n4355 vp_n.n4354 0.319
R56479 vp_n.n4365 vp_n.n4364 0.319
R56480 vp_n.n4375 vp_n.n4374 0.319
R56481 vp_n.n4385 vp_n.n4384 0.319
R56482 vp_n.n4395 vp_n.n4394 0.319
R56483 vp_n.n4405 vp_n.n4404 0.319
R56484 vp_n.n4415 vp_n.n4414 0.319
R56485 vp_n.n4425 vp_n.n4424 0.319
R56486 vp_n.n4435 vp_n.n4434 0.319
R56487 vp_n.n4445 vp_n.n4444 0.319
R56488 vp_n.n4455 vp_n.n4454 0.319
R56489 vp_n.n4465 vp_n.n4464 0.319
R56490 vp_n.n4475 vp_n.n4474 0.319
R56491 vp_n.n4485 vp_n.n4484 0.319
R56492 vp_n.n4495 vp_n.n4494 0.319
R56493 vp_n.n4505 vp_n.n4504 0.319
R56494 vp_n.n4515 vp_n.n4514 0.319
R56495 vp_n.n4525 vp_n.n4524 0.319
R56496 vp_n.n4535 vp_n.n4534 0.319
R56497 vp_n.n4545 vp_n.n4544 0.319
R56498 vp_n.n4555 vp_n.n4554 0.319
R56499 vp_n.n4565 vp_n.n4564 0.319
R56500 vp_n.n4575 vp_n.n4574 0.319
R56501 vp_n.n4585 vp_n.n4584 0.319
R56502 vp_n.n4595 vp_n.n4594 0.319
R56503 vp_n.n4605 vp_n.n4604 0.319
R56504 vp_n.n4615 vp_n.n4614 0.319
R56505 vp_n.n4625 vp_n.n4624 0.319
R56506 vp_n.n4635 vp_n.n4634 0.319
R56507 vp_n.n4645 vp_n.n4644 0.319
R56508 vp_n.n4655 vp_n.n4654 0.319
R56509 vp_n.n4665 vp_n.n4664 0.319
R56510 vp_n.n4675 vp_n.n4674 0.319
R56511 vp_n.n4685 vp_n.n4684 0.319
R56512 vp_n.n4695 vp_n.n4694 0.319
R56513 vp_n.n3153 vp_n.n3152 0.179
R56514 vp_n vp_n.n3153 0.104
R56515 vp_n vp_n.n4805 0.075
R56516 vp_n.n10 vp_n.n9 0.014
R56517 vp_n.n20 vp_n.n19 0.014
R56518 vp_n.n30 vp_n.n29 0.014
R56519 vp_n.n40 vp_n.n39 0.014
R56520 vp_n.n50 vp_n.n49 0.014
R56521 vp_n.n60 vp_n.n59 0.014
R56522 vp_n.n70 vp_n.n69 0.014
R56523 vp_n.n80 vp_n.n79 0.014
R56524 vp_n.n90 vp_n.n89 0.014
R56525 vp_n.n100 vp_n.n99 0.014
R56526 vp_n.n110 vp_n.n109 0.014
R56527 vp_n.n120 vp_n.n119 0.014
R56528 vp_n.n130 vp_n.n129 0.014
R56529 vp_n.n140 vp_n.n139 0.014
R56530 vp_n.n150 vp_n.n149 0.014
R56531 vp_n.n160 vp_n.n159 0.014
R56532 vp_n.n170 vp_n.n169 0.014
R56533 vp_n.n180 vp_n.n179 0.014
R56534 vp_n.n190 vp_n.n189 0.014
R56535 vp_n.n200 vp_n.n199 0.014
R56536 vp_n.n210 vp_n.n209 0.014
R56537 vp_n.n220 vp_n.n219 0.014
R56538 vp_n.n230 vp_n.n229 0.014
R56539 vp_n.n240 vp_n.n239 0.014
R56540 vp_n.n250 vp_n.n249 0.014
R56541 vp_n.n260 vp_n.n259 0.014
R56542 vp_n.n270 vp_n.n269 0.014
R56543 vp_n.n280 vp_n.n279 0.014
R56544 vp_n.n290 vp_n.n289 0.014
R56545 vp_n.n300 vp_n.n299 0.014
R56546 vp_n.n310 vp_n.n309 0.014
R56547 vp_n.n320 vp_n.n319 0.014
R56548 vp_n.n330 vp_n.n329 0.014
R56549 vp_n.n340 vp_n.n339 0.014
R56550 vp_n.n350 vp_n.n349 0.014
R56551 vp_n.n360 vp_n.n359 0.014
R56552 vp_n.n370 vp_n.n369 0.014
R56553 vp_n.n380 vp_n.n379 0.014
R56554 vp_n.n390 vp_n.n389 0.014
R56555 vp_n.n400 vp_n.n399 0.014
R56556 vp_n.n410 vp_n.n409 0.014
R56557 vp_n.n420 vp_n.n419 0.014
R56558 vp_n.n430 vp_n.n429 0.014
R56559 vp_n.n440 vp_n.n439 0.014
R56560 vp_n.n450 vp_n.n449 0.014
R56561 vp_n.n460 vp_n.n459 0.014
R56562 vp_n.n470 vp_n.n469 0.014
R56563 vp_n.n480 vp_n.n479 0.014
R56564 vp_n.n490 vp_n.n489 0.014
R56565 vp_n.n500 vp_n.n499 0.014
R56566 vp_n.n510 vp_n.n509 0.014
R56567 vp_n.n520 vp_n.n519 0.014
R56568 vp_n.n530 vp_n.n529 0.014
R56569 vp_n.n540 vp_n.n539 0.014
R56570 vp_n.n550 vp_n.n549 0.014
R56571 vp_n.n560 vp_n.n559 0.014
R56572 vp_n.n570 vp_n.n569 0.014
R56573 vp_n.n580 vp_n.n579 0.014
R56574 vp_n.n590 vp_n.n589 0.014
R56575 vp_n.n600 vp_n.n599 0.014
R56576 vp_n.n610 vp_n.n609 0.014
R56577 vp_n.n620 vp_n.n619 0.014
R56578 vp_n.n630 vp_n.n629 0.014
R56579 vp_n.n640 vp_n.n639 0.014
R56580 vp_n.n650 vp_n.n649 0.014
R56581 vp_n.n660 vp_n.n659 0.014
R56582 vp_n.n670 vp_n.n669 0.014
R56583 vp_n.n680 vp_n.n679 0.014
R56584 vp_n.n690 vp_n.n689 0.014
R56585 vp_n.n700 vp_n.n699 0.014
R56586 vp_n.n710 vp_n.n709 0.014
R56587 vp_n.n720 vp_n.n719 0.014
R56588 vp_n.n730 vp_n.n729 0.014
R56589 vp_n.n740 vp_n.n739 0.014
R56590 vp_n.n750 vp_n.n749 0.014
R56591 vp_n.n760 vp_n.n759 0.014
R56592 vp_n.n770 vp_n.n769 0.014
R56593 vp_n.n780 vp_n.n779 0.014
R56594 vp_n.n790 vp_n.n789 0.014
R56595 vp_n.n800 vp_n.n799 0.014
R56596 vp_n.n810 vp_n.n809 0.014
R56597 vp_n.n820 vp_n.n819 0.014
R56598 vp_n.n830 vp_n.n829 0.014
R56599 vp_n.n840 vp_n.n839 0.014
R56600 vp_n.n850 vp_n.n849 0.014
R56601 vp_n.n860 vp_n.n859 0.014
R56602 vp_n.n870 vp_n.n869 0.014
R56603 vp_n.n880 vp_n.n879 0.014
R56604 vp_n.n890 vp_n.n889 0.014
R56605 vp_n.n900 vp_n.n899 0.014
R56606 vp_n.n910 vp_n.n909 0.014
R56607 vp_n.n920 vp_n.n919 0.014
R56608 vp_n.n930 vp_n.n929 0.014
R56609 vp_n.n940 vp_n.n939 0.014
R56610 vp_n.n950 vp_n.n949 0.014
R56611 vp_n.n960 vp_n.n959 0.014
R56612 vp_n.n970 vp_n.n969 0.014
R56613 vp_n.n980 vp_n.n979 0.014
R56614 vp_n.n990 vp_n.n989 0.014
R56615 vp_n.n1000 vp_n.n999 0.014
R56616 vp_n.n1010 vp_n.n1009 0.014
R56617 vp_n.n1020 vp_n.n1019 0.014
R56618 vp_n.n1030 vp_n.n1029 0.014
R56619 vp_n.n1040 vp_n.n1039 0.014
R56620 vp_n.n1050 vp_n.n1049 0.014
R56621 vp_n.n1060 vp_n.n1059 0.014
R56622 vp_n.n1070 vp_n.n1069 0.014
R56623 vp_n.n1080 vp_n.n1079 0.014
R56624 vp_n.n1090 vp_n.n1089 0.014
R56625 vp_n.n1100 vp_n.n1099 0.014
R56626 vp_n.n1110 vp_n.n1109 0.014
R56627 vp_n.n1120 vp_n.n1119 0.014
R56628 vp_n.n1130 vp_n.n1129 0.014
R56629 vp_n.n1140 vp_n.n1139 0.014
R56630 vp_n.n1150 vp_n.n1149 0.014
R56631 vp_n.n1160 vp_n.n1159 0.014
R56632 vp_n.n1170 vp_n.n1169 0.014
R56633 vp_n.n1180 vp_n.n1179 0.014
R56634 vp_n.n1190 vp_n.n1189 0.014
R56635 vp_n.n1200 vp_n.n1199 0.014
R56636 vp_n.n1210 vp_n.n1209 0.014
R56637 vp_n.n1220 vp_n.n1219 0.014
R56638 vp_n.n1230 vp_n.n1229 0.014
R56639 vp_n.n1240 vp_n.n1239 0.014
R56640 vp_n.n1250 vp_n.n1249 0.014
R56641 vp_n.n1260 vp_n.n1259 0.014
R56642 vp_n.n1270 vp_n.n1269 0.014
R56643 vp_n.n1280 vp_n.n1279 0.014
R56644 vp_n.n1290 vp_n.n1289 0.014
R56645 vp_n.n1300 vp_n.n1299 0.014
R56646 vp_n.n1310 vp_n.n1309 0.014
R56647 vp_n.n1320 vp_n.n1319 0.014
R56648 vp_n.n1330 vp_n.n1329 0.014
R56649 vp_n.n1340 vp_n.n1339 0.014
R56650 vp_n.n1350 vp_n.n1349 0.014
R56651 vp_n.n1360 vp_n.n1359 0.014
R56652 vp_n.n1370 vp_n.n1369 0.014
R56653 vp_n.n1380 vp_n.n1379 0.014
R56654 vp_n.n1390 vp_n.n1389 0.014
R56655 vp_n.n1400 vp_n.n1399 0.014
R56656 vp_n.n1410 vp_n.n1409 0.014
R56657 vp_n.n1420 vp_n.n1419 0.014
R56658 vp_n.n1430 vp_n.n1429 0.014
R56659 vp_n.n1440 vp_n.n1439 0.014
R56660 vp_n.n1450 vp_n.n1449 0.014
R56661 vp_n.n1460 vp_n.n1459 0.014
R56662 vp_n.n1470 vp_n.n1469 0.014
R56663 vp_n.n1480 vp_n.n1479 0.014
R56664 vp_n.n1490 vp_n.n1489 0.014
R56665 vp_n.n1500 vp_n.n1499 0.014
R56666 vp_n.n1561 vp_n.n1560 0.014
R56667 vp_n.n1571 vp_n.n1570 0.014
R56668 vp_n.n1581 vp_n.n1580 0.014
R56669 vp_n.n1591 vp_n.n1590 0.014
R56670 vp_n.n1601 vp_n.n1600 0.014
R56671 vp_n.n1611 vp_n.n1610 0.014
R56672 vp_n.n1621 vp_n.n1620 0.014
R56673 vp_n.n1631 vp_n.n1630 0.014
R56674 vp_n.n1641 vp_n.n1640 0.014
R56675 vp_n.n1651 vp_n.n1650 0.014
R56676 vp_n.n1661 vp_n.n1660 0.014
R56677 vp_n.n1671 vp_n.n1670 0.014
R56678 vp_n.n1681 vp_n.n1680 0.014
R56679 vp_n.n1691 vp_n.n1690 0.014
R56680 vp_n.n1701 vp_n.n1700 0.014
R56681 vp_n.n1711 vp_n.n1710 0.014
R56682 vp_n.n1721 vp_n.n1720 0.014
R56683 vp_n.n1731 vp_n.n1730 0.014
R56684 vp_n.n1741 vp_n.n1740 0.014
R56685 vp_n.n1751 vp_n.n1750 0.014
R56686 vp_n.n1761 vp_n.n1760 0.014
R56687 vp_n.n1771 vp_n.n1770 0.014
R56688 vp_n.n1781 vp_n.n1780 0.014
R56689 vp_n.n1791 vp_n.n1790 0.014
R56690 vp_n.n1801 vp_n.n1800 0.014
R56691 vp_n.n1811 vp_n.n1810 0.014
R56692 vp_n.n1821 vp_n.n1820 0.014
R56693 vp_n.n1831 vp_n.n1830 0.014
R56694 vp_n.n1841 vp_n.n1840 0.014
R56695 vp_n.n1851 vp_n.n1850 0.014
R56696 vp_n.n1861 vp_n.n1860 0.014
R56697 vp_n.n1871 vp_n.n1870 0.014
R56698 vp_n.n1881 vp_n.n1880 0.014
R56699 vp_n.n1891 vp_n.n1890 0.014
R56700 vp_n.n1901 vp_n.n1900 0.014
R56701 vp_n.n1911 vp_n.n1910 0.014
R56702 vp_n.n1921 vp_n.n1920 0.014
R56703 vp_n.n1931 vp_n.n1930 0.014
R56704 vp_n.n1941 vp_n.n1940 0.014
R56705 vp_n.n1951 vp_n.n1950 0.014
R56706 vp_n.n1961 vp_n.n1960 0.014
R56707 vp_n.n1971 vp_n.n1970 0.014
R56708 vp_n.n1981 vp_n.n1980 0.014
R56709 vp_n.n1991 vp_n.n1990 0.014
R56710 vp_n.n2001 vp_n.n2000 0.014
R56711 vp_n.n2011 vp_n.n2010 0.014
R56712 vp_n.n2021 vp_n.n2020 0.014
R56713 vp_n.n2031 vp_n.n2030 0.014
R56714 vp_n.n2041 vp_n.n2040 0.014
R56715 vp_n.n2051 vp_n.n2050 0.014
R56716 vp_n.n2061 vp_n.n2060 0.014
R56717 vp_n.n2071 vp_n.n2070 0.014
R56718 vp_n.n2081 vp_n.n2080 0.014
R56719 vp_n.n2091 vp_n.n2090 0.014
R56720 vp_n.n2101 vp_n.n2100 0.014
R56721 vp_n.n2111 vp_n.n2110 0.014
R56722 vp_n.n2121 vp_n.n2120 0.014
R56723 vp_n.n2131 vp_n.n2130 0.014
R56724 vp_n.n2141 vp_n.n2140 0.014
R56725 vp_n.n2151 vp_n.n2150 0.014
R56726 vp_n.n2161 vp_n.n2160 0.014
R56727 vp_n.n2171 vp_n.n2170 0.014
R56728 vp_n.n2181 vp_n.n2180 0.014
R56729 vp_n.n2191 vp_n.n2190 0.014
R56730 vp_n.n2201 vp_n.n2200 0.014
R56731 vp_n.n2211 vp_n.n2210 0.014
R56732 vp_n.n2221 vp_n.n2220 0.014
R56733 vp_n.n2231 vp_n.n2230 0.014
R56734 vp_n.n2241 vp_n.n2240 0.014
R56735 vp_n.n2251 vp_n.n2250 0.014
R56736 vp_n.n2261 vp_n.n2260 0.014
R56737 vp_n.n2271 vp_n.n2270 0.014
R56738 vp_n.n2281 vp_n.n2280 0.014
R56739 vp_n.n2291 vp_n.n2290 0.014
R56740 vp_n.n2301 vp_n.n2300 0.014
R56741 vp_n.n2311 vp_n.n2310 0.014
R56742 vp_n.n2321 vp_n.n2320 0.014
R56743 vp_n.n2331 vp_n.n2330 0.014
R56744 vp_n.n2341 vp_n.n2340 0.014
R56745 vp_n.n2351 vp_n.n2350 0.014
R56746 vp_n.n2361 vp_n.n2360 0.014
R56747 vp_n.n2371 vp_n.n2370 0.014
R56748 vp_n.n2381 vp_n.n2380 0.014
R56749 vp_n.n2391 vp_n.n2390 0.014
R56750 vp_n.n2401 vp_n.n2400 0.014
R56751 vp_n.n2411 vp_n.n2410 0.014
R56752 vp_n.n2421 vp_n.n2420 0.014
R56753 vp_n.n2431 vp_n.n2430 0.014
R56754 vp_n.n2441 vp_n.n2440 0.014
R56755 vp_n.n2451 vp_n.n2450 0.014
R56756 vp_n.n2461 vp_n.n2460 0.014
R56757 vp_n.n2471 vp_n.n2470 0.014
R56758 vp_n.n2481 vp_n.n2480 0.014
R56759 vp_n.n2491 vp_n.n2490 0.014
R56760 vp_n.n2501 vp_n.n2500 0.014
R56761 vp_n.n2511 vp_n.n2510 0.014
R56762 vp_n.n2521 vp_n.n2520 0.014
R56763 vp_n.n2531 vp_n.n2530 0.014
R56764 vp_n.n2541 vp_n.n2540 0.014
R56765 vp_n.n2551 vp_n.n2550 0.014
R56766 vp_n.n2561 vp_n.n2560 0.014
R56767 vp_n.n2571 vp_n.n2570 0.014
R56768 vp_n.n2581 vp_n.n2580 0.014
R56769 vp_n.n2591 vp_n.n2590 0.014
R56770 vp_n.n2601 vp_n.n2600 0.014
R56771 vp_n.n2611 vp_n.n2610 0.014
R56772 vp_n.n2621 vp_n.n2620 0.014
R56773 vp_n.n2631 vp_n.n2630 0.014
R56774 vp_n.n2641 vp_n.n2640 0.014
R56775 vp_n.n2651 vp_n.n2650 0.014
R56776 vp_n.n2661 vp_n.n2660 0.014
R56777 vp_n.n2671 vp_n.n2670 0.014
R56778 vp_n.n2681 vp_n.n2680 0.014
R56779 vp_n.n2691 vp_n.n2690 0.014
R56780 vp_n.n2701 vp_n.n2700 0.014
R56781 vp_n.n2711 vp_n.n2710 0.014
R56782 vp_n.n2721 vp_n.n2720 0.014
R56783 vp_n.n2731 vp_n.n2730 0.014
R56784 vp_n.n2741 vp_n.n2740 0.014
R56785 vp_n.n2751 vp_n.n2750 0.014
R56786 vp_n.n2761 vp_n.n2760 0.014
R56787 vp_n.n2771 vp_n.n2770 0.014
R56788 vp_n.n2781 vp_n.n2780 0.014
R56789 vp_n.n2791 vp_n.n2790 0.014
R56790 vp_n.n2801 vp_n.n2800 0.014
R56791 vp_n.n2811 vp_n.n2810 0.014
R56792 vp_n.n2821 vp_n.n2820 0.014
R56793 vp_n.n2831 vp_n.n2830 0.014
R56794 vp_n.n2841 vp_n.n2840 0.014
R56795 vp_n.n2851 vp_n.n2850 0.014
R56796 vp_n.n2861 vp_n.n2860 0.014
R56797 vp_n.n2871 vp_n.n2870 0.014
R56798 vp_n.n2881 vp_n.n2880 0.014
R56799 vp_n.n2891 vp_n.n2890 0.014
R56800 vp_n.n2901 vp_n.n2900 0.014
R56801 vp_n.n2911 vp_n.n2910 0.014
R56802 vp_n.n2921 vp_n.n2920 0.014
R56803 vp_n.n2931 vp_n.n2930 0.014
R56804 vp_n.n2941 vp_n.n2940 0.014
R56805 vp_n.n2951 vp_n.n2950 0.014
R56806 vp_n.n2961 vp_n.n2960 0.014
R56807 vp_n.n2971 vp_n.n2970 0.014
R56808 vp_n.n2981 vp_n.n2980 0.014
R56809 vp_n.n2991 vp_n.n2990 0.014
R56810 vp_n.n3001 vp_n.n3000 0.014
R56811 vp_n.n3011 vp_n.n3010 0.014
R56812 vp_n.n3021 vp_n.n3020 0.014
R56813 vp_n.n3031 vp_n.n3030 0.014
R56814 vp_n.n3041 vp_n.n3040 0.014
R56815 vp_n.n3051 vp_n.n3050 0.014
R56816 vp_n.n3214 vp_n.n3213 0.014
R56817 vp_n.n3224 vp_n.n3223 0.014
R56818 vp_n.n3234 vp_n.n3233 0.014
R56819 vp_n.n3244 vp_n.n3243 0.014
R56820 vp_n.n3254 vp_n.n3253 0.014
R56821 vp_n.n3264 vp_n.n3263 0.014
R56822 vp_n.n3274 vp_n.n3273 0.014
R56823 vp_n.n3284 vp_n.n3283 0.014
R56824 vp_n.n3294 vp_n.n3293 0.014
R56825 vp_n.n3304 vp_n.n3303 0.014
R56826 vp_n.n3314 vp_n.n3313 0.014
R56827 vp_n.n3324 vp_n.n3323 0.014
R56828 vp_n.n3334 vp_n.n3333 0.014
R56829 vp_n.n3344 vp_n.n3343 0.014
R56830 vp_n.n3354 vp_n.n3353 0.014
R56831 vp_n.n3364 vp_n.n3363 0.014
R56832 vp_n.n3374 vp_n.n3373 0.014
R56833 vp_n.n3384 vp_n.n3383 0.014
R56834 vp_n.n3394 vp_n.n3393 0.014
R56835 vp_n.n3404 vp_n.n3403 0.014
R56836 vp_n.n3414 vp_n.n3413 0.014
R56837 vp_n.n3424 vp_n.n3423 0.014
R56838 vp_n.n3434 vp_n.n3433 0.014
R56839 vp_n.n3444 vp_n.n3443 0.014
R56840 vp_n.n3454 vp_n.n3453 0.014
R56841 vp_n.n3464 vp_n.n3463 0.014
R56842 vp_n.n3474 vp_n.n3473 0.014
R56843 vp_n.n3484 vp_n.n3483 0.014
R56844 vp_n.n3494 vp_n.n3493 0.014
R56845 vp_n.n3504 vp_n.n3503 0.014
R56846 vp_n.n3514 vp_n.n3513 0.014
R56847 vp_n.n3524 vp_n.n3523 0.014
R56848 vp_n.n3534 vp_n.n3533 0.014
R56849 vp_n.n3544 vp_n.n3543 0.014
R56850 vp_n.n3554 vp_n.n3553 0.014
R56851 vp_n.n3564 vp_n.n3563 0.014
R56852 vp_n.n3574 vp_n.n3573 0.014
R56853 vp_n.n3584 vp_n.n3583 0.014
R56854 vp_n.n3594 vp_n.n3593 0.014
R56855 vp_n.n3604 vp_n.n3603 0.014
R56856 vp_n.n3614 vp_n.n3613 0.014
R56857 vp_n.n3624 vp_n.n3623 0.014
R56858 vp_n.n3634 vp_n.n3633 0.014
R56859 vp_n.n3644 vp_n.n3643 0.014
R56860 vp_n.n3654 vp_n.n3653 0.014
R56861 vp_n.n3664 vp_n.n3663 0.014
R56862 vp_n.n3674 vp_n.n3673 0.014
R56863 vp_n.n3684 vp_n.n3683 0.014
R56864 vp_n.n3694 vp_n.n3693 0.014
R56865 vp_n.n3704 vp_n.n3703 0.014
R56866 vp_n.n3714 vp_n.n3713 0.014
R56867 vp_n.n3724 vp_n.n3723 0.014
R56868 vp_n.n3734 vp_n.n3733 0.014
R56869 vp_n.n3744 vp_n.n3743 0.014
R56870 vp_n.n3754 vp_n.n3753 0.014
R56871 vp_n.n3764 vp_n.n3763 0.014
R56872 vp_n.n3774 vp_n.n3773 0.014
R56873 vp_n.n3784 vp_n.n3783 0.014
R56874 vp_n.n3794 vp_n.n3793 0.014
R56875 vp_n.n3804 vp_n.n3803 0.014
R56876 vp_n.n3814 vp_n.n3813 0.014
R56877 vp_n.n3824 vp_n.n3823 0.014
R56878 vp_n.n3834 vp_n.n3833 0.014
R56879 vp_n.n3844 vp_n.n3843 0.014
R56880 vp_n.n3854 vp_n.n3853 0.014
R56881 vp_n.n3864 vp_n.n3863 0.014
R56882 vp_n.n3874 vp_n.n3873 0.014
R56883 vp_n.n3884 vp_n.n3883 0.014
R56884 vp_n.n3894 vp_n.n3893 0.014
R56885 vp_n.n3904 vp_n.n3903 0.014
R56886 vp_n.n3914 vp_n.n3913 0.014
R56887 vp_n.n3924 vp_n.n3923 0.014
R56888 vp_n.n3934 vp_n.n3933 0.014
R56889 vp_n.n3944 vp_n.n3943 0.014
R56890 vp_n.n3954 vp_n.n3953 0.014
R56891 vp_n.n3964 vp_n.n3963 0.014
R56892 vp_n.n3974 vp_n.n3973 0.014
R56893 vp_n.n3984 vp_n.n3983 0.014
R56894 vp_n.n3994 vp_n.n3993 0.014
R56895 vp_n.n4004 vp_n.n4003 0.014
R56896 vp_n.n4014 vp_n.n4013 0.014
R56897 vp_n.n4024 vp_n.n4023 0.014
R56898 vp_n.n4034 vp_n.n4033 0.014
R56899 vp_n.n4044 vp_n.n4043 0.014
R56900 vp_n.n4054 vp_n.n4053 0.014
R56901 vp_n.n4064 vp_n.n4063 0.014
R56902 vp_n.n4074 vp_n.n4073 0.014
R56903 vp_n.n4084 vp_n.n4083 0.014
R56904 vp_n.n4094 vp_n.n4093 0.014
R56905 vp_n.n4104 vp_n.n4103 0.014
R56906 vp_n.n4114 vp_n.n4113 0.014
R56907 vp_n.n4124 vp_n.n4123 0.014
R56908 vp_n.n4134 vp_n.n4133 0.014
R56909 vp_n.n4144 vp_n.n4143 0.014
R56910 vp_n.n4154 vp_n.n4153 0.014
R56911 vp_n.n4164 vp_n.n4163 0.014
R56912 vp_n.n4174 vp_n.n4173 0.014
R56913 vp_n.n4184 vp_n.n4183 0.014
R56914 vp_n.n4194 vp_n.n4193 0.014
R56915 vp_n.n4204 vp_n.n4203 0.014
R56916 vp_n.n4214 vp_n.n4213 0.014
R56917 vp_n.n4224 vp_n.n4223 0.014
R56918 vp_n.n4234 vp_n.n4233 0.014
R56919 vp_n.n4244 vp_n.n4243 0.014
R56920 vp_n.n4254 vp_n.n4253 0.014
R56921 vp_n.n4264 vp_n.n4263 0.014
R56922 vp_n.n4274 vp_n.n4273 0.014
R56923 vp_n.n4284 vp_n.n4283 0.014
R56924 vp_n.n4294 vp_n.n4293 0.014
R56925 vp_n.n4304 vp_n.n4303 0.014
R56926 vp_n.n4314 vp_n.n4313 0.014
R56927 vp_n.n4324 vp_n.n4323 0.014
R56928 vp_n.n4334 vp_n.n4333 0.014
R56929 vp_n.n4344 vp_n.n4343 0.014
R56930 vp_n.n4354 vp_n.n4353 0.014
R56931 vp_n.n4364 vp_n.n4363 0.014
R56932 vp_n.n4374 vp_n.n4373 0.014
R56933 vp_n.n4384 vp_n.n4383 0.014
R56934 vp_n.n4394 vp_n.n4393 0.014
R56935 vp_n.n4404 vp_n.n4403 0.014
R56936 vp_n.n4414 vp_n.n4413 0.014
R56937 vp_n.n4424 vp_n.n4423 0.014
R56938 vp_n.n4434 vp_n.n4433 0.014
R56939 vp_n.n4444 vp_n.n4443 0.014
R56940 vp_n.n4454 vp_n.n4453 0.014
R56941 vp_n.n4464 vp_n.n4463 0.014
R56942 vp_n.n4474 vp_n.n4473 0.014
R56943 vp_n.n4484 vp_n.n4483 0.014
R56944 vp_n.n4494 vp_n.n4493 0.014
R56945 vp_n.n4504 vp_n.n4503 0.014
R56946 vp_n.n4514 vp_n.n4513 0.014
R56947 vp_n.n4524 vp_n.n4523 0.014
R56948 vp_n.n4534 vp_n.n4533 0.014
R56949 vp_n.n4544 vp_n.n4543 0.014
R56950 vp_n.n4554 vp_n.n4553 0.014
R56951 vp_n.n4564 vp_n.n4563 0.014
R56952 vp_n.n4574 vp_n.n4573 0.014
R56953 vp_n.n4584 vp_n.n4583 0.014
R56954 vp_n.n4594 vp_n.n4593 0.014
R56955 vp_n.n4604 vp_n.n4603 0.014
R56956 vp_n.n4614 vp_n.n4613 0.014
R56957 vp_n.n4624 vp_n.n4623 0.014
R56958 vp_n.n4634 vp_n.n4633 0.014
R56959 vp_n.n4644 vp_n.n4643 0.014
R56960 vp_n.n4654 vp_n.n4653 0.014
R56961 vp_n.n4664 vp_n.n4663 0.014
R56962 vp_n.n4674 vp_n.n4673 0.014
R56963 vp_n.n4684 vp_n.n4683 0.014
R56964 vp_n.n4694 vp_n.n4693 0.014
R56965 vp_n.n4704 vp_n.n4703 0.014
R56966 vp_n.n9 vp_n.n1 0.013
R56967 vp_n.n19 vp_n.n11 0.013
R56968 vp_n.n29 vp_n.n21 0.013
R56969 vp_n.n39 vp_n.n31 0.013
R56970 vp_n.n49 vp_n.n41 0.013
R56971 vp_n.n59 vp_n.n51 0.013
R56972 vp_n.n69 vp_n.n61 0.013
R56973 vp_n.n79 vp_n.n71 0.013
R56974 vp_n.n89 vp_n.n81 0.013
R56975 vp_n.n99 vp_n.n91 0.013
R56976 vp_n.n109 vp_n.n101 0.013
R56977 vp_n.n119 vp_n.n111 0.013
R56978 vp_n.n129 vp_n.n121 0.013
R56979 vp_n.n139 vp_n.n131 0.013
R56980 vp_n.n149 vp_n.n141 0.013
R56981 vp_n.n159 vp_n.n151 0.013
R56982 vp_n.n169 vp_n.n161 0.013
R56983 vp_n.n179 vp_n.n171 0.013
R56984 vp_n.n189 vp_n.n181 0.013
R56985 vp_n.n199 vp_n.n191 0.013
R56986 vp_n.n209 vp_n.n201 0.013
R56987 vp_n.n219 vp_n.n211 0.013
R56988 vp_n.n229 vp_n.n221 0.013
R56989 vp_n.n239 vp_n.n231 0.013
R56990 vp_n.n249 vp_n.n241 0.013
R56991 vp_n.n259 vp_n.n251 0.013
R56992 vp_n.n269 vp_n.n261 0.013
R56993 vp_n.n279 vp_n.n271 0.013
R56994 vp_n.n289 vp_n.n281 0.013
R56995 vp_n.n299 vp_n.n291 0.013
R56996 vp_n.n309 vp_n.n301 0.013
R56997 vp_n.n319 vp_n.n311 0.013
R56998 vp_n.n329 vp_n.n321 0.013
R56999 vp_n.n339 vp_n.n331 0.013
R57000 vp_n.n349 vp_n.n341 0.013
R57001 vp_n.n359 vp_n.n351 0.013
R57002 vp_n.n369 vp_n.n361 0.013
R57003 vp_n.n379 vp_n.n371 0.013
R57004 vp_n.n389 vp_n.n381 0.013
R57005 vp_n.n399 vp_n.n391 0.013
R57006 vp_n.n409 vp_n.n401 0.013
R57007 vp_n.n419 vp_n.n411 0.013
R57008 vp_n.n429 vp_n.n421 0.013
R57009 vp_n.n439 vp_n.n431 0.013
R57010 vp_n.n449 vp_n.n441 0.013
R57011 vp_n.n459 vp_n.n451 0.013
R57012 vp_n.n469 vp_n.n461 0.013
R57013 vp_n.n479 vp_n.n471 0.013
R57014 vp_n.n489 vp_n.n481 0.013
R57015 vp_n.n499 vp_n.n491 0.013
R57016 vp_n.n509 vp_n.n501 0.013
R57017 vp_n.n519 vp_n.n511 0.013
R57018 vp_n.n529 vp_n.n521 0.013
R57019 vp_n.n539 vp_n.n531 0.013
R57020 vp_n.n549 vp_n.n541 0.013
R57021 vp_n.n559 vp_n.n551 0.013
R57022 vp_n.n569 vp_n.n561 0.013
R57023 vp_n.n579 vp_n.n571 0.013
R57024 vp_n.n589 vp_n.n581 0.013
R57025 vp_n.n599 vp_n.n591 0.013
R57026 vp_n.n609 vp_n.n601 0.013
R57027 vp_n.n619 vp_n.n611 0.013
R57028 vp_n.n629 vp_n.n621 0.013
R57029 vp_n.n639 vp_n.n631 0.013
R57030 vp_n.n649 vp_n.n641 0.013
R57031 vp_n.n659 vp_n.n651 0.013
R57032 vp_n.n669 vp_n.n661 0.013
R57033 vp_n.n679 vp_n.n671 0.013
R57034 vp_n.n689 vp_n.n681 0.013
R57035 vp_n.n699 vp_n.n691 0.013
R57036 vp_n.n709 vp_n.n701 0.013
R57037 vp_n.n719 vp_n.n711 0.013
R57038 vp_n.n729 vp_n.n721 0.013
R57039 vp_n.n739 vp_n.n731 0.013
R57040 vp_n.n749 vp_n.n741 0.013
R57041 vp_n.n759 vp_n.n751 0.013
R57042 vp_n.n769 vp_n.n761 0.013
R57043 vp_n.n779 vp_n.n771 0.013
R57044 vp_n.n789 vp_n.n781 0.013
R57045 vp_n.n799 vp_n.n791 0.013
R57046 vp_n.n809 vp_n.n801 0.013
R57047 vp_n.n819 vp_n.n811 0.013
R57048 vp_n.n829 vp_n.n821 0.013
R57049 vp_n.n839 vp_n.n831 0.013
R57050 vp_n.n849 vp_n.n841 0.013
R57051 vp_n.n859 vp_n.n851 0.013
R57052 vp_n.n869 vp_n.n861 0.013
R57053 vp_n.n879 vp_n.n871 0.013
R57054 vp_n.n889 vp_n.n881 0.013
R57055 vp_n.n899 vp_n.n891 0.013
R57056 vp_n.n909 vp_n.n901 0.013
R57057 vp_n.n919 vp_n.n911 0.013
R57058 vp_n.n929 vp_n.n921 0.013
R57059 vp_n.n939 vp_n.n931 0.013
R57060 vp_n.n949 vp_n.n941 0.013
R57061 vp_n.n959 vp_n.n951 0.013
R57062 vp_n.n969 vp_n.n961 0.013
R57063 vp_n.n979 vp_n.n971 0.013
R57064 vp_n.n989 vp_n.n981 0.013
R57065 vp_n.n999 vp_n.n991 0.013
R57066 vp_n.n1009 vp_n.n1001 0.013
R57067 vp_n.n1019 vp_n.n1011 0.013
R57068 vp_n.n1029 vp_n.n1021 0.013
R57069 vp_n.n1039 vp_n.n1031 0.013
R57070 vp_n.n1049 vp_n.n1041 0.013
R57071 vp_n.n1059 vp_n.n1051 0.013
R57072 vp_n.n1069 vp_n.n1061 0.013
R57073 vp_n.n1079 vp_n.n1071 0.013
R57074 vp_n.n1089 vp_n.n1081 0.013
R57075 vp_n.n1099 vp_n.n1091 0.013
R57076 vp_n.n1109 vp_n.n1101 0.013
R57077 vp_n.n1119 vp_n.n1111 0.013
R57078 vp_n.n1129 vp_n.n1121 0.013
R57079 vp_n.n1139 vp_n.n1131 0.013
R57080 vp_n.n1149 vp_n.n1141 0.013
R57081 vp_n.n1159 vp_n.n1151 0.013
R57082 vp_n.n1169 vp_n.n1161 0.013
R57083 vp_n.n1179 vp_n.n1171 0.013
R57084 vp_n.n1189 vp_n.n1181 0.013
R57085 vp_n.n1199 vp_n.n1191 0.013
R57086 vp_n.n1209 vp_n.n1201 0.013
R57087 vp_n.n1219 vp_n.n1211 0.013
R57088 vp_n.n1229 vp_n.n1221 0.013
R57089 vp_n.n1239 vp_n.n1231 0.013
R57090 vp_n.n1249 vp_n.n1241 0.013
R57091 vp_n.n1259 vp_n.n1251 0.013
R57092 vp_n.n1269 vp_n.n1261 0.013
R57093 vp_n.n1279 vp_n.n1271 0.013
R57094 vp_n.n1289 vp_n.n1281 0.013
R57095 vp_n.n1299 vp_n.n1291 0.013
R57096 vp_n.n1309 vp_n.n1301 0.013
R57097 vp_n.n1319 vp_n.n1311 0.013
R57098 vp_n.n1329 vp_n.n1321 0.013
R57099 vp_n.n1339 vp_n.n1331 0.013
R57100 vp_n.n1349 vp_n.n1341 0.013
R57101 vp_n.n1359 vp_n.n1351 0.013
R57102 vp_n.n1369 vp_n.n1361 0.013
R57103 vp_n.n1379 vp_n.n1371 0.013
R57104 vp_n.n1389 vp_n.n1381 0.013
R57105 vp_n.n1399 vp_n.n1391 0.013
R57106 vp_n.n1409 vp_n.n1401 0.013
R57107 vp_n.n1419 vp_n.n1411 0.013
R57108 vp_n.n1429 vp_n.n1421 0.013
R57109 vp_n.n1439 vp_n.n1431 0.013
R57110 vp_n.n1449 vp_n.n1441 0.013
R57111 vp_n.n1459 vp_n.n1451 0.013
R57112 vp_n.n1469 vp_n.n1461 0.013
R57113 vp_n.n1479 vp_n.n1471 0.013
R57114 vp_n.n1489 vp_n.n1481 0.013
R57115 vp_n.n1499 vp_n.n1491 0.013
R57116 vp_n.n1560 vp_n.n1552 0.013
R57117 vp_n.n1570 vp_n.n1562 0.013
R57118 vp_n.n1580 vp_n.n1572 0.013
R57119 vp_n.n1590 vp_n.n1582 0.013
R57120 vp_n.n1600 vp_n.n1592 0.013
R57121 vp_n.n1610 vp_n.n1602 0.013
R57122 vp_n.n1620 vp_n.n1612 0.013
R57123 vp_n.n1630 vp_n.n1622 0.013
R57124 vp_n.n1640 vp_n.n1632 0.013
R57125 vp_n.n1650 vp_n.n1642 0.013
R57126 vp_n.n1660 vp_n.n1652 0.013
R57127 vp_n.n1670 vp_n.n1662 0.013
R57128 vp_n.n1680 vp_n.n1672 0.013
R57129 vp_n.n1690 vp_n.n1682 0.013
R57130 vp_n.n1700 vp_n.n1692 0.013
R57131 vp_n.n1710 vp_n.n1702 0.013
R57132 vp_n.n1720 vp_n.n1712 0.013
R57133 vp_n.n1730 vp_n.n1722 0.013
R57134 vp_n.n1740 vp_n.n1732 0.013
R57135 vp_n.n1750 vp_n.n1742 0.013
R57136 vp_n.n1760 vp_n.n1752 0.013
R57137 vp_n.n1770 vp_n.n1762 0.013
R57138 vp_n.n1780 vp_n.n1772 0.013
R57139 vp_n.n1790 vp_n.n1782 0.013
R57140 vp_n.n1800 vp_n.n1792 0.013
R57141 vp_n.n1810 vp_n.n1802 0.013
R57142 vp_n.n1820 vp_n.n1812 0.013
R57143 vp_n.n1830 vp_n.n1822 0.013
R57144 vp_n.n1840 vp_n.n1832 0.013
R57145 vp_n.n1850 vp_n.n1842 0.013
R57146 vp_n.n1860 vp_n.n1852 0.013
R57147 vp_n.n1870 vp_n.n1862 0.013
R57148 vp_n.n1880 vp_n.n1872 0.013
R57149 vp_n.n1890 vp_n.n1882 0.013
R57150 vp_n.n1900 vp_n.n1892 0.013
R57151 vp_n.n1910 vp_n.n1902 0.013
R57152 vp_n.n1920 vp_n.n1912 0.013
R57153 vp_n.n1930 vp_n.n1922 0.013
R57154 vp_n.n1940 vp_n.n1932 0.013
R57155 vp_n.n1950 vp_n.n1942 0.013
R57156 vp_n.n1960 vp_n.n1952 0.013
R57157 vp_n.n1970 vp_n.n1962 0.013
R57158 vp_n.n1980 vp_n.n1972 0.013
R57159 vp_n.n1990 vp_n.n1982 0.013
R57160 vp_n.n2000 vp_n.n1992 0.013
R57161 vp_n.n2010 vp_n.n2002 0.013
R57162 vp_n.n2020 vp_n.n2012 0.013
R57163 vp_n.n2030 vp_n.n2022 0.013
R57164 vp_n.n2040 vp_n.n2032 0.013
R57165 vp_n.n2050 vp_n.n2042 0.013
R57166 vp_n.n2060 vp_n.n2052 0.013
R57167 vp_n.n2070 vp_n.n2062 0.013
R57168 vp_n.n2080 vp_n.n2072 0.013
R57169 vp_n.n2090 vp_n.n2082 0.013
R57170 vp_n.n2100 vp_n.n2092 0.013
R57171 vp_n.n2110 vp_n.n2102 0.013
R57172 vp_n.n2120 vp_n.n2112 0.013
R57173 vp_n.n2130 vp_n.n2122 0.013
R57174 vp_n.n2140 vp_n.n2132 0.013
R57175 vp_n.n2150 vp_n.n2142 0.013
R57176 vp_n.n2160 vp_n.n2152 0.013
R57177 vp_n.n2170 vp_n.n2162 0.013
R57178 vp_n.n2180 vp_n.n2172 0.013
R57179 vp_n.n2190 vp_n.n2182 0.013
R57180 vp_n.n2200 vp_n.n2192 0.013
R57181 vp_n.n2210 vp_n.n2202 0.013
R57182 vp_n.n2220 vp_n.n2212 0.013
R57183 vp_n.n2230 vp_n.n2222 0.013
R57184 vp_n.n2240 vp_n.n2232 0.013
R57185 vp_n.n2250 vp_n.n2242 0.013
R57186 vp_n.n2260 vp_n.n2252 0.013
R57187 vp_n.n2270 vp_n.n2262 0.013
R57188 vp_n.n2280 vp_n.n2272 0.013
R57189 vp_n.n2290 vp_n.n2282 0.013
R57190 vp_n.n2300 vp_n.n2292 0.013
R57191 vp_n.n2310 vp_n.n2302 0.013
R57192 vp_n.n2320 vp_n.n2312 0.013
R57193 vp_n.n2330 vp_n.n2322 0.013
R57194 vp_n.n2340 vp_n.n2332 0.013
R57195 vp_n.n2350 vp_n.n2342 0.013
R57196 vp_n.n2360 vp_n.n2352 0.013
R57197 vp_n.n2370 vp_n.n2362 0.013
R57198 vp_n.n2380 vp_n.n2372 0.013
R57199 vp_n.n2390 vp_n.n2382 0.013
R57200 vp_n.n2400 vp_n.n2392 0.013
R57201 vp_n.n2410 vp_n.n2402 0.013
R57202 vp_n.n2420 vp_n.n2412 0.013
R57203 vp_n.n2430 vp_n.n2422 0.013
R57204 vp_n.n2440 vp_n.n2432 0.013
R57205 vp_n.n2450 vp_n.n2442 0.013
R57206 vp_n.n2460 vp_n.n2452 0.013
R57207 vp_n.n2470 vp_n.n2462 0.013
R57208 vp_n.n2480 vp_n.n2472 0.013
R57209 vp_n.n2490 vp_n.n2482 0.013
R57210 vp_n.n2500 vp_n.n2492 0.013
R57211 vp_n.n2510 vp_n.n2502 0.013
R57212 vp_n.n2520 vp_n.n2512 0.013
R57213 vp_n.n2530 vp_n.n2522 0.013
R57214 vp_n.n2540 vp_n.n2532 0.013
R57215 vp_n.n2550 vp_n.n2542 0.013
R57216 vp_n.n2560 vp_n.n2552 0.013
R57217 vp_n.n2570 vp_n.n2562 0.013
R57218 vp_n.n2580 vp_n.n2572 0.013
R57219 vp_n.n2590 vp_n.n2582 0.013
R57220 vp_n.n2600 vp_n.n2592 0.013
R57221 vp_n.n2610 vp_n.n2602 0.013
R57222 vp_n.n2620 vp_n.n2612 0.013
R57223 vp_n.n2630 vp_n.n2622 0.013
R57224 vp_n.n2640 vp_n.n2632 0.013
R57225 vp_n.n2650 vp_n.n2642 0.013
R57226 vp_n.n2660 vp_n.n2652 0.013
R57227 vp_n.n2670 vp_n.n2662 0.013
R57228 vp_n.n2680 vp_n.n2672 0.013
R57229 vp_n.n2690 vp_n.n2682 0.013
R57230 vp_n.n2700 vp_n.n2692 0.013
R57231 vp_n.n2710 vp_n.n2702 0.013
R57232 vp_n.n2720 vp_n.n2712 0.013
R57233 vp_n.n2730 vp_n.n2722 0.013
R57234 vp_n.n2740 vp_n.n2732 0.013
R57235 vp_n.n2750 vp_n.n2742 0.013
R57236 vp_n.n2760 vp_n.n2752 0.013
R57237 vp_n.n2770 vp_n.n2762 0.013
R57238 vp_n.n2780 vp_n.n2772 0.013
R57239 vp_n.n2790 vp_n.n2782 0.013
R57240 vp_n.n2800 vp_n.n2792 0.013
R57241 vp_n.n2810 vp_n.n2802 0.013
R57242 vp_n.n2820 vp_n.n2812 0.013
R57243 vp_n.n2830 vp_n.n2822 0.013
R57244 vp_n.n2840 vp_n.n2832 0.013
R57245 vp_n.n2850 vp_n.n2842 0.013
R57246 vp_n.n2860 vp_n.n2852 0.013
R57247 vp_n.n2870 vp_n.n2862 0.013
R57248 vp_n.n2880 vp_n.n2872 0.013
R57249 vp_n.n2890 vp_n.n2882 0.013
R57250 vp_n.n2900 vp_n.n2892 0.013
R57251 vp_n.n2910 vp_n.n2902 0.013
R57252 vp_n.n2920 vp_n.n2912 0.013
R57253 vp_n.n2930 vp_n.n2922 0.013
R57254 vp_n.n2940 vp_n.n2932 0.013
R57255 vp_n.n2950 vp_n.n2942 0.013
R57256 vp_n.n2960 vp_n.n2952 0.013
R57257 vp_n.n2970 vp_n.n2962 0.013
R57258 vp_n.n2980 vp_n.n2972 0.013
R57259 vp_n.n2990 vp_n.n2982 0.013
R57260 vp_n.n3000 vp_n.n2992 0.013
R57261 vp_n.n3010 vp_n.n3002 0.013
R57262 vp_n.n3020 vp_n.n3012 0.013
R57263 vp_n.n3030 vp_n.n3022 0.013
R57264 vp_n.n3040 vp_n.n3032 0.013
R57265 vp_n.n3050 vp_n.n3042 0.013
R57266 vp_n.n3213 vp_n.n3205 0.013
R57267 vp_n.n3223 vp_n.n3215 0.013
R57268 vp_n.n3233 vp_n.n3225 0.013
R57269 vp_n.n3243 vp_n.n3235 0.013
R57270 vp_n.n3253 vp_n.n3245 0.013
R57271 vp_n.n3263 vp_n.n3255 0.013
R57272 vp_n.n3273 vp_n.n3265 0.013
R57273 vp_n.n3283 vp_n.n3275 0.013
R57274 vp_n.n3293 vp_n.n3285 0.013
R57275 vp_n.n3303 vp_n.n3295 0.013
R57276 vp_n.n3313 vp_n.n3305 0.013
R57277 vp_n.n3323 vp_n.n3315 0.013
R57278 vp_n.n3333 vp_n.n3325 0.013
R57279 vp_n.n3343 vp_n.n3335 0.013
R57280 vp_n.n3353 vp_n.n3345 0.013
R57281 vp_n.n3363 vp_n.n3355 0.013
R57282 vp_n.n3373 vp_n.n3365 0.013
R57283 vp_n.n3383 vp_n.n3375 0.013
R57284 vp_n.n3393 vp_n.n3385 0.013
R57285 vp_n.n3403 vp_n.n3395 0.013
R57286 vp_n.n3413 vp_n.n3405 0.013
R57287 vp_n.n3423 vp_n.n3415 0.013
R57288 vp_n.n3433 vp_n.n3425 0.013
R57289 vp_n.n3443 vp_n.n3435 0.013
R57290 vp_n.n3453 vp_n.n3445 0.013
R57291 vp_n.n3463 vp_n.n3455 0.013
R57292 vp_n.n3473 vp_n.n3465 0.013
R57293 vp_n.n3483 vp_n.n3475 0.013
R57294 vp_n.n3493 vp_n.n3485 0.013
R57295 vp_n.n3503 vp_n.n3495 0.013
R57296 vp_n.n3513 vp_n.n3505 0.013
R57297 vp_n.n3523 vp_n.n3515 0.013
R57298 vp_n.n3533 vp_n.n3525 0.013
R57299 vp_n.n3543 vp_n.n3535 0.013
R57300 vp_n.n3553 vp_n.n3545 0.013
R57301 vp_n.n3563 vp_n.n3555 0.013
R57302 vp_n.n3573 vp_n.n3565 0.013
R57303 vp_n.n3583 vp_n.n3575 0.013
R57304 vp_n.n3593 vp_n.n3585 0.013
R57305 vp_n.n3603 vp_n.n3595 0.013
R57306 vp_n.n3613 vp_n.n3605 0.013
R57307 vp_n.n3623 vp_n.n3615 0.013
R57308 vp_n.n3633 vp_n.n3625 0.013
R57309 vp_n.n3643 vp_n.n3635 0.013
R57310 vp_n.n3653 vp_n.n3645 0.013
R57311 vp_n.n3663 vp_n.n3655 0.013
R57312 vp_n.n3673 vp_n.n3665 0.013
R57313 vp_n.n3683 vp_n.n3675 0.013
R57314 vp_n.n3693 vp_n.n3685 0.013
R57315 vp_n.n3703 vp_n.n3695 0.013
R57316 vp_n.n3713 vp_n.n3705 0.013
R57317 vp_n.n3723 vp_n.n3715 0.013
R57318 vp_n.n3733 vp_n.n3725 0.013
R57319 vp_n.n3743 vp_n.n3735 0.013
R57320 vp_n.n3753 vp_n.n3745 0.013
R57321 vp_n.n3763 vp_n.n3755 0.013
R57322 vp_n.n3773 vp_n.n3765 0.013
R57323 vp_n.n3783 vp_n.n3775 0.013
R57324 vp_n.n3793 vp_n.n3785 0.013
R57325 vp_n.n3803 vp_n.n3795 0.013
R57326 vp_n.n3813 vp_n.n3805 0.013
R57327 vp_n.n3823 vp_n.n3815 0.013
R57328 vp_n.n3833 vp_n.n3825 0.013
R57329 vp_n.n3843 vp_n.n3835 0.013
R57330 vp_n.n3853 vp_n.n3845 0.013
R57331 vp_n.n3863 vp_n.n3855 0.013
R57332 vp_n.n3873 vp_n.n3865 0.013
R57333 vp_n.n3883 vp_n.n3875 0.013
R57334 vp_n.n3893 vp_n.n3885 0.013
R57335 vp_n.n3903 vp_n.n3895 0.013
R57336 vp_n.n3913 vp_n.n3905 0.013
R57337 vp_n.n3923 vp_n.n3915 0.013
R57338 vp_n.n3933 vp_n.n3925 0.013
R57339 vp_n.n3943 vp_n.n3935 0.013
R57340 vp_n.n3953 vp_n.n3945 0.013
R57341 vp_n.n3963 vp_n.n3955 0.013
R57342 vp_n.n3973 vp_n.n3965 0.013
R57343 vp_n.n3983 vp_n.n3975 0.013
R57344 vp_n.n3993 vp_n.n3985 0.013
R57345 vp_n.n4003 vp_n.n3995 0.013
R57346 vp_n.n4013 vp_n.n4005 0.013
R57347 vp_n.n4023 vp_n.n4015 0.013
R57348 vp_n.n4033 vp_n.n4025 0.013
R57349 vp_n.n4043 vp_n.n4035 0.013
R57350 vp_n.n4053 vp_n.n4045 0.013
R57351 vp_n.n4063 vp_n.n4055 0.013
R57352 vp_n.n4073 vp_n.n4065 0.013
R57353 vp_n.n4083 vp_n.n4075 0.013
R57354 vp_n.n4093 vp_n.n4085 0.013
R57355 vp_n.n4103 vp_n.n4095 0.013
R57356 vp_n.n4113 vp_n.n4105 0.013
R57357 vp_n.n4123 vp_n.n4115 0.013
R57358 vp_n.n4133 vp_n.n4125 0.013
R57359 vp_n.n4143 vp_n.n4135 0.013
R57360 vp_n.n4153 vp_n.n4145 0.013
R57361 vp_n.n4163 vp_n.n4155 0.013
R57362 vp_n.n4173 vp_n.n4165 0.013
R57363 vp_n.n4183 vp_n.n4175 0.013
R57364 vp_n.n4193 vp_n.n4185 0.013
R57365 vp_n.n4203 vp_n.n4195 0.013
R57366 vp_n.n4213 vp_n.n4205 0.013
R57367 vp_n.n4223 vp_n.n4215 0.013
R57368 vp_n.n4233 vp_n.n4225 0.013
R57369 vp_n.n4243 vp_n.n4235 0.013
R57370 vp_n.n4253 vp_n.n4245 0.013
R57371 vp_n.n4263 vp_n.n4255 0.013
R57372 vp_n.n4273 vp_n.n4265 0.013
R57373 vp_n.n4283 vp_n.n4275 0.013
R57374 vp_n.n4293 vp_n.n4285 0.013
R57375 vp_n.n4303 vp_n.n4295 0.013
R57376 vp_n.n4313 vp_n.n4305 0.013
R57377 vp_n.n4323 vp_n.n4315 0.013
R57378 vp_n.n4333 vp_n.n4325 0.013
R57379 vp_n.n4343 vp_n.n4335 0.013
R57380 vp_n.n4353 vp_n.n4345 0.013
R57381 vp_n.n4363 vp_n.n4355 0.013
R57382 vp_n.n4373 vp_n.n4365 0.013
R57383 vp_n.n4383 vp_n.n4375 0.013
R57384 vp_n.n4393 vp_n.n4385 0.013
R57385 vp_n.n4403 vp_n.n4395 0.013
R57386 vp_n.n4413 vp_n.n4405 0.013
R57387 vp_n.n4423 vp_n.n4415 0.013
R57388 vp_n.n4433 vp_n.n4425 0.013
R57389 vp_n.n4443 vp_n.n4435 0.013
R57390 vp_n.n4453 vp_n.n4445 0.013
R57391 vp_n.n4463 vp_n.n4455 0.013
R57392 vp_n.n4473 vp_n.n4465 0.013
R57393 vp_n.n4483 vp_n.n4475 0.013
R57394 vp_n.n4493 vp_n.n4485 0.013
R57395 vp_n.n4503 vp_n.n4495 0.013
R57396 vp_n.n4513 vp_n.n4505 0.013
R57397 vp_n.n4523 vp_n.n4515 0.013
R57398 vp_n.n4533 vp_n.n4525 0.013
R57399 vp_n.n4543 vp_n.n4535 0.013
R57400 vp_n.n4553 vp_n.n4545 0.013
R57401 vp_n.n4563 vp_n.n4555 0.013
R57402 vp_n.n4573 vp_n.n4565 0.013
R57403 vp_n.n4583 vp_n.n4575 0.013
R57404 vp_n.n4593 vp_n.n4585 0.013
R57405 vp_n.n4603 vp_n.n4595 0.013
R57406 vp_n.n4613 vp_n.n4605 0.013
R57407 vp_n.n4623 vp_n.n4615 0.013
R57408 vp_n.n4633 vp_n.n4625 0.013
R57409 vp_n.n4643 vp_n.n4635 0.013
R57410 vp_n.n4653 vp_n.n4645 0.013
R57411 vp_n.n4663 vp_n.n4655 0.013
R57412 vp_n.n4673 vp_n.n4665 0.013
R57413 vp_n.n4683 vp_n.n4675 0.013
R57414 vp_n.n4693 vp_n.n4685 0.013
R57415 vp_n.n4703 vp_n.n4695 0.013
R57416 vp_n.n9 vp_n.n8 0.002
R57417 vp_n.n19 vp_n.n18 0.002
R57418 vp_n.n29 vp_n.n28 0.002
R57419 vp_n.n39 vp_n.n38 0.002
R57420 vp_n.n49 vp_n.n48 0.002
R57421 vp_n.n59 vp_n.n58 0.002
R57422 vp_n.n69 vp_n.n68 0.002
R57423 vp_n.n79 vp_n.n78 0.002
R57424 vp_n.n89 vp_n.n88 0.002
R57425 vp_n.n99 vp_n.n98 0.002
R57426 vp_n.n109 vp_n.n108 0.002
R57427 vp_n.n119 vp_n.n118 0.002
R57428 vp_n.n129 vp_n.n128 0.002
R57429 vp_n.n139 vp_n.n138 0.002
R57430 vp_n.n149 vp_n.n148 0.002
R57431 vp_n.n159 vp_n.n158 0.002
R57432 vp_n.n169 vp_n.n168 0.002
R57433 vp_n.n179 vp_n.n178 0.002
R57434 vp_n.n189 vp_n.n188 0.002
R57435 vp_n.n199 vp_n.n198 0.002
R57436 vp_n.n209 vp_n.n208 0.002
R57437 vp_n.n219 vp_n.n218 0.002
R57438 vp_n.n229 vp_n.n228 0.002
R57439 vp_n.n239 vp_n.n238 0.002
R57440 vp_n.n249 vp_n.n248 0.002
R57441 vp_n.n259 vp_n.n258 0.002
R57442 vp_n.n269 vp_n.n268 0.002
R57443 vp_n.n279 vp_n.n278 0.002
R57444 vp_n.n289 vp_n.n288 0.002
R57445 vp_n.n299 vp_n.n298 0.002
R57446 vp_n.n309 vp_n.n308 0.002
R57447 vp_n.n319 vp_n.n318 0.002
R57448 vp_n.n329 vp_n.n328 0.002
R57449 vp_n.n339 vp_n.n338 0.002
R57450 vp_n.n349 vp_n.n348 0.002
R57451 vp_n.n359 vp_n.n358 0.002
R57452 vp_n.n369 vp_n.n368 0.002
R57453 vp_n.n379 vp_n.n378 0.002
R57454 vp_n.n389 vp_n.n388 0.002
R57455 vp_n.n399 vp_n.n398 0.002
R57456 vp_n.n409 vp_n.n408 0.002
R57457 vp_n.n419 vp_n.n418 0.002
R57458 vp_n.n429 vp_n.n428 0.002
R57459 vp_n.n439 vp_n.n438 0.002
R57460 vp_n.n449 vp_n.n448 0.002
R57461 vp_n.n459 vp_n.n458 0.002
R57462 vp_n.n469 vp_n.n468 0.002
R57463 vp_n.n479 vp_n.n478 0.002
R57464 vp_n.n489 vp_n.n488 0.002
R57465 vp_n.n499 vp_n.n498 0.002
R57466 vp_n.n509 vp_n.n508 0.002
R57467 vp_n.n519 vp_n.n518 0.002
R57468 vp_n.n529 vp_n.n528 0.002
R57469 vp_n.n539 vp_n.n538 0.002
R57470 vp_n.n549 vp_n.n548 0.002
R57471 vp_n.n559 vp_n.n558 0.002
R57472 vp_n.n569 vp_n.n568 0.002
R57473 vp_n.n579 vp_n.n578 0.002
R57474 vp_n.n589 vp_n.n588 0.002
R57475 vp_n.n599 vp_n.n598 0.002
R57476 vp_n.n609 vp_n.n608 0.002
R57477 vp_n.n619 vp_n.n618 0.002
R57478 vp_n.n629 vp_n.n628 0.002
R57479 vp_n.n639 vp_n.n638 0.002
R57480 vp_n.n649 vp_n.n648 0.002
R57481 vp_n.n659 vp_n.n658 0.002
R57482 vp_n.n669 vp_n.n668 0.002
R57483 vp_n.n679 vp_n.n678 0.002
R57484 vp_n.n689 vp_n.n688 0.002
R57485 vp_n.n699 vp_n.n698 0.002
R57486 vp_n.n709 vp_n.n708 0.002
R57487 vp_n.n719 vp_n.n718 0.002
R57488 vp_n.n729 vp_n.n728 0.002
R57489 vp_n.n739 vp_n.n738 0.002
R57490 vp_n.n749 vp_n.n748 0.002
R57491 vp_n.n759 vp_n.n758 0.002
R57492 vp_n.n769 vp_n.n768 0.002
R57493 vp_n.n779 vp_n.n778 0.002
R57494 vp_n.n789 vp_n.n788 0.002
R57495 vp_n.n799 vp_n.n798 0.002
R57496 vp_n.n809 vp_n.n808 0.002
R57497 vp_n.n819 vp_n.n818 0.002
R57498 vp_n.n829 vp_n.n828 0.002
R57499 vp_n.n839 vp_n.n838 0.002
R57500 vp_n.n849 vp_n.n848 0.002
R57501 vp_n.n859 vp_n.n858 0.002
R57502 vp_n.n869 vp_n.n868 0.002
R57503 vp_n.n879 vp_n.n878 0.002
R57504 vp_n.n889 vp_n.n888 0.002
R57505 vp_n.n899 vp_n.n898 0.002
R57506 vp_n.n909 vp_n.n908 0.002
R57507 vp_n.n919 vp_n.n918 0.002
R57508 vp_n.n929 vp_n.n928 0.002
R57509 vp_n.n939 vp_n.n938 0.002
R57510 vp_n.n949 vp_n.n948 0.002
R57511 vp_n.n959 vp_n.n958 0.002
R57512 vp_n.n969 vp_n.n968 0.002
R57513 vp_n.n979 vp_n.n978 0.002
R57514 vp_n.n989 vp_n.n988 0.002
R57515 vp_n.n999 vp_n.n998 0.002
R57516 vp_n.n1009 vp_n.n1008 0.002
R57517 vp_n.n1019 vp_n.n1018 0.002
R57518 vp_n.n1029 vp_n.n1028 0.002
R57519 vp_n.n1039 vp_n.n1038 0.002
R57520 vp_n.n1049 vp_n.n1048 0.002
R57521 vp_n.n1059 vp_n.n1058 0.002
R57522 vp_n.n1069 vp_n.n1068 0.002
R57523 vp_n.n1079 vp_n.n1078 0.002
R57524 vp_n.n1089 vp_n.n1088 0.002
R57525 vp_n.n1099 vp_n.n1098 0.002
R57526 vp_n.n1109 vp_n.n1108 0.002
R57527 vp_n.n1119 vp_n.n1118 0.002
R57528 vp_n.n1129 vp_n.n1128 0.002
R57529 vp_n.n1139 vp_n.n1138 0.002
R57530 vp_n.n1149 vp_n.n1148 0.002
R57531 vp_n.n1159 vp_n.n1158 0.002
R57532 vp_n.n1169 vp_n.n1168 0.002
R57533 vp_n.n1179 vp_n.n1178 0.002
R57534 vp_n.n1189 vp_n.n1188 0.002
R57535 vp_n.n1199 vp_n.n1198 0.002
R57536 vp_n.n1209 vp_n.n1208 0.002
R57537 vp_n.n1219 vp_n.n1218 0.002
R57538 vp_n.n1229 vp_n.n1228 0.002
R57539 vp_n.n1239 vp_n.n1238 0.002
R57540 vp_n.n1249 vp_n.n1248 0.002
R57541 vp_n.n1259 vp_n.n1258 0.002
R57542 vp_n.n1269 vp_n.n1268 0.002
R57543 vp_n.n1279 vp_n.n1278 0.002
R57544 vp_n.n1289 vp_n.n1288 0.002
R57545 vp_n.n1299 vp_n.n1298 0.002
R57546 vp_n.n1309 vp_n.n1308 0.002
R57547 vp_n.n1319 vp_n.n1318 0.002
R57548 vp_n.n1329 vp_n.n1328 0.002
R57549 vp_n.n1339 vp_n.n1338 0.002
R57550 vp_n.n1349 vp_n.n1348 0.002
R57551 vp_n.n1359 vp_n.n1358 0.002
R57552 vp_n.n1369 vp_n.n1368 0.002
R57553 vp_n.n1379 vp_n.n1378 0.002
R57554 vp_n.n1389 vp_n.n1388 0.002
R57555 vp_n.n1399 vp_n.n1398 0.002
R57556 vp_n.n1409 vp_n.n1408 0.002
R57557 vp_n.n1419 vp_n.n1418 0.002
R57558 vp_n.n1429 vp_n.n1428 0.002
R57559 vp_n.n1439 vp_n.n1438 0.002
R57560 vp_n.n1449 vp_n.n1448 0.002
R57561 vp_n.n1459 vp_n.n1458 0.002
R57562 vp_n.n1469 vp_n.n1468 0.002
R57563 vp_n.n1479 vp_n.n1478 0.002
R57564 vp_n.n1489 vp_n.n1488 0.002
R57565 vp_n.n1499 vp_n.n1498 0.002
R57566 vp_n.n1560 vp_n.n1559 0.002
R57567 vp_n.n1580 vp_n.n1579 0.002
R57568 vp_n.n1590 vp_n.n1589 0.002
R57569 vp_n.n1600 vp_n.n1599 0.002
R57570 vp_n.n1610 vp_n.n1609 0.002
R57571 vp_n.n1620 vp_n.n1619 0.002
R57572 vp_n.n1630 vp_n.n1629 0.002
R57573 vp_n.n1640 vp_n.n1639 0.002
R57574 vp_n.n1650 vp_n.n1649 0.002
R57575 vp_n.n1660 vp_n.n1659 0.002
R57576 vp_n.n1670 vp_n.n1669 0.002
R57577 vp_n.n1680 vp_n.n1679 0.002
R57578 vp_n.n1690 vp_n.n1689 0.002
R57579 vp_n.n1700 vp_n.n1699 0.002
R57580 vp_n.n1710 vp_n.n1709 0.002
R57581 vp_n.n1720 vp_n.n1719 0.002
R57582 vp_n.n1730 vp_n.n1729 0.002
R57583 vp_n.n1740 vp_n.n1739 0.002
R57584 vp_n.n1750 vp_n.n1749 0.002
R57585 vp_n.n1760 vp_n.n1759 0.002
R57586 vp_n.n1770 vp_n.n1769 0.002
R57587 vp_n.n1780 vp_n.n1779 0.002
R57588 vp_n.n1790 vp_n.n1789 0.002
R57589 vp_n.n1800 vp_n.n1799 0.002
R57590 vp_n.n1810 vp_n.n1809 0.002
R57591 vp_n.n1820 vp_n.n1819 0.002
R57592 vp_n.n1830 vp_n.n1829 0.002
R57593 vp_n.n1840 vp_n.n1839 0.002
R57594 vp_n.n1850 vp_n.n1849 0.002
R57595 vp_n.n1860 vp_n.n1859 0.002
R57596 vp_n.n1870 vp_n.n1869 0.002
R57597 vp_n.n1880 vp_n.n1879 0.002
R57598 vp_n.n1890 vp_n.n1889 0.002
R57599 vp_n.n1900 vp_n.n1899 0.002
R57600 vp_n.n1910 vp_n.n1909 0.002
R57601 vp_n.n1920 vp_n.n1919 0.002
R57602 vp_n.n1930 vp_n.n1929 0.002
R57603 vp_n.n1940 vp_n.n1939 0.002
R57604 vp_n.n1950 vp_n.n1949 0.002
R57605 vp_n.n1960 vp_n.n1959 0.002
R57606 vp_n.n1970 vp_n.n1969 0.002
R57607 vp_n.n1980 vp_n.n1979 0.002
R57608 vp_n.n1990 vp_n.n1989 0.002
R57609 vp_n.n2000 vp_n.n1999 0.002
R57610 vp_n.n2010 vp_n.n2009 0.002
R57611 vp_n.n2020 vp_n.n2019 0.002
R57612 vp_n.n2030 vp_n.n2029 0.002
R57613 vp_n.n2040 vp_n.n2039 0.002
R57614 vp_n.n2050 vp_n.n2049 0.002
R57615 vp_n.n2060 vp_n.n2059 0.002
R57616 vp_n.n2070 vp_n.n2069 0.002
R57617 vp_n.n2080 vp_n.n2079 0.002
R57618 vp_n.n2090 vp_n.n2089 0.002
R57619 vp_n.n2100 vp_n.n2099 0.002
R57620 vp_n.n2110 vp_n.n2109 0.002
R57621 vp_n.n2120 vp_n.n2119 0.002
R57622 vp_n.n2130 vp_n.n2129 0.002
R57623 vp_n.n2140 vp_n.n2139 0.002
R57624 vp_n.n2150 vp_n.n2149 0.002
R57625 vp_n.n2160 vp_n.n2159 0.002
R57626 vp_n.n2170 vp_n.n2169 0.002
R57627 vp_n.n2180 vp_n.n2179 0.002
R57628 vp_n.n2190 vp_n.n2189 0.002
R57629 vp_n.n2200 vp_n.n2199 0.002
R57630 vp_n.n2210 vp_n.n2209 0.002
R57631 vp_n.n2220 vp_n.n2219 0.002
R57632 vp_n.n2230 vp_n.n2229 0.002
R57633 vp_n.n2240 vp_n.n2239 0.002
R57634 vp_n.n2250 vp_n.n2249 0.002
R57635 vp_n.n2260 vp_n.n2259 0.002
R57636 vp_n.n2270 vp_n.n2269 0.002
R57637 vp_n.n2280 vp_n.n2279 0.002
R57638 vp_n.n2290 vp_n.n2289 0.002
R57639 vp_n.n2300 vp_n.n2299 0.002
R57640 vp_n.n2310 vp_n.n2309 0.002
R57641 vp_n.n2320 vp_n.n2319 0.002
R57642 vp_n.n2330 vp_n.n2329 0.002
R57643 vp_n.n2340 vp_n.n2339 0.002
R57644 vp_n.n2350 vp_n.n2349 0.002
R57645 vp_n.n2360 vp_n.n2359 0.002
R57646 vp_n.n2370 vp_n.n2369 0.002
R57647 vp_n.n2380 vp_n.n2379 0.002
R57648 vp_n.n2390 vp_n.n2389 0.002
R57649 vp_n.n2400 vp_n.n2399 0.002
R57650 vp_n.n2410 vp_n.n2409 0.002
R57651 vp_n.n2420 vp_n.n2419 0.002
R57652 vp_n.n2430 vp_n.n2429 0.002
R57653 vp_n.n2440 vp_n.n2439 0.002
R57654 vp_n.n2450 vp_n.n2449 0.002
R57655 vp_n.n2460 vp_n.n2459 0.002
R57656 vp_n.n2470 vp_n.n2469 0.002
R57657 vp_n.n2480 vp_n.n2479 0.002
R57658 vp_n.n2490 vp_n.n2489 0.002
R57659 vp_n.n2500 vp_n.n2499 0.002
R57660 vp_n.n2510 vp_n.n2509 0.002
R57661 vp_n.n2520 vp_n.n2519 0.002
R57662 vp_n.n2530 vp_n.n2529 0.002
R57663 vp_n.n2540 vp_n.n2539 0.002
R57664 vp_n.n2550 vp_n.n2549 0.002
R57665 vp_n.n2560 vp_n.n2559 0.002
R57666 vp_n.n2570 vp_n.n2569 0.002
R57667 vp_n.n2580 vp_n.n2579 0.002
R57668 vp_n.n2590 vp_n.n2589 0.002
R57669 vp_n.n2600 vp_n.n2599 0.002
R57670 vp_n.n2610 vp_n.n2609 0.002
R57671 vp_n.n2620 vp_n.n2619 0.002
R57672 vp_n.n2630 vp_n.n2629 0.002
R57673 vp_n.n2640 vp_n.n2639 0.002
R57674 vp_n.n2650 vp_n.n2649 0.002
R57675 vp_n.n2660 vp_n.n2659 0.002
R57676 vp_n.n2670 vp_n.n2669 0.002
R57677 vp_n.n2680 vp_n.n2679 0.002
R57678 vp_n.n2690 vp_n.n2689 0.002
R57679 vp_n.n2700 vp_n.n2699 0.002
R57680 vp_n.n2710 vp_n.n2709 0.002
R57681 vp_n.n2720 vp_n.n2719 0.002
R57682 vp_n.n2730 vp_n.n2729 0.002
R57683 vp_n.n2740 vp_n.n2739 0.002
R57684 vp_n.n2750 vp_n.n2749 0.002
R57685 vp_n.n2760 vp_n.n2759 0.002
R57686 vp_n.n2770 vp_n.n2769 0.002
R57687 vp_n.n2780 vp_n.n2779 0.002
R57688 vp_n.n2790 vp_n.n2789 0.002
R57689 vp_n.n2800 vp_n.n2799 0.002
R57690 vp_n.n2810 vp_n.n2809 0.002
R57691 vp_n.n2820 vp_n.n2819 0.002
R57692 vp_n.n2830 vp_n.n2829 0.002
R57693 vp_n.n2840 vp_n.n2839 0.002
R57694 vp_n.n2850 vp_n.n2849 0.002
R57695 vp_n.n2860 vp_n.n2859 0.002
R57696 vp_n.n2870 vp_n.n2869 0.002
R57697 vp_n.n2880 vp_n.n2879 0.002
R57698 vp_n.n2890 vp_n.n2889 0.002
R57699 vp_n.n2900 vp_n.n2899 0.002
R57700 vp_n.n2910 vp_n.n2909 0.002
R57701 vp_n.n2920 vp_n.n2919 0.002
R57702 vp_n.n2930 vp_n.n2929 0.002
R57703 vp_n.n2940 vp_n.n2939 0.002
R57704 vp_n.n2950 vp_n.n2949 0.002
R57705 vp_n.n2960 vp_n.n2959 0.002
R57706 vp_n.n2970 vp_n.n2969 0.002
R57707 vp_n.n2980 vp_n.n2979 0.002
R57708 vp_n.n2990 vp_n.n2989 0.002
R57709 vp_n.n3000 vp_n.n2999 0.002
R57710 vp_n.n3010 vp_n.n3009 0.002
R57711 vp_n.n3020 vp_n.n3019 0.002
R57712 vp_n.n3030 vp_n.n3029 0.002
R57713 vp_n.n3040 vp_n.n3039 0.002
R57714 vp_n.n3050 vp_n.n3049 0.002
R57715 vp_n.n1570 vp_n.n1569 0.002
R57716 vp_n.n4703 vp_n.n4702 0.002
R57717 vp_n.n4693 vp_n.n4692 0.002
R57718 vp_n.n4683 vp_n.n4682 0.002
R57719 vp_n.n4673 vp_n.n4672 0.002
R57720 vp_n.n4663 vp_n.n4662 0.002
R57721 vp_n.n4653 vp_n.n4652 0.002
R57722 vp_n.n4643 vp_n.n4642 0.002
R57723 vp_n.n4633 vp_n.n4632 0.002
R57724 vp_n.n4623 vp_n.n4622 0.002
R57725 vp_n.n4613 vp_n.n4612 0.002
R57726 vp_n.n4603 vp_n.n4602 0.002
R57727 vp_n.n4593 vp_n.n4592 0.002
R57728 vp_n.n4583 vp_n.n4582 0.002
R57729 vp_n.n4573 vp_n.n4572 0.002
R57730 vp_n.n4563 vp_n.n4562 0.002
R57731 vp_n.n4553 vp_n.n4552 0.002
R57732 vp_n.n4543 vp_n.n4542 0.002
R57733 vp_n.n4533 vp_n.n4532 0.002
R57734 vp_n.n4523 vp_n.n4522 0.002
R57735 vp_n.n4513 vp_n.n4512 0.002
R57736 vp_n.n4503 vp_n.n4502 0.002
R57737 vp_n.n4493 vp_n.n4492 0.002
R57738 vp_n.n4483 vp_n.n4482 0.002
R57739 vp_n.n4473 vp_n.n4472 0.002
R57740 vp_n.n4463 vp_n.n4462 0.002
R57741 vp_n.n4453 vp_n.n4452 0.002
R57742 vp_n.n4443 vp_n.n4442 0.002
R57743 vp_n.n4433 vp_n.n4432 0.002
R57744 vp_n.n4423 vp_n.n4422 0.002
R57745 vp_n.n4413 vp_n.n4412 0.002
R57746 vp_n.n4403 vp_n.n4402 0.002
R57747 vp_n.n4393 vp_n.n4392 0.002
R57748 vp_n.n4383 vp_n.n4382 0.002
R57749 vp_n.n4373 vp_n.n4372 0.002
R57750 vp_n.n4363 vp_n.n4362 0.002
R57751 vp_n.n4353 vp_n.n4352 0.002
R57752 vp_n.n4343 vp_n.n4342 0.002
R57753 vp_n.n4333 vp_n.n4332 0.002
R57754 vp_n.n4323 vp_n.n4322 0.002
R57755 vp_n.n4313 vp_n.n4312 0.002
R57756 vp_n.n4303 vp_n.n4302 0.002
R57757 vp_n.n4293 vp_n.n4292 0.002
R57758 vp_n.n4283 vp_n.n4282 0.002
R57759 vp_n.n4273 vp_n.n4272 0.002
R57760 vp_n.n4263 vp_n.n4262 0.002
R57761 vp_n.n4253 vp_n.n4252 0.002
R57762 vp_n.n4243 vp_n.n4242 0.002
R57763 vp_n.n4233 vp_n.n4232 0.002
R57764 vp_n.n4223 vp_n.n4222 0.002
R57765 vp_n.n4213 vp_n.n4212 0.002
R57766 vp_n.n4203 vp_n.n4202 0.002
R57767 vp_n.n4193 vp_n.n4192 0.002
R57768 vp_n.n4183 vp_n.n4182 0.002
R57769 vp_n.n4173 vp_n.n4172 0.002
R57770 vp_n.n4163 vp_n.n4162 0.002
R57771 vp_n.n4153 vp_n.n4152 0.002
R57772 vp_n.n4143 vp_n.n4142 0.002
R57773 vp_n.n4133 vp_n.n4132 0.002
R57774 vp_n.n4123 vp_n.n4122 0.002
R57775 vp_n.n4113 vp_n.n4112 0.002
R57776 vp_n.n4103 vp_n.n4102 0.002
R57777 vp_n.n4093 vp_n.n4092 0.002
R57778 vp_n.n4083 vp_n.n4082 0.002
R57779 vp_n.n4073 vp_n.n4072 0.002
R57780 vp_n.n4063 vp_n.n4062 0.002
R57781 vp_n.n4053 vp_n.n4052 0.002
R57782 vp_n.n4043 vp_n.n4042 0.002
R57783 vp_n.n4033 vp_n.n4032 0.002
R57784 vp_n.n4023 vp_n.n4022 0.002
R57785 vp_n.n4013 vp_n.n4012 0.002
R57786 vp_n.n4003 vp_n.n4002 0.002
R57787 vp_n.n3993 vp_n.n3992 0.002
R57788 vp_n.n3983 vp_n.n3982 0.002
R57789 vp_n.n3973 vp_n.n3972 0.002
R57790 vp_n.n3963 vp_n.n3962 0.002
R57791 vp_n.n3953 vp_n.n3952 0.002
R57792 vp_n.n3943 vp_n.n3942 0.002
R57793 vp_n.n3933 vp_n.n3932 0.002
R57794 vp_n.n3923 vp_n.n3922 0.002
R57795 vp_n.n3913 vp_n.n3912 0.002
R57796 vp_n.n3903 vp_n.n3902 0.002
R57797 vp_n.n3893 vp_n.n3892 0.002
R57798 vp_n.n3883 vp_n.n3882 0.002
R57799 vp_n.n3873 vp_n.n3872 0.002
R57800 vp_n.n3863 vp_n.n3862 0.002
R57801 vp_n.n3853 vp_n.n3852 0.002
R57802 vp_n.n3843 vp_n.n3842 0.002
R57803 vp_n.n3833 vp_n.n3832 0.002
R57804 vp_n.n3823 vp_n.n3822 0.002
R57805 vp_n.n3813 vp_n.n3812 0.002
R57806 vp_n.n3803 vp_n.n3802 0.002
R57807 vp_n.n3793 vp_n.n3792 0.002
R57808 vp_n.n3783 vp_n.n3782 0.002
R57809 vp_n.n3773 vp_n.n3772 0.002
R57810 vp_n.n3763 vp_n.n3762 0.002
R57811 vp_n.n3753 vp_n.n3752 0.002
R57812 vp_n.n3743 vp_n.n3742 0.002
R57813 vp_n.n3733 vp_n.n3732 0.002
R57814 vp_n.n3723 vp_n.n3722 0.002
R57815 vp_n.n3713 vp_n.n3712 0.002
R57816 vp_n.n3703 vp_n.n3702 0.002
R57817 vp_n.n3693 vp_n.n3692 0.002
R57818 vp_n.n3683 vp_n.n3682 0.002
R57819 vp_n.n3673 vp_n.n3672 0.002
R57820 vp_n.n3663 vp_n.n3662 0.002
R57821 vp_n.n3653 vp_n.n3652 0.002
R57822 vp_n.n3643 vp_n.n3642 0.002
R57823 vp_n.n3633 vp_n.n3632 0.002
R57824 vp_n.n3623 vp_n.n3622 0.002
R57825 vp_n.n3613 vp_n.n3612 0.002
R57826 vp_n.n3603 vp_n.n3602 0.002
R57827 vp_n.n3593 vp_n.n3592 0.002
R57828 vp_n.n3583 vp_n.n3582 0.002
R57829 vp_n.n3573 vp_n.n3572 0.002
R57830 vp_n.n3563 vp_n.n3562 0.002
R57831 vp_n.n3553 vp_n.n3552 0.002
R57832 vp_n.n3543 vp_n.n3542 0.002
R57833 vp_n.n3533 vp_n.n3532 0.002
R57834 vp_n.n3523 vp_n.n3522 0.002
R57835 vp_n.n3513 vp_n.n3512 0.002
R57836 vp_n.n3503 vp_n.n3502 0.002
R57837 vp_n.n3493 vp_n.n3492 0.002
R57838 vp_n.n3483 vp_n.n3482 0.002
R57839 vp_n.n3473 vp_n.n3472 0.002
R57840 vp_n.n3463 vp_n.n3462 0.002
R57841 vp_n.n3453 vp_n.n3452 0.002
R57842 vp_n.n3443 vp_n.n3442 0.002
R57843 vp_n.n3433 vp_n.n3432 0.002
R57844 vp_n.n3423 vp_n.n3422 0.002
R57845 vp_n.n3413 vp_n.n3412 0.002
R57846 vp_n.n3403 vp_n.n3402 0.002
R57847 vp_n.n3393 vp_n.n3392 0.002
R57848 vp_n.n3383 vp_n.n3382 0.002
R57849 vp_n.n3373 vp_n.n3372 0.002
R57850 vp_n.n3363 vp_n.n3362 0.002
R57851 vp_n.n3353 vp_n.n3352 0.002
R57852 vp_n.n3343 vp_n.n3342 0.002
R57853 vp_n.n3333 vp_n.n3332 0.002
R57854 vp_n.n3323 vp_n.n3322 0.002
R57855 vp_n.n3313 vp_n.n3312 0.002
R57856 vp_n.n3303 vp_n.n3302 0.002
R57857 vp_n.n3293 vp_n.n3292 0.002
R57858 vp_n.n3283 vp_n.n3282 0.002
R57859 vp_n.n3273 vp_n.n3272 0.002
R57860 vp_n.n3263 vp_n.n3262 0.002
R57861 vp_n.n3253 vp_n.n3252 0.002
R57862 vp_n.n3243 vp_n.n3242 0.002
R57863 vp_n.n3233 vp_n.n3232 0.002
R57864 vp_n.n3223 vp_n.n3222 0.002
R57865 vp_n.n3213 vp_n.n3212 0.002
R57866 vss.n3195 vss.n3193 109.642
R57867 vss.n3187 vss.n3185 109.642
R57868 vss.n2408 vss.n2406 100.602
R57869 vss.n2400 vss.n2398 100.602
R57870 vss.n3149 vss.n3146 69.611
R57871 vss.n3149 vss.n3148 69.611
R57872 vss.n3164 vss.n3163 69.611
R57873 vss.n3164 vss.n3161 69.611
R57874 vss.n3107 vss.n3104 69.611
R57875 vss.n3107 vss.n3106 69.611
R57876 vss.n3122 vss.n3121 69.611
R57877 vss.n3122 vss.n3119 69.611
R57878 vss.n3065 vss.n3062 69.611
R57879 vss.n3065 vss.n3064 69.611
R57880 vss.n3080 vss.n3079 69.611
R57881 vss.n3080 vss.n3077 69.611
R57882 vss.n3023 vss.n3020 69.611
R57883 vss.n3023 vss.n3022 69.611
R57884 vss.n3038 vss.n3037 69.611
R57885 vss.n3038 vss.n3035 69.611
R57886 vss.n2981 vss.n2978 69.611
R57887 vss.n2981 vss.n2980 69.611
R57888 vss.n2996 vss.n2995 69.611
R57889 vss.n2996 vss.n2993 69.611
R57890 vss.n2939 vss.n2936 69.611
R57891 vss.n2939 vss.n2938 69.611
R57892 vss.n2954 vss.n2953 69.611
R57893 vss.n2954 vss.n2951 69.611
R57894 vss.n2897 vss.n2894 69.611
R57895 vss.n2897 vss.n2896 69.611
R57896 vss.n2912 vss.n2911 69.611
R57897 vss.n2912 vss.n2909 69.611
R57898 vss.n2855 vss.n2852 69.611
R57899 vss.n2855 vss.n2854 69.611
R57900 vss.n2870 vss.n2869 69.611
R57901 vss.n2870 vss.n2867 69.611
R57902 vss.n2813 vss.n2810 69.611
R57903 vss.n2813 vss.n2812 69.611
R57904 vss.n2828 vss.n2827 69.611
R57905 vss.n2828 vss.n2825 69.611
R57906 vss.n2771 vss.n2768 69.611
R57907 vss.n2771 vss.n2770 69.611
R57908 vss.n2786 vss.n2785 69.611
R57909 vss.n2786 vss.n2783 69.611
R57910 vss.n2729 vss.n2726 69.611
R57911 vss.n2729 vss.n2728 69.611
R57912 vss.n2744 vss.n2743 69.611
R57913 vss.n2744 vss.n2741 69.611
R57914 vss.n2687 vss.n2684 69.611
R57915 vss.n2687 vss.n2686 69.611
R57916 vss.n2702 vss.n2701 69.611
R57917 vss.n2702 vss.n2699 69.611
R57918 vss.n2645 vss.n2642 69.611
R57919 vss.n2645 vss.n2644 69.611
R57920 vss.n2660 vss.n2659 69.611
R57921 vss.n2660 vss.n2657 69.611
R57922 vss.n2603 vss.n2600 69.611
R57923 vss.n2603 vss.n2602 69.611
R57924 vss.n2618 vss.n2617 69.611
R57925 vss.n2618 vss.n2615 69.611
R57926 vss.n2561 vss.n2558 69.611
R57927 vss.n2561 vss.n2560 69.611
R57928 vss.n2576 vss.n2575 69.611
R57929 vss.n2576 vss.n2573 69.611
R57930 vss.n2519 vss.n2516 69.611
R57931 vss.n2519 vss.n2518 69.611
R57932 vss.n2534 vss.n2533 69.611
R57933 vss.n2534 vss.n2531 69.611
R57934 vss.n2477 vss.n2474 69.611
R57935 vss.n2477 vss.n2476 69.611
R57936 vss.n2492 vss.n2491 69.611
R57937 vss.n2492 vss.n2489 69.611
R57938 vss.n10 vss.n7 69.611
R57939 vss.n10 vss.n9 69.611
R57940 vss.n25 vss.n24 69.611
R57941 vss.n25 vss.n22 69.611
R57942 vss.n52 vss.n49 69.611
R57943 vss.n52 vss.n51 69.611
R57944 vss.n67 vss.n66 69.611
R57945 vss.n67 vss.n64 69.611
R57946 vss.n94 vss.n91 69.611
R57947 vss.n94 vss.n93 69.611
R57948 vss.n109 vss.n108 69.611
R57949 vss.n109 vss.n106 69.611
R57950 vss.n136 vss.n133 69.611
R57951 vss.n136 vss.n135 69.611
R57952 vss.n151 vss.n150 69.611
R57953 vss.n151 vss.n148 69.611
R57954 vss.n178 vss.n175 69.611
R57955 vss.n178 vss.n177 69.611
R57956 vss.n193 vss.n192 69.611
R57957 vss.n193 vss.n190 69.611
R57958 vss.n220 vss.n217 69.611
R57959 vss.n220 vss.n219 69.611
R57960 vss.n235 vss.n234 69.611
R57961 vss.n235 vss.n232 69.611
R57962 vss.n262 vss.n259 69.611
R57963 vss.n262 vss.n261 69.611
R57964 vss.n277 vss.n276 69.611
R57965 vss.n277 vss.n274 69.611
R57966 vss.n304 vss.n301 69.611
R57967 vss.n304 vss.n303 69.611
R57968 vss.n319 vss.n318 69.611
R57969 vss.n319 vss.n316 69.611
R57970 vss.n346 vss.n343 69.611
R57971 vss.n346 vss.n345 69.611
R57972 vss.n361 vss.n360 69.611
R57973 vss.n361 vss.n358 69.611
R57974 vss.n388 vss.n385 69.611
R57975 vss.n388 vss.n387 69.611
R57976 vss.n403 vss.n402 69.611
R57977 vss.n403 vss.n400 69.611
R57978 vss.n430 vss.n427 69.611
R57979 vss.n430 vss.n429 69.611
R57980 vss.n445 vss.n444 69.611
R57981 vss.n445 vss.n442 69.611
R57982 vss.n472 vss.n469 69.611
R57983 vss.n472 vss.n471 69.611
R57984 vss.n487 vss.n486 69.611
R57985 vss.n487 vss.n484 69.611
R57986 vss.n514 vss.n511 69.611
R57987 vss.n514 vss.n513 69.611
R57988 vss.n529 vss.n528 69.611
R57989 vss.n529 vss.n526 69.611
R57990 vss.n556 vss.n553 69.611
R57991 vss.n556 vss.n555 69.611
R57992 vss.n571 vss.n570 69.611
R57993 vss.n571 vss.n568 69.611
R57994 vss.n598 vss.n595 69.611
R57995 vss.n598 vss.n597 69.611
R57996 vss.n613 vss.n612 69.611
R57997 vss.n613 vss.n610 69.611
R57998 vss.n640 vss.n637 69.611
R57999 vss.n640 vss.n639 69.611
R58000 vss.n655 vss.n654 69.611
R58001 vss.n655 vss.n652 69.611
R58002 vss.n682 vss.n679 69.611
R58003 vss.n682 vss.n681 69.611
R58004 vss.n697 vss.n696 69.611
R58005 vss.n697 vss.n694 69.611
R58006 vss.n724 vss.n721 69.611
R58007 vss.n724 vss.n723 69.611
R58008 vss.n739 vss.n738 69.611
R58009 vss.n739 vss.n736 69.611
R58010 vss.n766 vss.n763 69.611
R58011 vss.n766 vss.n765 69.611
R58012 vss.n781 vss.n780 69.611
R58013 vss.n781 vss.n778 69.611
R58014 vss.n808 vss.n805 69.611
R58015 vss.n808 vss.n807 69.611
R58016 vss.n823 vss.n822 69.611
R58017 vss.n823 vss.n820 69.611
R58018 vss.n850 vss.n847 69.611
R58019 vss.n850 vss.n849 69.611
R58020 vss.n865 vss.n864 69.611
R58021 vss.n865 vss.n862 69.611
R58022 vss.n892 vss.n889 69.611
R58023 vss.n892 vss.n891 69.611
R58024 vss.n907 vss.n906 69.611
R58025 vss.n907 vss.n904 69.611
R58026 vss.n934 vss.n931 69.611
R58027 vss.n934 vss.n933 69.611
R58028 vss.n949 vss.n948 69.611
R58029 vss.n949 vss.n946 69.611
R58030 vss.n976 vss.n973 69.611
R58031 vss.n976 vss.n975 69.611
R58032 vss.n991 vss.n990 69.611
R58033 vss.n991 vss.n988 69.611
R58034 vss.n1018 vss.n1015 69.611
R58035 vss.n1018 vss.n1017 69.611
R58036 vss.n1033 vss.n1032 69.611
R58037 vss.n1033 vss.n1030 69.611
R58038 vss.n1060 vss.n1057 69.611
R58039 vss.n1060 vss.n1059 69.611
R58040 vss.n1075 vss.n1074 69.611
R58041 vss.n1075 vss.n1072 69.611
R58042 vss.n1102 vss.n1099 69.611
R58043 vss.n1102 vss.n1101 69.611
R58044 vss.n1117 vss.n1116 69.611
R58045 vss.n1117 vss.n1114 69.611
R58046 vss.n1144 vss.n1141 69.611
R58047 vss.n1144 vss.n1143 69.611
R58048 vss.n1159 vss.n1158 69.611
R58049 vss.n1159 vss.n1156 69.611
R58050 vss.n1186 vss.n1183 69.611
R58051 vss.n1186 vss.n1185 69.611
R58052 vss.n1201 vss.n1200 69.611
R58053 vss.n1201 vss.n1198 69.611
R58054 vss.n1228 vss.n1225 69.611
R58055 vss.n1228 vss.n1227 69.611
R58056 vss.n1243 vss.n1242 69.611
R58057 vss.n1243 vss.n1240 69.611
R58058 vss.n1270 vss.n1267 69.611
R58059 vss.n1270 vss.n1269 69.611
R58060 vss.n1285 vss.n1284 69.611
R58061 vss.n1285 vss.n1282 69.611
R58062 vss.n1312 vss.n1309 69.611
R58063 vss.n1312 vss.n1311 69.611
R58064 vss.n1327 vss.n1326 69.611
R58065 vss.n1327 vss.n1324 69.611
R58066 vss.n1354 vss.n1351 69.611
R58067 vss.n1354 vss.n1353 69.611
R58068 vss.n1369 vss.n1368 69.611
R58069 vss.n1369 vss.n1366 69.611
R58070 vss.n1396 vss.n1393 69.611
R58071 vss.n1396 vss.n1395 69.611
R58072 vss.n1411 vss.n1410 69.611
R58073 vss.n1411 vss.n1408 69.611
R58074 vss.n1438 vss.n1435 69.611
R58075 vss.n1438 vss.n1437 69.611
R58076 vss.n1453 vss.n1452 69.611
R58077 vss.n1453 vss.n1450 69.611
R58078 vss.n1480 vss.n1477 69.611
R58079 vss.n1480 vss.n1479 69.611
R58080 vss.n1495 vss.n1494 69.611
R58081 vss.n1495 vss.n1492 69.611
R58082 vss.n1522 vss.n1519 69.611
R58083 vss.n1522 vss.n1521 69.611
R58084 vss.n1537 vss.n1536 69.611
R58085 vss.n1537 vss.n1534 69.611
R58086 vss.n1564 vss.n1561 69.611
R58087 vss.n1564 vss.n1563 69.611
R58088 vss.n1579 vss.n1578 69.611
R58089 vss.n1579 vss.n1576 69.611
R58090 vss.n1606 vss.n1603 69.611
R58091 vss.n1606 vss.n1605 69.611
R58092 vss.n1621 vss.n1620 69.611
R58093 vss.n1621 vss.n1618 69.611
R58094 vss.n1648 vss.n1645 69.611
R58095 vss.n1648 vss.n1647 69.611
R58096 vss.n1663 vss.n1662 69.611
R58097 vss.n1663 vss.n1660 69.611
R58098 vss.n1690 vss.n1687 69.611
R58099 vss.n1690 vss.n1689 69.611
R58100 vss.n1705 vss.n1704 69.611
R58101 vss.n1705 vss.n1702 69.611
R58102 vss.n1732 vss.n1729 69.611
R58103 vss.n1732 vss.n1731 69.611
R58104 vss.n1747 vss.n1746 69.611
R58105 vss.n1747 vss.n1744 69.611
R58106 vss.n1774 vss.n1771 69.611
R58107 vss.n1774 vss.n1773 69.611
R58108 vss.n1789 vss.n1788 69.611
R58109 vss.n1789 vss.n1786 69.611
R58110 vss.n1816 vss.n1813 69.611
R58111 vss.n1816 vss.n1815 69.611
R58112 vss.n1831 vss.n1830 69.611
R58113 vss.n1831 vss.n1828 69.611
R58114 vss.n1858 vss.n1855 69.611
R58115 vss.n1858 vss.n1857 69.611
R58116 vss.n1873 vss.n1872 69.611
R58117 vss.n1873 vss.n1870 69.611
R58118 vss.n1900 vss.n1897 69.611
R58119 vss.n1900 vss.n1899 69.611
R58120 vss.n1915 vss.n1914 69.611
R58121 vss.n1915 vss.n1912 69.611
R58122 vss.n1942 vss.n1939 69.611
R58123 vss.n1942 vss.n1941 69.611
R58124 vss.n1957 vss.n1956 69.611
R58125 vss.n1957 vss.n1954 69.611
R58126 vss.n1984 vss.n1981 69.611
R58127 vss.n1984 vss.n1983 69.611
R58128 vss.n1999 vss.n1998 69.611
R58129 vss.n1999 vss.n1996 69.611
R58130 vss.n2026 vss.n2023 69.611
R58131 vss.n2026 vss.n2025 69.611
R58132 vss.n2041 vss.n2040 69.611
R58133 vss.n2041 vss.n2038 69.611
R58134 vss.n2068 vss.n2065 69.611
R58135 vss.n2068 vss.n2067 69.611
R58136 vss.n2083 vss.n2082 69.611
R58137 vss.n2083 vss.n2080 69.611
R58138 vss.n2110 vss.n2107 69.611
R58139 vss.n2110 vss.n2109 69.611
R58140 vss.n2125 vss.n2124 69.611
R58141 vss.n2125 vss.n2122 69.611
R58142 vss.n2152 vss.n2149 69.611
R58143 vss.n2152 vss.n2151 69.611
R58144 vss.n2167 vss.n2166 69.611
R58145 vss.n2167 vss.n2164 69.611
R58146 vss.n2194 vss.n2191 69.611
R58147 vss.n2194 vss.n2193 69.611
R58148 vss.n2209 vss.n2208 69.611
R58149 vss.n2209 vss.n2206 69.611
R58150 vss.n2236 vss.n2233 69.611
R58151 vss.n2236 vss.n2235 69.611
R58152 vss.n2251 vss.n2250 69.611
R58153 vss.n2251 vss.n2248 69.611
R58154 vss.n2278 vss.n2275 69.611
R58155 vss.n2278 vss.n2277 69.611
R58156 vss.n2293 vss.n2292 69.611
R58157 vss.n2293 vss.n2290 69.611
R58158 vss.n2320 vss.n2317 69.611
R58159 vss.n2320 vss.n2319 69.611
R58160 vss.n2335 vss.n2334 69.611
R58161 vss.n2335 vss.n2332 69.611
R58162 vss.n2362 vss.n2359 69.611
R58163 vss.n2362 vss.n2361 69.611
R58164 vss.n2377 vss.n2376 69.611
R58165 vss.n2377 vss.n2374 69.611
R58166 vss.n3174 vss.n3173 66.741
R58167 vss.n3174 vss.n3171 66.741
R58168 vss.n3132 vss.n3131 66.741
R58169 vss.n3132 vss.n3129 66.741
R58170 vss.n3090 vss.n3089 66.741
R58171 vss.n3090 vss.n3087 66.741
R58172 vss.n3048 vss.n3047 66.741
R58173 vss.n3048 vss.n3045 66.741
R58174 vss.n3006 vss.n3005 66.741
R58175 vss.n3006 vss.n3003 66.741
R58176 vss.n2964 vss.n2963 66.741
R58177 vss.n2964 vss.n2961 66.741
R58178 vss.n2922 vss.n2921 66.741
R58179 vss.n2922 vss.n2919 66.741
R58180 vss.n2880 vss.n2879 66.741
R58181 vss.n2880 vss.n2877 66.741
R58182 vss.n2838 vss.n2837 66.741
R58183 vss.n2838 vss.n2835 66.741
R58184 vss.n2796 vss.n2795 66.741
R58185 vss.n2796 vss.n2793 66.741
R58186 vss.n2754 vss.n2753 66.741
R58187 vss.n2754 vss.n2751 66.741
R58188 vss.n2712 vss.n2711 66.741
R58189 vss.n2712 vss.n2709 66.741
R58190 vss.n2670 vss.n2669 66.741
R58191 vss.n2670 vss.n2667 66.741
R58192 vss.n2628 vss.n2627 66.741
R58193 vss.n2628 vss.n2625 66.741
R58194 vss.n2586 vss.n2585 66.741
R58195 vss.n2586 vss.n2583 66.741
R58196 vss.n2544 vss.n2543 66.741
R58197 vss.n2544 vss.n2541 66.741
R58198 vss.n2502 vss.n2501 66.741
R58199 vss.n2502 vss.n2499 66.741
R58200 vss.n35 vss.n34 66.741
R58201 vss.n35 vss.n32 66.741
R58202 vss.n77 vss.n76 66.741
R58203 vss.n77 vss.n74 66.741
R58204 vss.n119 vss.n118 66.741
R58205 vss.n119 vss.n116 66.741
R58206 vss.n161 vss.n160 66.741
R58207 vss.n161 vss.n158 66.741
R58208 vss.n203 vss.n202 66.741
R58209 vss.n203 vss.n200 66.741
R58210 vss.n245 vss.n244 66.741
R58211 vss.n245 vss.n242 66.741
R58212 vss.n287 vss.n286 66.741
R58213 vss.n287 vss.n284 66.741
R58214 vss.n329 vss.n328 66.741
R58215 vss.n329 vss.n326 66.741
R58216 vss.n371 vss.n370 66.741
R58217 vss.n371 vss.n368 66.741
R58218 vss.n413 vss.n412 66.741
R58219 vss.n413 vss.n410 66.741
R58220 vss.n455 vss.n454 66.741
R58221 vss.n455 vss.n452 66.741
R58222 vss.n497 vss.n496 66.741
R58223 vss.n497 vss.n494 66.741
R58224 vss.n539 vss.n538 66.741
R58225 vss.n539 vss.n536 66.741
R58226 vss.n581 vss.n580 66.741
R58227 vss.n581 vss.n578 66.741
R58228 vss.n623 vss.n622 66.741
R58229 vss.n623 vss.n620 66.741
R58230 vss.n665 vss.n664 66.741
R58231 vss.n665 vss.n662 66.741
R58232 vss.n707 vss.n706 66.741
R58233 vss.n707 vss.n704 66.741
R58234 vss.n749 vss.n748 66.741
R58235 vss.n749 vss.n746 66.741
R58236 vss.n791 vss.n790 66.741
R58237 vss.n791 vss.n788 66.741
R58238 vss.n833 vss.n832 66.741
R58239 vss.n833 vss.n830 66.741
R58240 vss.n875 vss.n874 66.741
R58241 vss.n875 vss.n872 66.741
R58242 vss.n917 vss.n916 66.741
R58243 vss.n917 vss.n914 66.741
R58244 vss.n959 vss.n958 66.741
R58245 vss.n959 vss.n956 66.741
R58246 vss.n1001 vss.n1000 66.741
R58247 vss.n1001 vss.n998 66.741
R58248 vss.n1043 vss.n1042 66.741
R58249 vss.n1043 vss.n1040 66.741
R58250 vss.n1085 vss.n1084 66.741
R58251 vss.n1085 vss.n1082 66.741
R58252 vss.n1127 vss.n1126 66.741
R58253 vss.n1127 vss.n1124 66.741
R58254 vss.n1169 vss.n1168 66.741
R58255 vss.n1169 vss.n1166 66.741
R58256 vss.n1211 vss.n1210 66.741
R58257 vss.n1211 vss.n1208 66.741
R58258 vss.n1253 vss.n1252 66.741
R58259 vss.n1253 vss.n1250 66.741
R58260 vss.n1295 vss.n1294 66.741
R58261 vss.n1295 vss.n1292 66.741
R58262 vss.n1337 vss.n1336 66.741
R58263 vss.n1337 vss.n1334 66.741
R58264 vss.n1379 vss.n1378 66.741
R58265 vss.n1379 vss.n1376 66.741
R58266 vss.n1421 vss.n1420 66.741
R58267 vss.n1421 vss.n1418 66.741
R58268 vss.n1463 vss.n1462 66.741
R58269 vss.n1463 vss.n1460 66.741
R58270 vss.n1505 vss.n1504 66.741
R58271 vss.n1505 vss.n1502 66.741
R58272 vss.n1547 vss.n1546 66.741
R58273 vss.n1547 vss.n1544 66.741
R58274 vss.n1589 vss.n1588 66.741
R58275 vss.n1589 vss.n1586 66.741
R58276 vss.n1631 vss.n1630 66.741
R58277 vss.n1631 vss.n1628 66.741
R58278 vss.n1673 vss.n1672 66.741
R58279 vss.n1673 vss.n1670 66.741
R58280 vss.n1715 vss.n1714 66.741
R58281 vss.n1715 vss.n1712 66.741
R58282 vss.n1757 vss.n1756 66.741
R58283 vss.n1757 vss.n1754 66.741
R58284 vss.n1799 vss.n1798 66.741
R58285 vss.n1799 vss.n1796 66.741
R58286 vss.n1841 vss.n1840 66.741
R58287 vss.n1841 vss.n1838 66.741
R58288 vss.n1883 vss.n1882 66.741
R58289 vss.n1883 vss.n1880 66.741
R58290 vss.n1925 vss.n1924 66.741
R58291 vss.n1925 vss.n1922 66.741
R58292 vss.n1967 vss.n1966 66.741
R58293 vss.n1967 vss.n1964 66.741
R58294 vss.n2009 vss.n2008 66.741
R58295 vss.n2009 vss.n2006 66.741
R58296 vss.n2051 vss.n2050 66.741
R58297 vss.n2051 vss.n2048 66.741
R58298 vss.n2093 vss.n2092 66.741
R58299 vss.n2093 vss.n2090 66.741
R58300 vss.n2135 vss.n2134 66.741
R58301 vss.n2135 vss.n2132 66.741
R58302 vss.n2177 vss.n2176 66.741
R58303 vss.n2177 vss.n2174 66.741
R58304 vss.n2219 vss.n2218 66.741
R58305 vss.n2219 vss.n2216 66.741
R58306 vss.n2261 vss.n2260 66.741
R58307 vss.n2261 vss.n2258 66.741
R58308 vss.n2303 vss.n2302 66.741
R58309 vss.n2303 vss.n2300 66.741
R58310 vss.n2345 vss.n2344 66.741
R58311 vss.n2345 vss.n2342 66.741
R58312 vss.n2387 vss.n2386 66.741
R58313 vss.n2387 vss.n2384 66.741
R58314 vss.n3142 vss.n3140 30.859
R58315 vss.n3142 vss.n3141 30.859
R58316 vss.n3100 vss.n3098 30.859
R58317 vss.n3100 vss.n3099 30.859
R58318 vss.n3058 vss.n3056 30.859
R58319 vss.n3058 vss.n3057 30.859
R58320 vss.n3016 vss.n3014 30.859
R58321 vss.n3016 vss.n3015 30.859
R58322 vss.n2974 vss.n2972 30.859
R58323 vss.n2974 vss.n2973 30.859
R58324 vss.n2932 vss.n2930 30.859
R58325 vss.n2932 vss.n2931 30.859
R58326 vss.n2890 vss.n2888 30.859
R58327 vss.n2890 vss.n2889 30.859
R58328 vss.n2848 vss.n2846 30.859
R58329 vss.n2848 vss.n2847 30.859
R58330 vss.n2806 vss.n2804 30.859
R58331 vss.n2806 vss.n2805 30.859
R58332 vss.n2764 vss.n2762 30.859
R58333 vss.n2764 vss.n2763 30.859
R58334 vss.n2722 vss.n2720 30.859
R58335 vss.n2722 vss.n2721 30.859
R58336 vss.n2680 vss.n2678 30.859
R58337 vss.n2680 vss.n2679 30.859
R58338 vss.n2638 vss.n2636 30.859
R58339 vss.n2638 vss.n2637 30.859
R58340 vss.n2596 vss.n2594 30.859
R58341 vss.n2596 vss.n2595 30.859
R58342 vss.n2554 vss.n2552 30.859
R58343 vss.n2554 vss.n2553 30.859
R58344 vss.n2512 vss.n2510 30.859
R58345 vss.n2512 vss.n2511 30.859
R58346 vss.n2470 vss.n2468 30.859
R58347 vss.n2470 vss.n2469 30.859
R58348 vss.n3 vss.n1 30.859
R58349 vss.n3 vss.n2 30.859
R58350 vss.n45 vss.n43 30.859
R58351 vss.n45 vss.n44 30.859
R58352 vss.n87 vss.n85 30.859
R58353 vss.n87 vss.n86 30.859
R58354 vss.n129 vss.n127 30.859
R58355 vss.n129 vss.n128 30.859
R58356 vss.n171 vss.n169 30.859
R58357 vss.n171 vss.n170 30.859
R58358 vss.n213 vss.n211 30.859
R58359 vss.n213 vss.n212 30.859
R58360 vss.n255 vss.n253 30.859
R58361 vss.n255 vss.n254 30.859
R58362 vss.n297 vss.n295 30.859
R58363 vss.n297 vss.n296 30.859
R58364 vss.n339 vss.n337 30.859
R58365 vss.n339 vss.n338 30.859
R58366 vss.n381 vss.n379 30.859
R58367 vss.n381 vss.n380 30.859
R58368 vss.n423 vss.n421 30.859
R58369 vss.n423 vss.n422 30.859
R58370 vss.n465 vss.n463 30.859
R58371 vss.n465 vss.n464 30.859
R58372 vss.n507 vss.n505 30.859
R58373 vss.n507 vss.n506 30.859
R58374 vss.n549 vss.n547 30.859
R58375 vss.n549 vss.n548 30.859
R58376 vss.n591 vss.n589 30.859
R58377 vss.n591 vss.n590 30.859
R58378 vss.n633 vss.n631 30.859
R58379 vss.n633 vss.n632 30.859
R58380 vss.n675 vss.n673 30.859
R58381 vss.n675 vss.n674 30.859
R58382 vss.n717 vss.n715 30.859
R58383 vss.n717 vss.n716 30.859
R58384 vss.n759 vss.n757 30.859
R58385 vss.n759 vss.n758 30.859
R58386 vss.n801 vss.n799 30.859
R58387 vss.n801 vss.n800 30.859
R58388 vss.n843 vss.n841 30.859
R58389 vss.n843 vss.n842 30.859
R58390 vss.n885 vss.n883 30.859
R58391 vss.n885 vss.n884 30.859
R58392 vss.n927 vss.n925 30.859
R58393 vss.n927 vss.n926 30.859
R58394 vss.n969 vss.n967 30.859
R58395 vss.n969 vss.n968 30.859
R58396 vss.n1011 vss.n1009 30.859
R58397 vss.n1011 vss.n1010 30.859
R58398 vss.n1053 vss.n1051 30.859
R58399 vss.n1053 vss.n1052 30.859
R58400 vss.n1095 vss.n1093 30.859
R58401 vss.n1095 vss.n1094 30.859
R58402 vss.n1137 vss.n1135 30.859
R58403 vss.n1137 vss.n1136 30.859
R58404 vss.n1179 vss.n1177 30.859
R58405 vss.n1179 vss.n1178 30.859
R58406 vss.n1221 vss.n1219 30.859
R58407 vss.n1221 vss.n1220 30.859
R58408 vss.n1263 vss.n1261 30.859
R58409 vss.n1263 vss.n1262 30.859
R58410 vss.n1305 vss.n1303 30.859
R58411 vss.n1305 vss.n1304 30.859
R58412 vss.n1347 vss.n1345 30.859
R58413 vss.n1347 vss.n1346 30.859
R58414 vss.n1389 vss.n1387 30.859
R58415 vss.n1389 vss.n1388 30.859
R58416 vss.n1431 vss.n1429 30.859
R58417 vss.n1431 vss.n1430 30.859
R58418 vss.n1473 vss.n1471 30.859
R58419 vss.n1473 vss.n1472 30.859
R58420 vss.n1515 vss.n1513 30.859
R58421 vss.n1515 vss.n1514 30.859
R58422 vss.n1557 vss.n1555 30.859
R58423 vss.n1557 vss.n1556 30.859
R58424 vss.n1599 vss.n1597 30.859
R58425 vss.n1599 vss.n1598 30.859
R58426 vss.n1641 vss.n1639 30.859
R58427 vss.n1641 vss.n1640 30.859
R58428 vss.n1683 vss.n1681 30.859
R58429 vss.n1683 vss.n1682 30.859
R58430 vss.n1725 vss.n1723 30.859
R58431 vss.n1725 vss.n1724 30.859
R58432 vss.n1767 vss.n1765 30.859
R58433 vss.n1767 vss.n1766 30.859
R58434 vss.n1809 vss.n1807 30.859
R58435 vss.n1809 vss.n1808 30.859
R58436 vss.n1851 vss.n1849 30.859
R58437 vss.n1851 vss.n1850 30.859
R58438 vss.n1893 vss.n1891 30.859
R58439 vss.n1893 vss.n1892 30.859
R58440 vss.n1935 vss.n1933 30.859
R58441 vss.n1935 vss.n1934 30.859
R58442 vss.n1977 vss.n1975 30.859
R58443 vss.n1977 vss.n1976 30.859
R58444 vss.n2019 vss.n2017 30.859
R58445 vss.n2019 vss.n2018 30.859
R58446 vss.n2061 vss.n2059 30.859
R58447 vss.n2061 vss.n2060 30.859
R58448 vss.n2103 vss.n2101 30.859
R58449 vss.n2103 vss.n2102 30.859
R58450 vss.n2145 vss.n2143 30.859
R58451 vss.n2145 vss.n2144 30.859
R58452 vss.n2187 vss.n2185 30.859
R58453 vss.n2187 vss.n2186 30.859
R58454 vss.n2229 vss.n2227 30.859
R58455 vss.n2229 vss.n2228 30.859
R58456 vss.n2271 vss.n2269 30.859
R58457 vss.n2271 vss.n2270 30.859
R58458 vss.n2313 vss.n2311 30.859
R58459 vss.n2313 vss.n2312 30.859
R58460 vss.n2355 vss.n2353 30.859
R58461 vss.n2355 vss.n2354 30.859
R58462 vss.n3154 vss.n3152 27.63
R58463 vss.n3154 vss.n3153 27.63
R58464 vss.n3112 vss.n3110 27.63
R58465 vss.n3112 vss.n3111 27.63
R58466 vss.n3070 vss.n3068 27.63
R58467 vss.n3070 vss.n3069 27.63
R58468 vss.n3028 vss.n3026 27.63
R58469 vss.n3028 vss.n3027 27.63
R58470 vss.n2986 vss.n2984 27.63
R58471 vss.n2986 vss.n2985 27.63
R58472 vss.n2944 vss.n2942 27.63
R58473 vss.n2944 vss.n2943 27.63
R58474 vss.n2902 vss.n2900 27.63
R58475 vss.n2902 vss.n2901 27.63
R58476 vss.n2860 vss.n2858 27.63
R58477 vss.n2860 vss.n2859 27.63
R58478 vss.n2818 vss.n2816 27.63
R58479 vss.n2818 vss.n2817 27.63
R58480 vss.n2776 vss.n2774 27.63
R58481 vss.n2776 vss.n2775 27.63
R58482 vss.n2734 vss.n2732 27.63
R58483 vss.n2734 vss.n2733 27.63
R58484 vss.n2692 vss.n2690 27.63
R58485 vss.n2692 vss.n2691 27.63
R58486 vss.n2650 vss.n2648 27.63
R58487 vss.n2650 vss.n2649 27.63
R58488 vss.n2608 vss.n2606 27.63
R58489 vss.n2608 vss.n2607 27.63
R58490 vss.n2566 vss.n2564 27.63
R58491 vss.n2566 vss.n2565 27.63
R58492 vss.n2524 vss.n2522 27.63
R58493 vss.n2524 vss.n2523 27.63
R58494 vss.n2482 vss.n2480 27.63
R58495 vss.n2482 vss.n2481 27.63
R58496 vss.n15 vss.n13 27.63
R58497 vss.n15 vss.n14 27.63
R58498 vss.n57 vss.n55 27.63
R58499 vss.n57 vss.n56 27.63
R58500 vss.n99 vss.n97 27.63
R58501 vss.n99 vss.n98 27.63
R58502 vss.n141 vss.n139 27.63
R58503 vss.n141 vss.n140 27.63
R58504 vss.n183 vss.n181 27.63
R58505 vss.n183 vss.n182 27.63
R58506 vss.n225 vss.n223 27.63
R58507 vss.n225 vss.n224 27.63
R58508 vss.n267 vss.n265 27.63
R58509 vss.n267 vss.n266 27.63
R58510 vss.n309 vss.n307 27.63
R58511 vss.n309 vss.n308 27.63
R58512 vss.n351 vss.n349 27.63
R58513 vss.n351 vss.n350 27.63
R58514 vss.n393 vss.n391 27.63
R58515 vss.n393 vss.n392 27.63
R58516 vss.n435 vss.n433 27.63
R58517 vss.n435 vss.n434 27.63
R58518 vss.n477 vss.n475 27.63
R58519 vss.n477 vss.n476 27.63
R58520 vss.n519 vss.n517 27.63
R58521 vss.n519 vss.n518 27.63
R58522 vss.n561 vss.n559 27.63
R58523 vss.n561 vss.n560 27.63
R58524 vss.n603 vss.n601 27.63
R58525 vss.n603 vss.n602 27.63
R58526 vss.n645 vss.n643 27.63
R58527 vss.n645 vss.n644 27.63
R58528 vss.n687 vss.n685 27.63
R58529 vss.n687 vss.n686 27.63
R58530 vss.n729 vss.n727 27.63
R58531 vss.n729 vss.n728 27.63
R58532 vss.n771 vss.n769 27.63
R58533 vss.n771 vss.n770 27.63
R58534 vss.n813 vss.n811 27.63
R58535 vss.n813 vss.n812 27.63
R58536 vss.n855 vss.n853 27.63
R58537 vss.n855 vss.n854 27.63
R58538 vss.n897 vss.n895 27.63
R58539 vss.n897 vss.n896 27.63
R58540 vss.n939 vss.n937 27.63
R58541 vss.n939 vss.n938 27.63
R58542 vss.n981 vss.n979 27.63
R58543 vss.n981 vss.n980 27.63
R58544 vss.n1023 vss.n1021 27.63
R58545 vss.n1023 vss.n1022 27.63
R58546 vss.n1065 vss.n1063 27.63
R58547 vss.n1065 vss.n1064 27.63
R58548 vss.n1107 vss.n1105 27.63
R58549 vss.n1107 vss.n1106 27.63
R58550 vss.n1149 vss.n1147 27.63
R58551 vss.n1149 vss.n1148 27.63
R58552 vss.n1191 vss.n1189 27.63
R58553 vss.n1191 vss.n1190 27.63
R58554 vss.n1233 vss.n1231 27.63
R58555 vss.n1233 vss.n1232 27.63
R58556 vss.n1275 vss.n1273 27.63
R58557 vss.n1275 vss.n1274 27.63
R58558 vss.n1317 vss.n1315 27.63
R58559 vss.n1317 vss.n1316 27.63
R58560 vss.n1359 vss.n1357 27.63
R58561 vss.n1359 vss.n1358 27.63
R58562 vss.n1401 vss.n1399 27.63
R58563 vss.n1401 vss.n1400 27.63
R58564 vss.n1443 vss.n1441 27.63
R58565 vss.n1443 vss.n1442 27.63
R58566 vss.n1485 vss.n1483 27.63
R58567 vss.n1485 vss.n1484 27.63
R58568 vss.n1527 vss.n1525 27.63
R58569 vss.n1527 vss.n1526 27.63
R58570 vss.n1569 vss.n1567 27.63
R58571 vss.n1569 vss.n1568 27.63
R58572 vss.n1611 vss.n1609 27.63
R58573 vss.n1611 vss.n1610 27.63
R58574 vss.n1653 vss.n1651 27.63
R58575 vss.n1653 vss.n1652 27.63
R58576 vss.n1695 vss.n1693 27.63
R58577 vss.n1695 vss.n1694 27.63
R58578 vss.n1737 vss.n1735 27.63
R58579 vss.n1737 vss.n1736 27.63
R58580 vss.n1779 vss.n1777 27.63
R58581 vss.n1779 vss.n1778 27.63
R58582 vss.n1821 vss.n1819 27.63
R58583 vss.n1821 vss.n1820 27.63
R58584 vss.n1863 vss.n1861 27.63
R58585 vss.n1863 vss.n1862 27.63
R58586 vss.n1905 vss.n1903 27.63
R58587 vss.n1905 vss.n1904 27.63
R58588 vss.n1947 vss.n1945 27.63
R58589 vss.n1947 vss.n1946 27.63
R58590 vss.n1989 vss.n1987 27.63
R58591 vss.n1989 vss.n1988 27.63
R58592 vss.n2031 vss.n2029 27.63
R58593 vss.n2031 vss.n2030 27.63
R58594 vss.n2073 vss.n2071 27.63
R58595 vss.n2073 vss.n2072 27.63
R58596 vss.n2115 vss.n2113 27.63
R58597 vss.n2115 vss.n2114 27.63
R58598 vss.n2157 vss.n2155 27.63
R58599 vss.n2157 vss.n2156 27.63
R58600 vss.n2199 vss.n2197 27.63
R58601 vss.n2199 vss.n2198 27.63
R58602 vss.n2241 vss.n2239 27.63
R58603 vss.n2241 vss.n2240 27.63
R58604 vss.n2283 vss.n2281 27.63
R58605 vss.n2283 vss.n2282 27.63
R58606 vss.n2325 vss.n2323 27.63
R58607 vss.n2325 vss.n2324 27.63
R58608 vss.n2367 vss.n2365 27.63
R58609 vss.n2367 vss.n2366 27.63
R58610 vss.n3178 vss.n3174 19.409
R58611 vss.n3178 vss.n3176 19.409
R58612 vss.n3168 vss.n3164 19.409
R58613 vss.n3168 vss.n3166 19.409
R58614 vss.n3158 vss.n3154 19.409
R58615 vss.n3158 vss.n3156 19.409
R58616 vss.n3150 vss.n3149 19.409
R58617 vss.n3150 vss.n3142 19.409
R58618 vss.n3136 vss.n3132 19.409
R58619 vss.n3136 vss.n3134 19.409
R58620 vss.n3126 vss.n3122 19.409
R58621 vss.n3126 vss.n3124 19.409
R58622 vss.n3116 vss.n3112 19.409
R58623 vss.n3116 vss.n3114 19.409
R58624 vss.n3108 vss.n3107 19.409
R58625 vss.n3108 vss.n3100 19.409
R58626 vss.n3094 vss.n3090 19.409
R58627 vss.n3094 vss.n3092 19.409
R58628 vss.n3084 vss.n3080 19.409
R58629 vss.n3084 vss.n3082 19.409
R58630 vss.n3074 vss.n3070 19.409
R58631 vss.n3074 vss.n3072 19.409
R58632 vss.n3066 vss.n3065 19.409
R58633 vss.n3066 vss.n3058 19.409
R58634 vss.n3052 vss.n3048 19.409
R58635 vss.n3052 vss.n3050 19.409
R58636 vss.n3042 vss.n3038 19.409
R58637 vss.n3042 vss.n3040 19.409
R58638 vss.n3032 vss.n3028 19.409
R58639 vss.n3032 vss.n3030 19.409
R58640 vss.n3024 vss.n3023 19.409
R58641 vss.n3024 vss.n3016 19.409
R58642 vss.n3010 vss.n3006 19.409
R58643 vss.n3010 vss.n3008 19.409
R58644 vss.n3000 vss.n2996 19.409
R58645 vss.n3000 vss.n2998 19.409
R58646 vss.n2990 vss.n2986 19.409
R58647 vss.n2990 vss.n2988 19.409
R58648 vss.n2982 vss.n2981 19.409
R58649 vss.n2982 vss.n2974 19.409
R58650 vss.n2968 vss.n2964 19.409
R58651 vss.n2968 vss.n2966 19.409
R58652 vss.n2958 vss.n2954 19.409
R58653 vss.n2958 vss.n2956 19.409
R58654 vss.n2948 vss.n2944 19.409
R58655 vss.n2948 vss.n2946 19.409
R58656 vss.n2940 vss.n2939 19.409
R58657 vss.n2940 vss.n2932 19.409
R58658 vss.n2926 vss.n2922 19.409
R58659 vss.n2926 vss.n2924 19.409
R58660 vss.n2916 vss.n2912 19.409
R58661 vss.n2916 vss.n2914 19.409
R58662 vss.n2906 vss.n2902 19.409
R58663 vss.n2906 vss.n2904 19.409
R58664 vss.n2898 vss.n2897 19.409
R58665 vss.n2898 vss.n2890 19.409
R58666 vss.n2884 vss.n2880 19.409
R58667 vss.n2884 vss.n2882 19.409
R58668 vss.n2874 vss.n2870 19.409
R58669 vss.n2874 vss.n2872 19.409
R58670 vss.n2864 vss.n2860 19.409
R58671 vss.n2864 vss.n2862 19.409
R58672 vss.n2856 vss.n2855 19.409
R58673 vss.n2856 vss.n2848 19.409
R58674 vss.n2842 vss.n2838 19.409
R58675 vss.n2842 vss.n2840 19.409
R58676 vss.n2832 vss.n2828 19.409
R58677 vss.n2832 vss.n2830 19.409
R58678 vss.n2822 vss.n2818 19.409
R58679 vss.n2822 vss.n2820 19.409
R58680 vss.n2814 vss.n2813 19.409
R58681 vss.n2814 vss.n2806 19.409
R58682 vss.n2800 vss.n2796 19.409
R58683 vss.n2800 vss.n2798 19.409
R58684 vss.n2790 vss.n2786 19.409
R58685 vss.n2790 vss.n2788 19.409
R58686 vss.n2780 vss.n2776 19.409
R58687 vss.n2780 vss.n2778 19.409
R58688 vss.n2772 vss.n2771 19.409
R58689 vss.n2772 vss.n2764 19.409
R58690 vss.n2758 vss.n2754 19.409
R58691 vss.n2758 vss.n2756 19.409
R58692 vss.n2748 vss.n2744 19.409
R58693 vss.n2748 vss.n2746 19.409
R58694 vss.n2738 vss.n2734 19.409
R58695 vss.n2738 vss.n2736 19.409
R58696 vss.n2730 vss.n2729 19.409
R58697 vss.n2730 vss.n2722 19.409
R58698 vss.n2716 vss.n2712 19.409
R58699 vss.n2716 vss.n2714 19.409
R58700 vss.n2706 vss.n2702 19.409
R58701 vss.n2706 vss.n2704 19.409
R58702 vss.n2696 vss.n2692 19.409
R58703 vss.n2696 vss.n2694 19.409
R58704 vss.n2688 vss.n2687 19.409
R58705 vss.n2688 vss.n2680 19.409
R58706 vss.n2674 vss.n2670 19.409
R58707 vss.n2674 vss.n2672 19.409
R58708 vss.n2664 vss.n2660 19.409
R58709 vss.n2664 vss.n2662 19.409
R58710 vss.n2654 vss.n2650 19.409
R58711 vss.n2654 vss.n2652 19.409
R58712 vss.n2646 vss.n2645 19.409
R58713 vss.n2646 vss.n2638 19.409
R58714 vss.n2632 vss.n2628 19.409
R58715 vss.n2632 vss.n2630 19.409
R58716 vss.n2622 vss.n2618 19.409
R58717 vss.n2622 vss.n2620 19.409
R58718 vss.n2612 vss.n2608 19.409
R58719 vss.n2612 vss.n2610 19.409
R58720 vss.n2604 vss.n2603 19.409
R58721 vss.n2604 vss.n2596 19.409
R58722 vss.n2590 vss.n2586 19.409
R58723 vss.n2590 vss.n2588 19.409
R58724 vss.n2580 vss.n2576 19.409
R58725 vss.n2580 vss.n2578 19.409
R58726 vss.n2570 vss.n2566 19.409
R58727 vss.n2570 vss.n2568 19.409
R58728 vss.n2562 vss.n2561 19.409
R58729 vss.n2562 vss.n2554 19.409
R58730 vss.n2548 vss.n2544 19.409
R58731 vss.n2548 vss.n2546 19.409
R58732 vss.n2538 vss.n2534 19.409
R58733 vss.n2538 vss.n2536 19.409
R58734 vss.n2528 vss.n2524 19.409
R58735 vss.n2528 vss.n2526 19.409
R58736 vss.n2520 vss.n2519 19.409
R58737 vss.n2520 vss.n2512 19.409
R58738 vss.n2506 vss.n2502 19.409
R58739 vss.n2506 vss.n2504 19.409
R58740 vss.n2496 vss.n2492 19.409
R58741 vss.n2496 vss.n2494 19.409
R58742 vss.n2486 vss.n2482 19.409
R58743 vss.n2486 vss.n2484 19.409
R58744 vss.n2478 vss.n2477 19.409
R58745 vss.n2478 vss.n2470 19.409
R58746 vss.n39 vss.n35 19.409
R58747 vss.n39 vss.n37 19.409
R58748 vss.n29 vss.n25 19.409
R58749 vss.n29 vss.n27 19.409
R58750 vss.n19 vss.n15 19.409
R58751 vss.n19 vss.n17 19.409
R58752 vss.n11 vss.n10 19.409
R58753 vss.n11 vss.n3 19.409
R58754 vss.n81 vss.n77 19.409
R58755 vss.n81 vss.n79 19.409
R58756 vss.n71 vss.n67 19.409
R58757 vss.n71 vss.n69 19.409
R58758 vss.n61 vss.n57 19.409
R58759 vss.n61 vss.n59 19.409
R58760 vss.n53 vss.n52 19.409
R58761 vss.n53 vss.n45 19.409
R58762 vss.n123 vss.n119 19.409
R58763 vss.n123 vss.n121 19.409
R58764 vss.n113 vss.n109 19.409
R58765 vss.n113 vss.n111 19.409
R58766 vss.n103 vss.n99 19.409
R58767 vss.n103 vss.n101 19.409
R58768 vss.n95 vss.n94 19.409
R58769 vss.n95 vss.n87 19.409
R58770 vss.n165 vss.n161 19.409
R58771 vss.n165 vss.n163 19.409
R58772 vss.n155 vss.n151 19.409
R58773 vss.n155 vss.n153 19.409
R58774 vss.n145 vss.n141 19.409
R58775 vss.n145 vss.n143 19.409
R58776 vss.n137 vss.n136 19.409
R58777 vss.n137 vss.n129 19.409
R58778 vss.n207 vss.n203 19.409
R58779 vss.n207 vss.n205 19.409
R58780 vss.n197 vss.n193 19.409
R58781 vss.n197 vss.n195 19.409
R58782 vss.n187 vss.n183 19.409
R58783 vss.n187 vss.n185 19.409
R58784 vss.n179 vss.n178 19.409
R58785 vss.n179 vss.n171 19.409
R58786 vss.n249 vss.n245 19.409
R58787 vss.n249 vss.n247 19.409
R58788 vss.n239 vss.n235 19.409
R58789 vss.n239 vss.n237 19.409
R58790 vss.n229 vss.n225 19.409
R58791 vss.n229 vss.n227 19.409
R58792 vss.n221 vss.n220 19.409
R58793 vss.n221 vss.n213 19.409
R58794 vss.n291 vss.n287 19.409
R58795 vss.n291 vss.n289 19.409
R58796 vss.n281 vss.n277 19.409
R58797 vss.n281 vss.n279 19.409
R58798 vss.n271 vss.n267 19.409
R58799 vss.n271 vss.n269 19.409
R58800 vss.n263 vss.n262 19.409
R58801 vss.n263 vss.n255 19.409
R58802 vss.n333 vss.n329 19.409
R58803 vss.n333 vss.n331 19.409
R58804 vss.n323 vss.n319 19.409
R58805 vss.n323 vss.n321 19.409
R58806 vss.n313 vss.n309 19.409
R58807 vss.n313 vss.n311 19.409
R58808 vss.n305 vss.n304 19.409
R58809 vss.n305 vss.n297 19.409
R58810 vss.n375 vss.n371 19.409
R58811 vss.n375 vss.n373 19.409
R58812 vss.n365 vss.n361 19.409
R58813 vss.n365 vss.n363 19.409
R58814 vss.n355 vss.n351 19.409
R58815 vss.n355 vss.n353 19.409
R58816 vss.n347 vss.n346 19.409
R58817 vss.n347 vss.n339 19.409
R58818 vss.n417 vss.n413 19.409
R58819 vss.n417 vss.n415 19.409
R58820 vss.n407 vss.n403 19.409
R58821 vss.n407 vss.n405 19.409
R58822 vss.n397 vss.n393 19.409
R58823 vss.n397 vss.n395 19.409
R58824 vss.n389 vss.n388 19.409
R58825 vss.n389 vss.n381 19.409
R58826 vss.n459 vss.n455 19.409
R58827 vss.n459 vss.n457 19.409
R58828 vss.n449 vss.n445 19.409
R58829 vss.n449 vss.n447 19.409
R58830 vss.n439 vss.n435 19.409
R58831 vss.n439 vss.n437 19.409
R58832 vss.n431 vss.n430 19.409
R58833 vss.n431 vss.n423 19.409
R58834 vss.n501 vss.n497 19.409
R58835 vss.n501 vss.n499 19.409
R58836 vss.n491 vss.n487 19.409
R58837 vss.n491 vss.n489 19.409
R58838 vss.n481 vss.n477 19.409
R58839 vss.n481 vss.n479 19.409
R58840 vss.n473 vss.n472 19.409
R58841 vss.n473 vss.n465 19.409
R58842 vss.n543 vss.n539 19.409
R58843 vss.n543 vss.n541 19.409
R58844 vss.n533 vss.n529 19.409
R58845 vss.n533 vss.n531 19.409
R58846 vss.n523 vss.n519 19.409
R58847 vss.n523 vss.n521 19.409
R58848 vss.n515 vss.n514 19.409
R58849 vss.n515 vss.n507 19.409
R58850 vss.n585 vss.n581 19.409
R58851 vss.n585 vss.n583 19.409
R58852 vss.n575 vss.n571 19.409
R58853 vss.n575 vss.n573 19.409
R58854 vss.n565 vss.n561 19.409
R58855 vss.n565 vss.n563 19.409
R58856 vss.n557 vss.n556 19.409
R58857 vss.n557 vss.n549 19.409
R58858 vss.n627 vss.n623 19.409
R58859 vss.n627 vss.n625 19.409
R58860 vss.n617 vss.n613 19.409
R58861 vss.n617 vss.n615 19.409
R58862 vss.n607 vss.n603 19.409
R58863 vss.n607 vss.n605 19.409
R58864 vss.n599 vss.n598 19.409
R58865 vss.n599 vss.n591 19.409
R58866 vss.n669 vss.n665 19.409
R58867 vss.n669 vss.n667 19.409
R58868 vss.n659 vss.n655 19.409
R58869 vss.n659 vss.n657 19.409
R58870 vss.n649 vss.n645 19.409
R58871 vss.n649 vss.n647 19.409
R58872 vss.n641 vss.n640 19.409
R58873 vss.n641 vss.n633 19.409
R58874 vss.n711 vss.n707 19.409
R58875 vss.n711 vss.n709 19.409
R58876 vss.n701 vss.n697 19.409
R58877 vss.n701 vss.n699 19.409
R58878 vss.n691 vss.n687 19.409
R58879 vss.n691 vss.n689 19.409
R58880 vss.n683 vss.n682 19.409
R58881 vss.n683 vss.n675 19.409
R58882 vss.n753 vss.n749 19.409
R58883 vss.n753 vss.n751 19.409
R58884 vss.n743 vss.n739 19.409
R58885 vss.n743 vss.n741 19.409
R58886 vss.n733 vss.n729 19.409
R58887 vss.n733 vss.n731 19.409
R58888 vss.n725 vss.n724 19.409
R58889 vss.n725 vss.n717 19.409
R58890 vss.n795 vss.n791 19.409
R58891 vss.n795 vss.n793 19.409
R58892 vss.n785 vss.n781 19.409
R58893 vss.n785 vss.n783 19.409
R58894 vss.n775 vss.n771 19.409
R58895 vss.n775 vss.n773 19.409
R58896 vss.n767 vss.n766 19.409
R58897 vss.n767 vss.n759 19.409
R58898 vss.n837 vss.n833 19.409
R58899 vss.n837 vss.n835 19.409
R58900 vss.n827 vss.n823 19.409
R58901 vss.n827 vss.n825 19.409
R58902 vss.n817 vss.n813 19.409
R58903 vss.n817 vss.n815 19.409
R58904 vss.n809 vss.n808 19.409
R58905 vss.n809 vss.n801 19.409
R58906 vss.n879 vss.n875 19.409
R58907 vss.n879 vss.n877 19.409
R58908 vss.n869 vss.n865 19.409
R58909 vss.n869 vss.n867 19.409
R58910 vss.n859 vss.n855 19.409
R58911 vss.n859 vss.n857 19.409
R58912 vss.n851 vss.n850 19.409
R58913 vss.n851 vss.n843 19.409
R58914 vss.n921 vss.n917 19.409
R58915 vss.n921 vss.n919 19.409
R58916 vss.n911 vss.n907 19.409
R58917 vss.n911 vss.n909 19.409
R58918 vss.n901 vss.n897 19.409
R58919 vss.n901 vss.n899 19.409
R58920 vss.n893 vss.n892 19.409
R58921 vss.n893 vss.n885 19.409
R58922 vss.n963 vss.n959 19.409
R58923 vss.n963 vss.n961 19.409
R58924 vss.n953 vss.n949 19.409
R58925 vss.n953 vss.n951 19.409
R58926 vss.n943 vss.n939 19.409
R58927 vss.n943 vss.n941 19.409
R58928 vss.n935 vss.n934 19.409
R58929 vss.n935 vss.n927 19.409
R58930 vss.n1005 vss.n1001 19.409
R58931 vss.n1005 vss.n1003 19.409
R58932 vss.n995 vss.n991 19.409
R58933 vss.n995 vss.n993 19.409
R58934 vss.n985 vss.n981 19.409
R58935 vss.n985 vss.n983 19.409
R58936 vss.n977 vss.n976 19.409
R58937 vss.n977 vss.n969 19.409
R58938 vss.n1047 vss.n1043 19.409
R58939 vss.n1047 vss.n1045 19.409
R58940 vss.n1037 vss.n1033 19.409
R58941 vss.n1037 vss.n1035 19.409
R58942 vss.n1027 vss.n1023 19.409
R58943 vss.n1027 vss.n1025 19.409
R58944 vss.n1019 vss.n1018 19.409
R58945 vss.n1019 vss.n1011 19.409
R58946 vss.n1089 vss.n1085 19.409
R58947 vss.n1089 vss.n1087 19.409
R58948 vss.n1079 vss.n1075 19.409
R58949 vss.n1079 vss.n1077 19.409
R58950 vss.n1069 vss.n1065 19.409
R58951 vss.n1069 vss.n1067 19.409
R58952 vss.n1061 vss.n1060 19.409
R58953 vss.n1061 vss.n1053 19.409
R58954 vss.n1131 vss.n1127 19.409
R58955 vss.n1131 vss.n1129 19.409
R58956 vss.n1121 vss.n1117 19.409
R58957 vss.n1121 vss.n1119 19.409
R58958 vss.n1111 vss.n1107 19.409
R58959 vss.n1111 vss.n1109 19.409
R58960 vss.n1103 vss.n1102 19.409
R58961 vss.n1103 vss.n1095 19.409
R58962 vss.n1173 vss.n1169 19.409
R58963 vss.n1173 vss.n1171 19.409
R58964 vss.n1163 vss.n1159 19.409
R58965 vss.n1163 vss.n1161 19.409
R58966 vss.n1153 vss.n1149 19.409
R58967 vss.n1153 vss.n1151 19.409
R58968 vss.n1145 vss.n1144 19.409
R58969 vss.n1145 vss.n1137 19.409
R58970 vss.n1215 vss.n1211 19.409
R58971 vss.n1215 vss.n1213 19.409
R58972 vss.n1205 vss.n1201 19.409
R58973 vss.n1205 vss.n1203 19.409
R58974 vss.n1195 vss.n1191 19.409
R58975 vss.n1195 vss.n1193 19.409
R58976 vss.n1187 vss.n1186 19.409
R58977 vss.n1187 vss.n1179 19.409
R58978 vss.n1257 vss.n1253 19.409
R58979 vss.n1257 vss.n1255 19.409
R58980 vss.n1247 vss.n1243 19.409
R58981 vss.n1247 vss.n1245 19.409
R58982 vss.n1237 vss.n1233 19.409
R58983 vss.n1237 vss.n1235 19.409
R58984 vss.n1229 vss.n1228 19.409
R58985 vss.n1229 vss.n1221 19.409
R58986 vss.n1299 vss.n1295 19.409
R58987 vss.n1299 vss.n1297 19.409
R58988 vss.n1289 vss.n1285 19.409
R58989 vss.n1289 vss.n1287 19.409
R58990 vss.n1279 vss.n1275 19.409
R58991 vss.n1279 vss.n1277 19.409
R58992 vss.n1271 vss.n1270 19.409
R58993 vss.n1271 vss.n1263 19.409
R58994 vss.n1341 vss.n1337 19.409
R58995 vss.n1341 vss.n1339 19.409
R58996 vss.n1331 vss.n1327 19.409
R58997 vss.n1331 vss.n1329 19.409
R58998 vss.n1321 vss.n1317 19.409
R58999 vss.n1321 vss.n1319 19.409
R59000 vss.n1313 vss.n1312 19.409
R59001 vss.n1313 vss.n1305 19.409
R59002 vss.n1383 vss.n1379 19.409
R59003 vss.n1383 vss.n1381 19.409
R59004 vss.n1373 vss.n1369 19.409
R59005 vss.n1373 vss.n1371 19.409
R59006 vss.n1363 vss.n1359 19.409
R59007 vss.n1363 vss.n1361 19.409
R59008 vss.n1355 vss.n1354 19.409
R59009 vss.n1355 vss.n1347 19.409
R59010 vss.n1425 vss.n1421 19.409
R59011 vss.n1425 vss.n1423 19.409
R59012 vss.n1415 vss.n1411 19.409
R59013 vss.n1415 vss.n1413 19.409
R59014 vss.n1405 vss.n1401 19.409
R59015 vss.n1405 vss.n1403 19.409
R59016 vss.n1397 vss.n1396 19.409
R59017 vss.n1397 vss.n1389 19.409
R59018 vss.n1467 vss.n1463 19.409
R59019 vss.n1467 vss.n1465 19.409
R59020 vss.n1457 vss.n1453 19.409
R59021 vss.n1457 vss.n1455 19.409
R59022 vss.n1447 vss.n1443 19.409
R59023 vss.n1447 vss.n1445 19.409
R59024 vss.n1439 vss.n1438 19.409
R59025 vss.n1439 vss.n1431 19.409
R59026 vss.n1509 vss.n1505 19.409
R59027 vss.n1509 vss.n1507 19.409
R59028 vss.n1499 vss.n1495 19.409
R59029 vss.n1499 vss.n1497 19.409
R59030 vss.n1489 vss.n1485 19.409
R59031 vss.n1489 vss.n1487 19.409
R59032 vss.n1481 vss.n1480 19.409
R59033 vss.n1481 vss.n1473 19.409
R59034 vss.n1551 vss.n1547 19.409
R59035 vss.n1551 vss.n1549 19.409
R59036 vss.n1541 vss.n1537 19.409
R59037 vss.n1541 vss.n1539 19.409
R59038 vss.n1531 vss.n1527 19.409
R59039 vss.n1531 vss.n1529 19.409
R59040 vss.n1523 vss.n1522 19.409
R59041 vss.n1523 vss.n1515 19.409
R59042 vss.n1593 vss.n1589 19.409
R59043 vss.n1593 vss.n1591 19.409
R59044 vss.n1583 vss.n1579 19.409
R59045 vss.n1583 vss.n1581 19.409
R59046 vss.n1573 vss.n1569 19.409
R59047 vss.n1573 vss.n1571 19.409
R59048 vss.n1565 vss.n1564 19.409
R59049 vss.n1565 vss.n1557 19.409
R59050 vss.n1635 vss.n1631 19.409
R59051 vss.n1635 vss.n1633 19.409
R59052 vss.n1625 vss.n1621 19.409
R59053 vss.n1625 vss.n1623 19.409
R59054 vss.n1615 vss.n1611 19.409
R59055 vss.n1615 vss.n1613 19.409
R59056 vss.n1607 vss.n1606 19.409
R59057 vss.n1607 vss.n1599 19.409
R59058 vss.n1677 vss.n1673 19.409
R59059 vss.n1677 vss.n1675 19.409
R59060 vss.n1667 vss.n1663 19.409
R59061 vss.n1667 vss.n1665 19.409
R59062 vss.n1657 vss.n1653 19.409
R59063 vss.n1657 vss.n1655 19.409
R59064 vss.n1649 vss.n1648 19.409
R59065 vss.n1649 vss.n1641 19.409
R59066 vss.n1719 vss.n1715 19.409
R59067 vss.n1719 vss.n1717 19.409
R59068 vss.n1709 vss.n1705 19.409
R59069 vss.n1709 vss.n1707 19.409
R59070 vss.n1699 vss.n1695 19.409
R59071 vss.n1699 vss.n1697 19.409
R59072 vss.n1691 vss.n1690 19.409
R59073 vss.n1691 vss.n1683 19.409
R59074 vss.n1761 vss.n1757 19.409
R59075 vss.n1761 vss.n1759 19.409
R59076 vss.n1751 vss.n1747 19.409
R59077 vss.n1751 vss.n1749 19.409
R59078 vss.n1741 vss.n1737 19.409
R59079 vss.n1741 vss.n1739 19.409
R59080 vss.n1733 vss.n1732 19.409
R59081 vss.n1733 vss.n1725 19.409
R59082 vss.n1803 vss.n1799 19.409
R59083 vss.n1803 vss.n1801 19.409
R59084 vss.n1793 vss.n1789 19.409
R59085 vss.n1793 vss.n1791 19.409
R59086 vss.n1783 vss.n1779 19.409
R59087 vss.n1783 vss.n1781 19.409
R59088 vss.n1775 vss.n1774 19.409
R59089 vss.n1775 vss.n1767 19.409
R59090 vss.n1845 vss.n1841 19.409
R59091 vss.n1845 vss.n1843 19.409
R59092 vss.n1835 vss.n1831 19.409
R59093 vss.n1835 vss.n1833 19.409
R59094 vss.n1825 vss.n1821 19.409
R59095 vss.n1825 vss.n1823 19.409
R59096 vss.n1817 vss.n1816 19.409
R59097 vss.n1817 vss.n1809 19.409
R59098 vss.n1887 vss.n1883 19.409
R59099 vss.n1887 vss.n1885 19.409
R59100 vss.n1877 vss.n1873 19.409
R59101 vss.n1877 vss.n1875 19.409
R59102 vss.n1867 vss.n1863 19.409
R59103 vss.n1867 vss.n1865 19.409
R59104 vss.n1859 vss.n1858 19.409
R59105 vss.n1859 vss.n1851 19.409
R59106 vss.n1929 vss.n1925 19.409
R59107 vss.n1929 vss.n1927 19.409
R59108 vss.n1919 vss.n1915 19.409
R59109 vss.n1919 vss.n1917 19.409
R59110 vss.n1909 vss.n1905 19.409
R59111 vss.n1909 vss.n1907 19.409
R59112 vss.n1901 vss.n1900 19.409
R59113 vss.n1901 vss.n1893 19.409
R59114 vss.n1971 vss.n1967 19.409
R59115 vss.n1971 vss.n1969 19.409
R59116 vss.n1961 vss.n1957 19.409
R59117 vss.n1961 vss.n1959 19.409
R59118 vss.n1951 vss.n1947 19.409
R59119 vss.n1951 vss.n1949 19.409
R59120 vss.n1943 vss.n1942 19.409
R59121 vss.n1943 vss.n1935 19.409
R59122 vss.n2013 vss.n2009 19.409
R59123 vss.n2013 vss.n2011 19.409
R59124 vss.n2003 vss.n1999 19.409
R59125 vss.n2003 vss.n2001 19.409
R59126 vss.n1993 vss.n1989 19.409
R59127 vss.n1993 vss.n1991 19.409
R59128 vss.n1985 vss.n1984 19.409
R59129 vss.n1985 vss.n1977 19.409
R59130 vss.n2055 vss.n2051 19.409
R59131 vss.n2055 vss.n2053 19.409
R59132 vss.n2045 vss.n2041 19.409
R59133 vss.n2045 vss.n2043 19.409
R59134 vss.n2035 vss.n2031 19.409
R59135 vss.n2035 vss.n2033 19.409
R59136 vss.n2027 vss.n2026 19.409
R59137 vss.n2027 vss.n2019 19.409
R59138 vss.n2097 vss.n2093 19.409
R59139 vss.n2097 vss.n2095 19.409
R59140 vss.n2087 vss.n2083 19.409
R59141 vss.n2087 vss.n2085 19.409
R59142 vss.n2077 vss.n2073 19.409
R59143 vss.n2077 vss.n2075 19.409
R59144 vss.n2069 vss.n2068 19.409
R59145 vss.n2069 vss.n2061 19.409
R59146 vss.n2139 vss.n2135 19.409
R59147 vss.n2139 vss.n2137 19.409
R59148 vss.n2129 vss.n2125 19.409
R59149 vss.n2129 vss.n2127 19.409
R59150 vss.n2119 vss.n2115 19.409
R59151 vss.n2119 vss.n2117 19.409
R59152 vss.n2111 vss.n2110 19.409
R59153 vss.n2111 vss.n2103 19.409
R59154 vss.n2181 vss.n2177 19.409
R59155 vss.n2181 vss.n2179 19.409
R59156 vss.n2171 vss.n2167 19.409
R59157 vss.n2171 vss.n2169 19.409
R59158 vss.n2161 vss.n2157 19.409
R59159 vss.n2161 vss.n2159 19.409
R59160 vss.n2153 vss.n2152 19.409
R59161 vss.n2153 vss.n2145 19.409
R59162 vss.n2223 vss.n2219 19.409
R59163 vss.n2223 vss.n2221 19.409
R59164 vss.n2213 vss.n2209 19.409
R59165 vss.n2213 vss.n2211 19.409
R59166 vss.n2203 vss.n2199 19.409
R59167 vss.n2203 vss.n2201 19.409
R59168 vss.n2195 vss.n2194 19.409
R59169 vss.n2195 vss.n2187 19.409
R59170 vss.n2265 vss.n2261 19.409
R59171 vss.n2265 vss.n2263 19.409
R59172 vss.n2255 vss.n2251 19.409
R59173 vss.n2255 vss.n2253 19.409
R59174 vss.n2245 vss.n2241 19.409
R59175 vss.n2245 vss.n2243 19.409
R59176 vss.n2237 vss.n2236 19.409
R59177 vss.n2237 vss.n2229 19.409
R59178 vss.n2307 vss.n2303 19.409
R59179 vss.n2307 vss.n2305 19.409
R59180 vss.n2297 vss.n2293 19.409
R59181 vss.n2297 vss.n2295 19.409
R59182 vss.n2287 vss.n2283 19.409
R59183 vss.n2287 vss.n2285 19.409
R59184 vss.n2279 vss.n2278 19.409
R59185 vss.n2279 vss.n2271 19.409
R59186 vss.n2349 vss.n2345 19.409
R59187 vss.n2349 vss.n2347 19.409
R59188 vss.n2339 vss.n2335 19.409
R59189 vss.n2339 vss.n2337 19.409
R59190 vss.n2329 vss.n2325 19.409
R59191 vss.n2329 vss.n2327 19.409
R59192 vss.n2321 vss.n2320 19.409
R59193 vss.n2321 vss.n2313 19.409
R59194 vss.n2391 vss.n2387 19.409
R59195 vss.n2391 vss.n2389 19.409
R59196 vss.n2381 vss.n2377 19.409
R59197 vss.n2381 vss.n2379 19.409
R59198 vss.n2371 vss.n2367 19.409
R59199 vss.n2371 vss.n2369 19.409
R59200 vss.n2363 vss.n2362 19.409
R59201 vss.n2363 vss.n2355 19.409
R59202 vss.n3183 vss.t580 4.356
R59203 vss.n2396 vss.t45 4.356
R59204 vss.n3188 vss.t328 4.355
R59205 vss.n3191 vss.t524 4.355
R59206 vss.n3196 vss.t115 4.355
R59207 vss.n3139 vss.t346 4.355
R59208 vss.n3139 vss.t144 4.355
R59209 vss.n3159 vss.t188 4.355
R59210 vss.n3159 vss.t591 4.355
R59211 vss.n3169 vss.t564 4.355
R59212 vss.n3169 vss.t357 4.355
R59213 vss.n3179 vss.t153 4.355
R59214 vss.n3179 vss.t556 4.355
R59215 vss.n3097 vss.t366 4.355
R59216 vss.n3097 vss.t340 4.355
R59217 vss.n3117 vss.t194 4.355
R59218 vss.n3117 vss.t187 4.355
R59219 vss.n3127 vss.t576 4.355
R59220 vss.n3127 vss.t558 4.355
R59221 vss.n3137 vss.t169 4.355
R59222 vss.n3137 vss.t148 4.355
R59223 vss.n3055 vss.t241 4.355
R59224 vss.n3055 vss.t361 4.355
R59225 vss.n3075 vss.t98 4.355
R59226 vss.n3075 vss.t193 4.355
R59227 vss.n3085 vss.t452 4.355
R59228 vss.n3085 vss.t571 4.355
R59229 vss.n3095 vss.t44 4.355
R59230 vss.n3095 vss.t163 4.355
R59231 vss.n3013 vss.t254 4.355
R59232 vss.n3013 vss.t582 4.355
R59233 vss.n3033 vss.t122 4.355
R59234 vss.n3033 vss.t399 4.355
R59235 vss.n3043 vss.t469 4.355
R59236 vss.n3043 vss.t185 4.355
R59237 vss.n3053 vss.t61 4.355
R59238 vss.n3053 vss.t382 4.355
R59239 vss.n2971 vss.t586 4.355
R59240 vss.n2971 vss.t459 4.355
R59241 vss.n2991 vss.t400 4.355
R59242 vss.n2991 vss.t320 4.355
R59243 vss.n3001 vss.t189 4.355
R59244 vss.n3001 vss.t70 4.355
R59245 vss.n3011 vss.t388 4.355
R59246 vss.n3011 vss.t262 4.355
R59247 vss.n2929 vss.t77 4.355
R59248 vss.n2929 vss.t480 4.355
R59249 vss.n2949 vss.t551 4.355
R59250 vss.n2949 vss.t347 4.355
R59251 vss.n2959 vss.t291 4.355
R59252 vss.n2959 vss.t87 4.355
R59253 vss.n2969 vss.t486 4.355
R59254 vss.n2969 vss.t283 4.355
R59255 vss.n2887 vss.t96 4.355
R59256 vss.n2887 vss.t495 4.355
R59257 vss.n2907 vss.t567 4.355
R59258 vss.n2907 vss.t367 4.355
R59259 vss.n2917 vss.t310 4.355
R59260 vss.n2917 vss.t105 4.355
R59261 vss.n2927 vss.t505 4.355
R59262 vss.n2927 vss.t299 4.355
R59263 vss.n2845 vss.t117 4.355
R59264 vss.n2845 vss.t407 4.355
R59265 vss.n2865 vss.t581 4.355
R59266 vss.n2865 vss.t242 4.355
R59267 vss.n2875 vss.t332 4.355
R59268 vss.n2875 vss.t9 4.355
R59269 vss.n2885 vss.t528 4.355
R59270 vss.n2885 vss.t206 4.355
R59271 vss.n2803 vss.t284 4.355
R59272 vss.n2803 vss.t316 4.355
R59273 vss.n2823 vss.t154 4.355
R59274 vss.n2823 vss.t178 4.355
R59275 vss.n2833 vss.t496 4.355
R59276 vss.n2833 vss.t538 4.355
R59277 vss.n2843 vss.t88 4.355
R59278 vss.n2843 vss.t126 4.355
R59279 vss.n2761 vss.t300 4.355
R59280 vss.n2761 vss.t596 4.355
R59281 vss.n2781 vss.t170 4.355
R59282 vss.n2781 vss.t401 4.355
R59283 vss.n2791 vss.t514 4.355
R59284 vss.n2791 vss.t196 4.355
R59285 vss.n2801 vss.t106 4.355
R59286 vss.n2801 vss.t396 4.355
R59287 vss.n2719 vss.t535 4.355
R59288 vss.n2719 vss.t506 4.355
R59289 vss.n2739 vss.t385 4.355
R59290 vss.n2739 vss.t371 4.355
R59291 vss.n2749 vss.t147 4.355
R59292 vss.n2749 vss.t118 4.355
R59293 vss.n2759 vss.t341 4.355
R59294 vss.n2759 vss.t311 4.355
R59295 vss.n2677 vss.t127 4.355
R59296 vss.n2677 vss.t529 4.355
R59297 vss.n2697 vss.t584 4.355
R59298 vss.n2697 vss.t383 4.355
R59299 vss.n2707 vss.t343 4.355
R59300 vss.n2707 vss.t140 4.355
R59301 vss.n2717 vss.t539 4.355
R59302 vss.n2717 vss.t334 4.355
R59303 vss.n2635 vss.t151 4.355
R59304 vss.n2635 vss.t552 4.355
R59305 vss.n2655 vss.t593 4.355
R59306 vss.n2655 vss.t391 4.355
R59307 vss.n2665 vss.t363 4.355
R59308 vss.n2665 vss.t158 4.355
R59309 vss.n2675 vss.t561 4.355
R59310 vss.n2675 vss.t353 4.355
R59311 vss.n2593 vss.t167 4.355
R59312 vss.n2593 vss.t35 4.355
R59313 vss.n2613 vss.t597 4.355
R59314 vss.n2613 vss.t489 4.355
R59315 vss.n2623 vss.t376 4.355
R59316 vss.n2623 vss.t244 4.355
R59317 vss.n2633 vss.t573 4.355
R59318 vss.n2633 vss.t440 4.355
R59319 vss.n2551 vss.t179 4.355
R59320 vss.n2551 vss.t48 4.355
R59321 vss.n2571 vss.t598 4.355
R59322 vss.n2571 vss.t509 4.355
R59323 vss.n2581 vss.t386 4.355
R59324 vss.n2581 vss.t257 4.355
R59325 vss.n2591 vss.t585 4.355
R59326 vss.n2591 vss.t454 4.355
R59327 vss.n2509 vss.t264 4.355
R59328 vss.n2509 vss.t64 4.355
R59329 vss.n2529 vss.t131 4.355
R59330 vss.n2529 vss.t536 4.355
R59331 vss.n2539 vss.t483 4.355
R59332 vss.n2539 vss.t275 4.355
R59333 vss.n2549 vss.t73 4.355
R59334 vss.n2549 vss.t473 4.355
R59335 vss.n2467 vss.t286 4.355
R59336 vss.n2467 vss.t389 4.355
R59337 vss.n2487 vss.t155 4.355
R59338 vss.n2487 vss.t198 4.355
R59339 vss.n2497 vss.t498 4.355
R59340 vss.n2497 vss.t594 4.355
R59341 vss.n2507 vss.t90 4.355
R59342 vss.n2507 vss.t190 4.355
R59343 vss.n0 vss.t304 4.355
R59344 vss.n0 vss.t278 4.355
R59345 vss.n20 vss.t173 4.355
R59346 vss.n20 vss.t150 4.355
R59347 vss.n30 vss.t517 4.355
R59348 vss.n30 vss.t492 4.355
R59349 vss.n40 vss.t109 4.355
R59350 vss.n40 vss.t83 4.355
R59351 vss.n42 vss.t208 4.355
R59352 vss.n42 vss.t507 4.355
R59353 vss.n62 vss.t47 4.355
R59354 vss.n62 vss.t373 4.355
R59355 vss.n72 vss.t416 4.355
R59356 vss.n72 vss.t120 4.355
R59357 vss.n82 vss.t11 4.355
R59358 vss.n82 vss.t312 4.355
R59359 vss.n84 vss.t521 4.355
R59360 vss.n84 vss.t531 4.355
R59361 vss.n104 vss.t379 4.355
R59362 vss.n104 vss.t384 4.355
R59363 vss.n114 vss.t134 4.355
R59364 vss.n114 vss.t142 4.355
R59365 vss.n124 vss.t326 4.355
R59366 vss.n124 vss.t335 4.355
R59367 vss.n126 vss.t398 4.355
R59368 vss.n126 vss.t91 4.355
R59369 vss.n146 vss.t199 4.355
R59370 vss.n146 vss.t565 4.355
R59371 vss.n156 vss.t599 4.355
R59372 vss.n156 vss.t303 4.355
R59373 vss.n166 vss.t197 4.355
R59374 vss.n166 vss.t499 4.355
R59375 vss.n168 vss.t314 4.355
R59376 vss.n168 vss.t110 4.355
R59377 vss.n188 vss.t177 4.355
R59378 vss.n188 vss.t578 4.355
R59379 vss.n198 vss.t532 4.355
R59380 vss.n198 vss.t324 4.355
R59381 vss.n208 vss.t121 4.355
R59382 vss.n208 vss.t518 4.355
R59383 vss.n210 vss.t337 4.355
R59384 vss.n210 vss.t132 4.355
R59385 vss.n230 vss.t186 4.355
R59386 vss.n230 vss.t587 4.355
R59387 vss.n240 vss.t555 4.355
R59388 vss.n240 vss.t349 4.355
R59389 vss.n250 vss.t143 4.355
R59390 vss.n250 vss.t544 4.355
R59391 vss.n252 vss.t356 4.355
R59392 vss.n252 vss.t541 4.355
R59393 vss.n272 vss.t191 4.355
R59394 vss.n272 vss.t387 4.355
R59395 vss.n282 vss.t569 4.355
R59396 vss.n282 vss.t152 4.355
R59397 vss.n292 vss.t160 4.355
R59398 vss.n292 vss.t345 4.355
R59399 vss.n294 vss.t234 4.355
R59400 vss.n294 vss.t562 4.355
R59401 vss.n314 vss.t92 4.355
R59402 vss.n314 vss.t394 4.355
R59403 vss.n324 vss.t444 4.355
R59404 vss.n324 vss.t168 4.355
R59405 vss.n334 vss.t37 4.355
R59406 vss.n334 vss.t364 4.355
R59407 vss.n336 vss.t456 4.355
R59408 vss.n336 vss.t574 4.355
R59409 vss.n356 vss.t317 4.355
R59410 vss.n356 vss.t397 4.355
R59411 vss.n366 vss.t67 4.355
R59412 vss.n366 vss.t181 4.355
R59413 vss.n376 vss.t259 4.355
R59414 vss.n376 vss.t377 4.355
R59415 vss.n378 vss.t476 4.355
R59416 vss.n378 vss.t451 4.355
R59417 vss.n398 vss.t342 4.355
R59418 vss.n398 vss.t313 4.355
R59419 vss.n408 vss.t84 4.355
R59420 vss.n408 vss.t60 4.355
R59421 vss.n418 vss.t279 4.355
R59422 vss.n418 vss.t253 4.355
R59423 vss.n420 vss.t69 4.355
R59424 vss.n420 vss.t468 4.355
R59425 vss.n440 vss.t542 4.355
R59426 vss.n440 vss.t336 4.355
R59427 vss.n450 vss.t282 4.355
R59428 vss.n450 vss.t78 4.355
R59429 vss.n460 vss.t479 4.355
R59430 vss.n460 vss.t271 4.355
R59431 vss.n462 vss.t86 4.355
R59432 vss.n462 vss.t95 4.355
R59433 vss.n482 vss.t563 4.355
R59434 vss.n482 vss.t566 4.355
R59435 vss.n492 vss.t298 4.355
R59436 vss.n492 vss.t307 4.355
R59437 vss.n502 vss.t493 4.355
R59438 vss.n502 vss.t502 4.355
R59439 vss.n504 vss.t104 4.355
R59440 vss.n504 vss.t5 4.355
R59441 vss.n524 vss.t575 4.355
R59442 vss.n524 vss.t441 4.355
R59443 vss.n534 vss.t319 4.355
R59444 vss.n534 vss.t210 4.355
R59445 vss.n544 vss.t513 4.355
R59446 vss.n544 vss.t409 4.355
R59447 vss.n546 vss.t213 4.355
R59448 vss.n546 vss.t13 4.355
R59449 vss.n566 vss.t53 4.355
R59450 vss.n566 vss.t457 4.355
R59451 vss.n576 vss.t425 4.355
R59452 vss.n576 vss.t219 4.355
R59453 vss.n586 vss.t18 4.355
R59454 vss.n586 vss.t419 4.355
R59455 vss.n588 vss.t503 4.355
R59456 vss.n588 vss.t331 4.355
R59457 vss.n608 vss.t370 4.355
R59458 vss.n608 vss.t184 4.355
R59459 vss.n618 vss.t114 4.355
R59460 vss.n618 vss.t548 4.355
R59461 vss.n628 vss.t306 4.355
R59462 vss.n628 vss.t139 4.355
R59463 vss.n630 vss.t523 4.355
R59464 vss.n630 vss.t494 4.355
R59465 vss.n650 vss.t380 4.355
R59466 vss.n650 vss.t365 4.355
R59467 vss.n660 vss.t135 4.355
R59468 vss.n660 vss.t103 4.355
R59469 vss.n670 vss.t327 4.355
R59470 vss.n670 vss.t297 4.355
R59471 vss.n672 vss.t418 4.355
R59472 vss.n672 vss.t124 4.355
R59473 vss.n692 vss.t260 4.355
R59474 vss.n692 vss.t583 4.355
R59475 vss.n702 vss.t24 4.355
R59476 vss.n702 vss.t339 4.355
R59477 vss.n712 vss.t220 4.355
R59478 vss.n712 vss.t534 4.355
R59479 vss.n714 vss.t138 4.355
R59480 vss.n714 vss.t146 4.355
R59481 vss.n734 vss.t589 4.355
R59482 vss.n734 vss.t592 4.355
R59483 vss.n744 vss.t352 4.355
R59484 vss.n744 vss.t360 4.355
R59485 vss.n754 vss.t550 4.355
R59486 vss.n754 vss.t557 4.355
R59487 vss.n756 vss.t369 4.355
R59488 vss.n756 vss.t31 4.355
R59489 vss.n776 vss.t195 4.355
R59490 vss.n776 vss.t484 4.355
R59491 vss.n786 vss.t577 4.355
R59492 vss.n786 vss.t237 4.355
R59493 vss.n796 vss.t172 4.355
R59494 vss.n796 vss.t436 4.355
R59495 vss.n798 vss.t243 4.355
R59496 vss.n798 vss.t40 4.355
R59497 vss.n818 vss.t101 4.355
R59498 vss.n818 vss.t501 4.355
R59499 vss.n828 vss.t453 4.355
R59500 vss.n828 vss.t248 4.355
R59501 vss.n838 vss.t46 4.355
R59502 vss.n838 vss.t446 4.355
R59503 vss.n840 vss.t256 4.355
R59504 vss.n840 vss.t54 4.355
R59505 vss.n860 vss.t123 4.355
R59506 vss.n860 vss.t522 4.355
R59507 vss.n870 vss.t472 4.355
R59508 vss.n870 vss.t266 4.355
R59509 vss.n880 vss.t63 4.355
R59510 vss.n880 vss.t463 4.355
R59511 vss.n882 vss.t274 4.355
R59512 vss.n882 vss.t461 4.355
R59513 vss.n902 vss.t145 4.355
R59514 vss.n902 vss.t322 4.355
R59515 vss.n912 vss.t488 4.355
R59516 vss.n912 vss.t72 4.355
R59517 vss.n922 vss.t80 4.355
R59518 vss.n922 vss.t263 4.355
R59519 vss.n924 vss.t293 4.355
R59520 vss.n924 vss.t482 4.355
R59521 vss.n944 vss.t162 4.355
R59522 vss.n944 vss.t348 4.355
R59523 vss.n954 vss.t508 4.355
R59524 vss.n954 vss.t89 4.355
R59525 vss.n964 vss.t100 4.355
R59526 vss.n964 vss.t285 4.355
R59527 vss.n966 vss.t411 4.355
R59528 vss.n966 vss.t497 4.355
R59529 vss.n986 vss.t246 4.355
R59530 vss.n986 vss.t368 4.355
R59531 vss.n996 vss.t15 4.355
R59532 vss.n996 vss.t107 4.355
R59533 vss.n1006 vss.t212 4.355
R59534 vss.n1006 vss.t302 4.355
R59535 vss.n1008 vss.t421 4.355
R59536 vss.n1008 vss.t516 4.355
R59537 vss.n1028 vss.t261 4.355
R59538 vss.n1028 vss.t378 4.355
R59539 vss.n1038 vss.t27 4.355
R59540 vss.n1038 vss.t129 4.355
R59541 vss.n1048 vss.t222 4.355
R59542 vss.n1048 vss.t321 4.355
R59543 vss.n1050 vss.t141 4.355
R59544 vss.n1050 vss.t415 4.355
R59545 vss.n1070 vss.t590 4.355
R59546 vss.n1070 vss.t255 4.355
R59547 vss.n1080 vss.t355 4.355
R59548 vss.n1080 vss.t21 4.355
R59549 vss.n1090 vss.t553 4.355
R59550 vss.n1090 vss.t217 4.355
R59551 vss.n1092 vss.t301 4.355
R59552 vss.n1092 vss.t309 4.355
R59553 vss.n1112 vss.t171 4.355
R59554 vss.n1112 vss.t175 4.355
R59555 vss.n1122 vss.t515 4.355
R59556 vss.n1122 vss.t527 4.355
R59557 vss.n1132 vss.t108 4.355
R59558 vss.n1132 vss.t116 4.355
R59559 vss.n1134 vss.t323 4.355
R59560 vss.n1134 vss.t333 4.355
R59561 vss.n1154 vss.t182 4.355
R59562 vss.n1154 vss.t183 4.355
R59563 vss.n1164 vss.t543 4.355
R59564 vss.n1164 vss.t549 4.355
R59565 vss.n1174 vss.t130 4.355
R59566 vss.n1174 vss.t137 4.355
R59567 vss.n1176 vss.t560 4.355
R59568 vss.n1176 vss.t223 4.355
R59569 vss.n1196 vss.t393 4.355
R59570 vss.n1196 vss.t68 4.355
R59571 vss.n1206 vss.t166 4.355
R59572 vss.n1206 vss.t432 4.355
R59573 vss.n1216 vss.t362 4.355
R59574 vss.n1216 vss.t26 4.355
R59575 vss.n1218 vss.t439 4.355
R59576 vss.n1218 vss.t554 4.355
R59577 vss.n1238 vss.t290 4.355
R59578 vss.n1238 vss.t392 4.355
R59579 vss.n1248 vss.t42 4.355
R59580 vss.n1248 vss.t159 4.355
R59581 vss.n1258 vss.t238 4.355
R59582 vss.n1258 vss.t354 4.355
R59583 vss.n1260 vss.t449 4.355
R59584 vss.n1260 vss.t568 4.355
R59585 vss.n1280 vss.t308 4.355
R59586 vss.n1280 vss.t395 4.355
R59587 vss.n1290 vss.t56 4.355
R59588 vss.n1290 vss.t176 4.355
R59589 vss.n1300 vss.t250 4.355
R59590 vss.n1300 vss.t372 4.355
R59591 vss.n1302 vss.t465 4.355
R59592 vss.n1302 vss.t50 4.355
R59593 vss.n1322 vss.t330 4.355
R59594 vss.n1322 vss.t511 4.355
R59595 vss.n1332 vss.t76 4.355
R59596 vss.n1332 vss.t258 4.355
R59597 vss.n1342 vss.t268 4.355
R59598 vss.n1342 vss.t455 4.355
R59599 vss.n1344 vss.t59 4.355
R59600 vss.n1344 vss.t66 4.355
R59601 vss.n1364 vss.t530 4.355
R59602 vss.n1364 vss.t537 4.355
R59603 vss.n1374 vss.t270 4.355
R59604 vss.n1374 vss.t277 4.355
R59605 vss.n1384 vss.t467 4.355
R59606 vss.n1384 vss.t475 4.355
R59607 vss.n1386 vss.t288 4.355
R59608 vss.n1386 vss.t82 4.355
R59609 vss.n1406 vss.t156 4.355
R59610 vss.n1406 vss.t559 4.355
R59611 vss.n1416 vss.t500 4.355
R59612 vss.n1416 vss.t295 4.355
R59613 vss.n1426 vss.t94 4.355
R59614 vss.n1426 vss.t491 4.355
R59615 vss.n1428 vss.t305 4.355
R59616 vss.n1428 vss.t2 4.355
R59617 vss.n1448 vss.t174 4.355
R59618 vss.n1448 vss.t438 4.355
R59619 vss.n1458 vss.t520 4.355
R59620 vss.n1458 vss.t204 4.355
R59621 vss.n1468 vss.t112 4.355
R59622 vss.n1468 vss.t405 4.355
R59623 vss.n1470 vss.t209 4.355
R59624 vss.n1470 vss.t7 4.355
R59625 vss.n1490 vss.t49 4.355
R59626 vss.n1490 vss.t448 4.355
R59627 vss.n1500 vss.t417 4.355
R59628 vss.n1500 vss.t214 4.355
R59629 vss.n1510 vss.t12 4.355
R59630 vss.n1510 vss.t412 4.355
R59631 vss.n1512 vss.t218 4.355
R59632 vss.n1512 vss.t225 4.355
R59633 vss.n1532 vss.t65 4.355
R59634 vss.n1532 vss.t71 4.355
R59635 vss.n1542 vss.t428 4.355
R59636 vss.n1542 vss.t433 4.355
R59637 vss.n1552 vss.t23 4.355
R59638 vss.n1552 vss.t29 4.355
R59639 vss.n1554 vss.t512 4.355
R59640 vss.n1554 vss.t424 4.355
R59641 vss.n1574 vss.t375 4.355
R59642 vss.n1574 vss.t265 4.355
R59643 vss.n1584 vss.t125 4.355
R59644 vss.n1584 vss.t30 4.355
R59645 vss.n1594 vss.t315 4.355
R59646 vss.n1594 vss.t226 4.355
R59647 vss.n1596 vss.t17 4.355
R59648 vss.n1596 vss.t113 4.355
R59649 vss.n1616 vss.t460 4.355
R59650 vss.n1616 vss.t579 4.355
R59651 vss.n1626 vss.t224 4.355
R59652 vss.n1626 vss.t325 4.355
R59653 vss.n1636 vss.t422 4.355
R59654 vss.n1636 vss.t519 4.355
R59655 vss.n1638 vss.t28 4.355
R59656 vss.n1638 vss.t133 4.355
R59657 vss.n1658 vss.t481 4.355
R59658 vss.n1658 vss.t588 4.355
R59659 vss.n1668 vss.t233 4.355
R59660 vss.n1668 vss.t350 4.355
R59661 vss.n1678 vss.t434 4.355
R59662 vss.n1678 vss.t545 4.355
R59663 vss.n1680 vss.t359 4.355
R59664 vss.n1680 vss.t22 4.355
R59665 vss.n1700 vss.t192 4.355
R59666 vss.n1700 vss.t474 4.355
R59667 vss.n1710 vss.t570 4.355
R59668 vss.n1710 vss.t230 4.355
R59669 vss.n1720 vss.t161 4.355
R59670 vss.n1720 vss.t429 4.355
R59671 vss.n1722 vss.t236 4.355
R59672 vss.n1722 vss.t240 4.355
R59673 vss.n1742 vss.t93 4.355
R59674 vss.n1742 vss.t97 4.355
R59675 vss.n1752 vss.t445 4.355
R59676 vss.n1752 vss.t450 4.355
R59677 vss.n1762 vss.t39 4.355
R59678 vss.n1762 vss.t43 4.355
R59679 vss.n1764 vss.t247 4.355
R59680 vss.n1764 vss.t252 4.355
R59681 vss.n1784 vss.t111 4.355
R59682 vss.n1784 vss.t119 4.355
R59683 vss.n1794 vss.t462 4.355
R59684 vss.n1794 vss.t466 4.355
R59685 vss.n1804 vss.t52 4.355
R59686 vss.n1804 vss.t58 4.355
R59687 vss.n1806 vss.t478 4.355
R59688 vss.n1806 vss.t200 4.355
R59689 vss.n1826 vss.t344 4.355
R59690 vss.n1826 vss.t16 4.355
R59691 vss.n1836 vss.t85 4.355
R59692 vss.n1836 vss.t402 4.355
R59693 vss.n1846 vss.t281 4.355
R59694 vss.n1846 vss.t0 4.355
R59695 vss.n1848 vss.t404 4.355
R59696 vss.n1848 vss.t471 4.355
R59697 vss.n1868 vss.t229 4.355
R59698 vss.n1868 vss.t338 4.355
R59699 vss.n1878 vss.t3 4.355
R59700 vss.n1878 vss.t79 4.355
R59701 vss.n1888 vss.t202 4.355
R59702 vss.n1888 vss.t273 4.355
R59703 vss.n1890 vss.t406 4.355
R59704 vss.n1890 vss.t487 4.355
R59705 vss.n1910 vss.t239 4.355
R59706 vss.n1910 vss.t358 4.355
R59707 vss.n1920 vss.t8 4.355
R59708 vss.n1920 vss.t99 4.355
R59709 vss.n1930 vss.t205 4.355
R59710 vss.n1930 vss.t292 4.355
R59711 vss.n1932 vss.t413 4.355
R59712 vss.n1932 vss.t6 4.355
R59713 vss.n1952 vss.t251 4.355
R59714 vss.n1952 vss.t442 4.355
R59715 vss.n1962 vss.t19 4.355
R59716 vss.n1962 vss.t211 4.355
R59717 vss.n1972 vss.t215 4.355
R59718 vss.n1972 vss.t410 4.355
R59719 vss.n1974 vss.t426 4.355
R59720 vss.n1974 vss.t14 4.355
R59721 vss.n1994 vss.t269 4.355
R59722 vss.n1994 vss.t458 4.355
R59723 vss.n2004 vss.t33 4.355
R59724 vss.n2004 vss.t221 4.355
R59725 vss.n2014 vss.t228 4.355
R59726 vss.n2014 vss.t420 4.355
R59727 vss.n2016 vss.t227 4.355
R59728 vss.n2016 vss.t25 4.355
R59729 vss.n2036 vss.t74 4.355
R59730 vss.n2036 vss.t477 4.355
R59731 vss.n2046 vss.t437 4.355
R59732 vss.n2046 vss.t231 4.355
R59733 vss.n2056 vss.t32 4.355
R59734 vss.n2056 vss.t430 4.355
R59735 vss.n2058 vss.t525 4.355
R59736 vss.n2058 vss.t318 4.355
R59737 vss.n2078 vss.t381 4.355
R59738 vss.n2078 vss.t180 4.355
R59739 vss.n2088 vss.t136 4.355
R59740 vss.n2088 vss.t540 4.355
R59741 vss.n2098 vss.t329 4.355
R59742 vss.n2098 vss.t128 4.355
R59743 vss.n2100 vss.t547 4.355
R59744 vss.n2100 vss.t216 4.355
R59745 vss.n2120 vss.t390 4.355
R59746 vss.n2120 vss.t57 4.355
R59747 vss.n2130 vss.t157 4.355
R59748 vss.n2130 vss.t427 4.355
R59749 vss.n2140 vss.t351 4.355
R59750 vss.n2140 vss.t20 4.355
R59751 vss.n2142 vss.t431 4.355
R59752 vss.n2142 vss.t435 4.355
R59753 vss.n2162 vss.t280 4.355
R59754 vss.n2162 vss.t287 4.355
R59755 vss.n2172 vss.t36 4.355
R59756 vss.n2172 vss.t38 4.355
R59757 vss.n2182 vss.t232 4.355
R59758 vss.n2182 vss.t235 4.355
R59759 vss.n2184 vss.t443 4.355
R59760 vss.n2184 vss.t165 4.355
R59761 vss.n2204 vss.t296 4.355
R59762 vss.n2204 vss.t595 4.355
R59763 vss.n2214 vss.t51 4.355
R59764 vss.n2214 vss.t374 4.355
R59765 vss.n2224 vss.t245 4.355
R59766 vss.n2224 vss.t572 4.355
R59767 vss.n2226 vss.t62 4.355
R59768 vss.n2226 vss.t41 4.355
R59769 vss.n2246 vss.t533 4.355
R59770 vss.n2246 vss.t504 4.355
R59771 vss.n2256 vss.t272 4.355
R59772 vss.n2256 vss.t249 4.355
R59773 vss.n2266 vss.t470 4.355
R59774 vss.n2266 vss.t447 4.355
R59775 vss.n2268 vss.t1 4.355
R59776 vss.n2268 vss.t55 4.355
R59777 vss.n2288 vss.t423 4.355
R59778 vss.n2288 vss.t526 4.355
R59779 vss.n2298 vss.t201 4.355
R59780 vss.n2298 vss.t267 4.355
R59781 vss.n2308 vss.t403 4.355
R59782 vss.n2308 vss.t464 4.355
R59783 vss.n2310 vss.t276 4.355
R59784 vss.n2310 vss.t75 4.355
R59785 vss.n2330 vss.t149 4.355
R59786 vss.n2330 vss.t546 4.355
R59787 vss.n2340 vss.t490 4.355
R59788 vss.n2340 vss.t289 4.355
R59789 vss.n2350 vss.t81 4.355
R59790 vss.n2350 vss.t485 4.355
R59791 vss.n2352 vss.t294 4.355
R59792 vss.n2352 vss.t203 4.355
R59793 vss.n2372 vss.t164 4.355
R59794 vss.n2372 vss.t34 4.355
R59795 vss.n2382 vss.t510 4.355
R59796 vss.n2382 vss.t408 4.355
R59797 vss.n2392 vss.t102 4.355
R59798 vss.n2392 vss.t4 4.355
R59799 vss.n2401 vss.t414 4.355
R59800 vss.n2404 vss.t10 4.355
R59801 vss.n2409 vss.t207 4.355
R59802 vss.n3173 vss.n3172 2.703
R59803 vss.n3171 vss.n3170 2.703
R59804 vss.n3131 vss.n3130 2.703
R59805 vss.n3129 vss.n3128 2.703
R59806 vss.n3089 vss.n3088 2.703
R59807 vss.n3087 vss.n3086 2.703
R59808 vss.n3047 vss.n3046 2.703
R59809 vss.n3045 vss.n3044 2.703
R59810 vss.n3005 vss.n3004 2.703
R59811 vss.n3003 vss.n3002 2.703
R59812 vss.n2963 vss.n2962 2.703
R59813 vss.n2961 vss.n2960 2.703
R59814 vss.n2921 vss.n2920 2.703
R59815 vss.n2919 vss.n2918 2.703
R59816 vss.n2879 vss.n2878 2.703
R59817 vss.n2877 vss.n2876 2.703
R59818 vss.n2837 vss.n2836 2.703
R59819 vss.n2835 vss.n2834 2.703
R59820 vss.n2795 vss.n2794 2.703
R59821 vss.n2793 vss.n2792 2.703
R59822 vss.n2753 vss.n2752 2.703
R59823 vss.n2751 vss.n2750 2.703
R59824 vss.n2711 vss.n2710 2.703
R59825 vss.n2709 vss.n2708 2.703
R59826 vss.n2669 vss.n2668 2.703
R59827 vss.n2667 vss.n2666 2.703
R59828 vss.n2627 vss.n2626 2.703
R59829 vss.n2625 vss.n2624 2.703
R59830 vss.n2585 vss.n2584 2.703
R59831 vss.n2583 vss.n2582 2.703
R59832 vss.n2543 vss.n2542 2.703
R59833 vss.n2541 vss.n2540 2.703
R59834 vss.n2501 vss.n2500 2.703
R59835 vss.n2499 vss.n2498 2.703
R59836 vss.n34 vss.n33 2.703
R59837 vss.n32 vss.n31 2.703
R59838 vss.n76 vss.n75 2.703
R59839 vss.n74 vss.n73 2.703
R59840 vss.n118 vss.n117 2.703
R59841 vss.n116 vss.n115 2.703
R59842 vss.n160 vss.n159 2.703
R59843 vss.n158 vss.n157 2.703
R59844 vss.n202 vss.n201 2.703
R59845 vss.n200 vss.n199 2.703
R59846 vss.n244 vss.n243 2.703
R59847 vss.n242 vss.n241 2.703
R59848 vss.n286 vss.n285 2.703
R59849 vss.n284 vss.n283 2.703
R59850 vss.n328 vss.n327 2.703
R59851 vss.n326 vss.n325 2.703
R59852 vss.n370 vss.n369 2.703
R59853 vss.n368 vss.n367 2.703
R59854 vss.n412 vss.n411 2.703
R59855 vss.n410 vss.n409 2.703
R59856 vss.n454 vss.n453 2.703
R59857 vss.n452 vss.n451 2.703
R59858 vss.n496 vss.n495 2.703
R59859 vss.n494 vss.n493 2.703
R59860 vss.n538 vss.n537 2.703
R59861 vss.n536 vss.n535 2.703
R59862 vss.n580 vss.n579 2.703
R59863 vss.n578 vss.n577 2.703
R59864 vss.n622 vss.n621 2.703
R59865 vss.n620 vss.n619 2.703
R59866 vss.n664 vss.n663 2.703
R59867 vss.n662 vss.n661 2.703
R59868 vss.n706 vss.n705 2.703
R59869 vss.n704 vss.n703 2.703
R59870 vss.n748 vss.n747 2.703
R59871 vss.n746 vss.n745 2.703
R59872 vss.n790 vss.n789 2.703
R59873 vss.n788 vss.n787 2.703
R59874 vss.n832 vss.n831 2.703
R59875 vss.n830 vss.n829 2.703
R59876 vss.n874 vss.n873 2.703
R59877 vss.n872 vss.n871 2.703
R59878 vss.n916 vss.n915 2.703
R59879 vss.n914 vss.n913 2.703
R59880 vss.n958 vss.n957 2.703
R59881 vss.n956 vss.n955 2.703
R59882 vss.n1000 vss.n999 2.703
R59883 vss.n998 vss.n997 2.703
R59884 vss.n1042 vss.n1041 2.703
R59885 vss.n1040 vss.n1039 2.703
R59886 vss.n1084 vss.n1083 2.703
R59887 vss.n1082 vss.n1081 2.703
R59888 vss.n1126 vss.n1125 2.703
R59889 vss.n1124 vss.n1123 2.703
R59890 vss.n1168 vss.n1167 2.703
R59891 vss.n1166 vss.n1165 2.703
R59892 vss.n1210 vss.n1209 2.703
R59893 vss.n1208 vss.n1207 2.703
R59894 vss.n1252 vss.n1251 2.703
R59895 vss.n1250 vss.n1249 2.703
R59896 vss.n1294 vss.n1293 2.703
R59897 vss.n1292 vss.n1291 2.703
R59898 vss.n1336 vss.n1335 2.703
R59899 vss.n1334 vss.n1333 2.703
R59900 vss.n1378 vss.n1377 2.703
R59901 vss.n1376 vss.n1375 2.703
R59902 vss.n1420 vss.n1419 2.703
R59903 vss.n1418 vss.n1417 2.703
R59904 vss.n1462 vss.n1461 2.703
R59905 vss.n1460 vss.n1459 2.703
R59906 vss.n1504 vss.n1503 2.703
R59907 vss.n1502 vss.n1501 2.703
R59908 vss.n1546 vss.n1545 2.703
R59909 vss.n1544 vss.n1543 2.703
R59910 vss.n1588 vss.n1587 2.703
R59911 vss.n1586 vss.n1585 2.703
R59912 vss.n1630 vss.n1629 2.703
R59913 vss.n1628 vss.n1627 2.703
R59914 vss.n1672 vss.n1671 2.703
R59915 vss.n1670 vss.n1669 2.703
R59916 vss.n1714 vss.n1713 2.703
R59917 vss.n1712 vss.n1711 2.703
R59918 vss.n1756 vss.n1755 2.703
R59919 vss.n1754 vss.n1753 2.703
R59920 vss.n1798 vss.n1797 2.703
R59921 vss.n1796 vss.n1795 2.703
R59922 vss.n1840 vss.n1839 2.703
R59923 vss.n1838 vss.n1837 2.703
R59924 vss.n1882 vss.n1881 2.703
R59925 vss.n1880 vss.n1879 2.703
R59926 vss.n1924 vss.n1923 2.703
R59927 vss.n1922 vss.n1921 2.703
R59928 vss.n1966 vss.n1965 2.703
R59929 vss.n1964 vss.n1963 2.703
R59930 vss.n2008 vss.n2007 2.703
R59931 vss.n2006 vss.n2005 2.703
R59932 vss.n2050 vss.n2049 2.703
R59933 vss.n2048 vss.n2047 2.703
R59934 vss.n2092 vss.n2091 2.703
R59935 vss.n2090 vss.n2089 2.703
R59936 vss.n2134 vss.n2133 2.703
R59937 vss.n2132 vss.n2131 2.703
R59938 vss.n2176 vss.n2175 2.703
R59939 vss.n2174 vss.n2173 2.703
R59940 vss.n2218 vss.n2217 2.703
R59941 vss.n2216 vss.n2215 2.703
R59942 vss.n2260 vss.n2259 2.703
R59943 vss.n2258 vss.n2257 2.703
R59944 vss.n2302 vss.n2301 2.703
R59945 vss.n2300 vss.n2299 2.703
R59946 vss.n2344 vss.n2343 2.703
R59947 vss.n2342 vss.n2341 2.703
R59948 vss.n2386 vss.n2385 2.703
R59949 vss.n2384 vss.n2383 2.703
R59950 vss.n3188 vss.n3183 0.196
R59951 vss.n3191 vss.n3188 0.195
R59952 vss.n3196 vss.n3191 0.195
R59953 vss.n3197 vss.n3196 0.193
R59954 vss.n2401 vss.n2396 0.17
R59955 vss.n2404 vss.n2401 0.169
R59956 vss.n2409 vss.n2404 0.169
R59957 vss.n2410 vss.n2409 0.152
R59958 vss.n3169 vss.n3159 0.144
R59959 vss.n3179 vss.n3169 0.144
R59960 vss.n3180 vss.n3179 0.144
R59961 vss.n3127 vss.n3117 0.144
R59962 vss.n3137 vss.n3127 0.144
R59963 vss.n3138 vss.n3137 0.144
R59964 vss.n3085 vss.n3075 0.144
R59965 vss.n3095 vss.n3085 0.144
R59966 vss.n3096 vss.n3095 0.144
R59967 vss.n3043 vss.n3033 0.144
R59968 vss.n3053 vss.n3043 0.144
R59969 vss.n3054 vss.n3053 0.144
R59970 vss.n3001 vss.n2991 0.144
R59971 vss.n3011 vss.n3001 0.144
R59972 vss.n3012 vss.n3011 0.144
R59973 vss.n2959 vss.n2949 0.144
R59974 vss.n2969 vss.n2959 0.144
R59975 vss.n2970 vss.n2969 0.144
R59976 vss.n2917 vss.n2907 0.144
R59977 vss.n2927 vss.n2917 0.144
R59978 vss.n2928 vss.n2927 0.144
R59979 vss.n2875 vss.n2865 0.144
R59980 vss.n2885 vss.n2875 0.144
R59981 vss.n2886 vss.n2885 0.144
R59982 vss.n2833 vss.n2823 0.144
R59983 vss.n2843 vss.n2833 0.144
R59984 vss.n2844 vss.n2843 0.144
R59985 vss.n2791 vss.n2781 0.144
R59986 vss.n2801 vss.n2791 0.144
R59987 vss.n2802 vss.n2801 0.144
R59988 vss.n2749 vss.n2739 0.144
R59989 vss.n2759 vss.n2749 0.144
R59990 vss.n2760 vss.n2759 0.144
R59991 vss.n2707 vss.n2697 0.144
R59992 vss.n2717 vss.n2707 0.144
R59993 vss.n2718 vss.n2717 0.144
R59994 vss.n2665 vss.n2655 0.144
R59995 vss.n2675 vss.n2665 0.144
R59996 vss.n2676 vss.n2675 0.144
R59997 vss.n2623 vss.n2613 0.144
R59998 vss.n2633 vss.n2623 0.144
R59999 vss.n2634 vss.n2633 0.144
R60000 vss.n2581 vss.n2571 0.144
R60001 vss.n2591 vss.n2581 0.144
R60002 vss.n2592 vss.n2591 0.144
R60003 vss.n2539 vss.n2529 0.144
R60004 vss.n2549 vss.n2539 0.144
R60005 vss.n2550 vss.n2549 0.144
R60006 vss.n2497 vss.n2487 0.144
R60007 vss.n2507 vss.n2497 0.144
R60008 vss.n2508 vss.n2507 0.144
R60009 vss.n30 vss.n20 0.144
R60010 vss.n40 vss.n30 0.144
R60011 vss.n41 vss.n40 0.144
R60012 vss.n72 vss.n62 0.144
R60013 vss.n82 vss.n72 0.144
R60014 vss.n83 vss.n82 0.144
R60015 vss.n114 vss.n104 0.144
R60016 vss.n124 vss.n114 0.144
R60017 vss.n125 vss.n124 0.144
R60018 vss.n156 vss.n146 0.144
R60019 vss.n166 vss.n156 0.144
R60020 vss.n167 vss.n166 0.144
R60021 vss.n198 vss.n188 0.144
R60022 vss.n208 vss.n198 0.144
R60023 vss.n209 vss.n208 0.144
R60024 vss.n240 vss.n230 0.144
R60025 vss.n250 vss.n240 0.144
R60026 vss.n251 vss.n250 0.144
R60027 vss.n282 vss.n272 0.144
R60028 vss.n292 vss.n282 0.144
R60029 vss.n293 vss.n292 0.144
R60030 vss.n324 vss.n314 0.144
R60031 vss.n334 vss.n324 0.144
R60032 vss.n335 vss.n334 0.144
R60033 vss.n366 vss.n356 0.144
R60034 vss.n376 vss.n366 0.144
R60035 vss.n377 vss.n376 0.144
R60036 vss.n408 vss.n398 0.144
R60037 vss.n418 vss.n408 0.144
R60038 vss.n419 vss.n418 0.144
R60039 vss.n450 vss.n440 0.144
R60040 vss.n460 vss.n450 0.144
R60041 vss.n461 vss.n460 0.144
R60042 vss.n492 vss.n482 0.144
R60043 vss.n502 vss.n492 0.144
R60044 vss.n503 vss.n502 0.144
R60045 vss.n534 vss.n524 0.144
R60046 vss.n544 vss.n534 0.144
R60047 vss.n545 vss.n544 0.144
R60048 vss.n576 vss.n566 0.144
R60049 vss.n586 vss.n576 0.144
R60050 vss.n587 vss.n586 0.144
R60051 vss.n618 vss.n608 0.144
R60052 vss.n628 vss.n618 0.144
R60053 vss.n629 vss.n628 0.144
R60054 vss.n660 vss.n650 0.144
R60055 vss.n670 vss.n660 0.144
R60056 vss.n671 vss.n670 0.144
R60057 vss.n702 vss.n692 0.144
R60058 vss.n712 vss.n702 0.144
R60059 vss.n713 vss.n712 0.144
R60060 vss.n744 vss.n734 0.144
R60061 vss.n754 vss.n744 0.144
R60062 vss.n755 vss.n754 0.144
R60063 vss.n786 vss.n776 0.144
R60064 vss.n796 vss.n786 0.144
R60065 vss.n797 vss.n796 0.144
R60066 vss.n828 vss.n818 0.144
R60067 vss.n838 vss.n828 0.144
R60068 vss.n839 vss.n838 0.144
R60069 vss.n870 vss.n860 0.144
R60070 vss.n880 vss.n870 0.144
R60071 vss.n881 vss.n880 0.144
R60072 vss.n912 vss.n902 0.144
R60073 vss.n922 vss.n912 0.144
R60074 vss.n923 vss.n922 0.144
R60075 vss.n954 vss.n944 0.144
R60076 vss.n964 vss.n954 0.144
R60077 vss.n965 vss.n964 0.144
R60078 vss.n996 vss.n986 0.144
R60079 vss.n1006 vss.n996 0.144
R60080 vss.n1007 vss.n1006 0.144
R60081 vss.n1038 vss.n1028 0.144
R60082 vss.n1048 vss.n1038 0.144
R60083 vss.n1049 vss.n1048 0.144
R60084 vss.n1080 vss.n1070 0.144
R60085 vss.n1090 vss.n1080 0.144
R60086 vss.n1091 vss.n1090 0.144
R60087 vss.n1122 vss.n1112 0.144
R60088 vss.n1132 vss.n1122 0.144
R60089 vss.n1133 vss.n1132 0.144
R60090 vss.n1164 vss.n1154 0.144
R60091 vss.n1174 vss.n1164 0.144
R60092 vss.n1175 vss.n1174 0.144
R60093 vss.n1206 vss.n1196 0.144
R60094 vss.n1216 vss.n1206 0.144
R60095 vss.n1217 vss.n1216 0.144
R60096 vss.n1248 vss.n1238 0.144
R60097 vss.n1258 vss.n1248 0.144
R60098 vss.n1259 vss.n1258 0.144
R60099 vss.n1290 vss.n1280 0.144
R60100 vss.n1300 vss.n1290 0.144
R60101 vss.n1301 vss.n1300 0.144
R60102 vss.n1332 vss.n1322 0.144
R60103 vss.n1342 vss.n1332 0.144
R60104 vss.n1343 vss.n1342 0.144
R60105 vss.n1374 vss.n1364 0.144
R60106 vss.n1384 vss.n1374 0.144
R60107 vss.n1385 vss.n1384 0.144
R60108 vss.n1416 vss.n1406 0.144
R60109 vss.n1426 vss.n1416 0.144
R60110 vss.n1427 vss.n1426 0.144
R60111 vss.n1458 vss.n1448 0.144
R60112 vss.n1468 vss.n1458 0.144
R60113 vss.n1469 vss.n1468 0.144
R60114 vss.n1500 vss.n1490 0.144
R60115 vss.n1510 vss.n1500 0.144
R60116 vss.n1511 vss.n1510 0.144
R60117 vss.n1542 vss.n1532 0.144
R60118 vss.n1552 vss.n1542 0.144
R60119 vss.n1553 vss.n1552 0.144
R60120 vss.n1584 vss.n1574 0.144
R60121 vss.n1594 vss.n1584 0.144
R60122 vss.n1595 vss.n1594 0.144
R60123 vss.n1626 vss.n1616 0.144
R60124 vss.n1636 vss.n1626 0.144
R60125 vss.n1637 vss.n1636 0.144
R60126 vss.n1668 vss.n1658 0.144
R60127 vss.n1678 vss.n1668 0.144
R60128 vss.n1679 vss.n1678 0.144
R60129 vss.n1710 vss.n1700 0.144
R60130 vss.n1720 vss.n1710 0.144
R60131 vss.n1721 vss.n1720 0.144
R60132 vss.n1752 vss.n1742 0.144
R60133 vss.n1762 vss.n1752 0.144
R60134 vss.n1763 vss.n1762 0.144
R60135 vss.n1794 vss.n1784 0.144
R60136 vss.n1804 vss.n1794 0.144
R60137 vss.n1805 vss.n1804 0.144
R60138 vss.n1836 vss.n1826 0.144
R60139 vss.n1846 vss.n1836 0.144
R60140 vss.n1847 vss.n1846 0.144
R60141 vss.n1878 vss.n1868 0.144
R60142 vss.n1888 vss.n1878 0.144
R60143 vss.n1889 vss.n1888 0.144
R60144 vss.n1920 vss.n1910 0.144
R60145 vss.n1930 vss.n1920 0.144
R60146 vss.n1931 vss.n1930 0.144
R60147 vss.n1962 vss.n1952 0.144
R60148 vss.n1972 vss.n1962 0.144
R60149 vss.n1973 vss.n1972 0.144
R60150 vss.n2004 vss.n1994 0.144
R60151 vss.n2014 vss.n2004 0.144
R60152 vss.n2015 vss.n2014 0.144
R60153 vss.n2046 vss.n2036 0.144
R60154 vss.n2056 vss.n2046 0.144
R60155 vss.n2057 vss.n2056 0.144
R60156 vss.n2088 vss.n2078 0.144
R60157 vss.n2098 vss.n2088 0.144
R60158 vss.n2099 vss.n2098 0.144
R60159 vss.n2130 vss.n2120 0.144
R60160 vss.n2140 vss.n2130 0.144
R60161 vss.n2141 vss.n2140 0.144
R60162 vss.n2172 vss.n2162 0.144
R60163 vss.n2182 vss.n2172 0.144
R60164 vss.n2183 vss.n2182 0.144
R60165 vss.n2214 vss.n2204 0.144
R60166 vss.n2224 vss.n2214 0.144
R60167 vss.n2225 vss.n2224 0.144
R60168 vss.n2256 vss.n2246 0.144
R60169 vss.n2266 vss.n2256 0.144
R60170 vss.n2267 vss.n2266 0.144
R60171 vss.n2298 vss.n2288 0.144
R60172 vss.n2308 vss.n2298 0.144
R60173 vss.n2309 vss.n2308 0.144
R60174 vss.n2340 vss.n2330 0.144
R60175 vss.n2350 vss.n2340 0.144
R60176 vss.n2351 vss.n2350 0.144
R60177 vss.n2382 vss.n2372 0.144
R60178 vss.n2392 vss.n2382 0.144
R60179 vss.n2393 vss.n2392 0.144
R60180 vss.n3197 vss.n3180 0.13
R60181 vss.n3198 vss.n3138 0.13
R60182 vss.n3199 vss.n3096 0.13
R60183 vss.n3200 vss.n3054 0.13
R60184 vss.n3201 vss.n3012 0.13
R60185 vss.n3202 vss.n2970 0.13
R60186 vss.n3203 vss.n2928 0.13
R60187 vss.n3204 vss.n2886 0.13
R60188 vss.n3205 vss.n2844 0.13
R60189 vss.n3206 vss.n2802 0.13
R60190 vss.n3207 vss.n2760 0.13
R60191 vss.n3208 vss.n2718 0.13
R60192 vss.n3209 vss.n2676 0.13
R60193 vss.n3210 vss.n2634 0.13
R60194 vss.n3211 vss.n2592 0.13
R60195 vss.n3212 vss.n2550 0.13
R60196 vss.n3213 vss.n2508 0.13
R60197 vss.n2466 vss.n41 0.13
R60198 vss.n2465 vss.n83 0.13
R60199 vss.n2464 vss.n125 0.13
R60200 vss.n2463 vss.n167 0.13
R60201 vss.n2462 vss.n209 0.13
R60202 vss.n2461 vss.n251 0.13
R60203 vss.n2460 vss.n293 0.13
R60204 vss.n2459 vss.n335 0.13
R60205 vss.n2458 vss.n377 0.13
R60206 vss.n2457 vss.n419 0.13
R60207 vss.n2456 vss.n461 0.13
R60208 vss.n2455 vss.n503 0.13
R60209 vss.n2454 vss.n545 0.13
R60210 vss.n2453 vss.n587 0.13
R60211 vss.n2452 vss.n629 0.13
R60212 vss.n2451 vss.n671 0.13
R60213 vss.n2450 vss.n713 0.13
R60214 vss.n2449 vss.n755 0.13
R60215 vss.n2448 vss.n797 0.13
R60216 vss.n2447 vss.n839 0.13
R60217 vss.n2446 vss.n881 0.13
R60218 vss.n2445 vss.n923 0.13
R60219 vss.n2444 vss.n965 0.13
R60220 vss.n2443 vss.n1007 0.13
R60221 vss.n2442 vss.n1049 0.13
R60222 vss.n2441 vss.n1091 0.13
R60223 vss.n2440 vss.n1133 0.13
R60224 vss.n2439 vss.n1175 0.13
R60225 vss.n2438 vss.n1217 0.13
R60226 vss.n2437 vss.n1259 0.13
R60227 vss.n2436 vss.n1301 0.13
R60228 vss.n2435 vss.n1343 0.13
R60229 vss.n2434 vss.n1385 0.13
R60230 vss.n2433 vss.n1427 0.13
R60231 vss.n2432 vss.n1469 0.13
R60232 vss.n2431 vss.n1511 0.13
R60233 vss.n2430 vss.n1553 0.13
R60234 vss.n2429 vss.n1595 0.13
R60235 vss.n2428 vss.n1637 0.13
R60236 vss.n2427 vss.n1679 0.13
R60237 vss.n2426 vss.n1721 0.13
R60238 vss.n2425 vss.n1763 0.13
R60239 vss.n2424 vss.n1805 0.13
R60240 vss.n2423 vss.n1847 0.13
R60241 vss.n2422 vss.n1889 0.13
R60242 vss.n2421 vss.n1931 0.13
R60243 vss.n2420 vss.n1973 0.13
R60244 vss.n2419 vss.n2015 0.13
R60245 vss.n2418 vss.n2057 0.13
R60246 vss.n2417 vss.n2099 0.13
R60247 vss.n2416 vss.n2141 0.13
R60248 vss.n2415 vss.n2183 0.13
R60249 vss.n2414 vss.n2225 0.13
R60250 vss.n2413 vss.n2267 0.13
R60251 vss.n2412 vss.n2309 0.13
R60252 vss.n2411 vss.n2351 0.13
R60253 vss.n2410 vss.n2393 0.13
R60254 vss.n3178 vss.n3175 0.011
R60255 vss.n3178 vss.n3177 0.011
R60256 vss.n3168 vss.n3165 0.011
R60257 vss.n3168 vss.n3167 0.011
R60258 vss.n3158 vss.n3155 0.011
R60259 vss.n3158 vss.n3157 0.011
R60260 vss.n3150 vss.n3143 0.011
R60261 vss.n3150 vss.n3144 0.011
R60262 vss.n3136 vss.n3133 0.011
R60263 vss.n3136 vss.n3135 0.011
R60264 vss.n3126 vss.n3123 0.011
R60265 vss.n3126 vss.n3125 0.011
R60266 vss.n3116 vss.n3113 0.011
R60267 vss.n3116 vss.n3115 0.011
R60268 vss.n3108 vss.n3101 0.011
R60269 vss.n3108 vss.n3102 0.011
R60270 vss.n3094 vss.n3091 0.011
R60271 vss.n3094 vss.n3093 0.011
R60272 vss.n3084 vss.n3081 0.011
R60273 vss.n3084 vss.n3083 0.011
R60274 vss.n3074 vss.n3071 0.011
R60275 vss.n3074 vss.n3073 0.011
R60276 vss.n3066 vss.n3059 0.011
R60277 vss.n3066 vss.n3060 0.011
R60278 vss.n3052 vss.n3049 0.011
R60279 vss.n3052 vss.n3051 0.011
R60280 vss.n3042 vss.n3039 0.011
R60281 vss.n3042 vss.n3041 0.011
R60282 vss.n3032 vss.n3029 0.011
R60283 vss.n3032 vss.n3031 0.011
R60284 vss.n3024 vss.n3017 0.011
R60285 vss.n3024 vss.n3018 0.011
R60286 vss.n3010 vss.n3007 0.011
R60287 vss.n3010 vss.n3009 0.011
R60288 vss.n3000 vss.n2997 0.011
R60289 vss.n3000 vss.n2999 0.011
R60290 vss.n2990 vss.n2987 0.011
R60291 vss.n2990 vss.n2989 0.011
R60292 vss.n2982 vss.n2975 0.011
R60293 vss.n2982 vss.n2976 0.011
R60294 vss.n2968 vss.n2965 0.011
R60295 vss.n2968 vss.n2967 0.011
R60296 vss.n2958 vss.n2955 0.011
R60297 vss.n2958 vss.n2957 0.011
R60298 vss.n2948 vss.n2945 0.011
R60299 vss.n2948 vss.n2947 0.011
R60300 vss.n2940 vss.n2933 0.011
R60301 vss.n2940 vss.n2934 0.011
R60302 vss.n2926 vss.n2923 0.011
R60303 vss.n2926 vss.n2925 0.011
R60304 vss.n2916 vss.n2913 0.011
R60305 vss.n2916 vss.n2915 0.011
R60306 vss.n2906 vss.n2903 0.011
R60307 vss.n2906 vss.n2905 0.011
R60308 vss.n2898 vss.n2891 0.011
R60309 vss.n2898 vss.n2892 0.011
R60310 vss.n2884 vss.n2881 0.011
R60311 vss.n2884 vss.n2883 0.011
R60312 vss.n2874 vss.n2871 0.011
R60313 vss.n2874 vss.n2873 0.011
R60314 vss.n2864 vss.n2861 0.011
R60315 vss.n2864 vss.n2863 0.011
R60316 vss.n2856 vss.n2849 0.011
R60317 vss.n2856 vss.n2850 0.011
R60318 vss.n2842 vss.n2839 0.011
R60319 vss.n2842 vss.n2841 0.011
R60320 vss.n2832 vss.n2829 0.011
R60321 vss.n2832 vss.n2831 0.011
R60322 vss.n2822 vss.n2819 0.011
R60323 vss.n2822 vss.n2821 0.011
R60324 vss.n2814 vss.n2807 0.011
R60325 vss.n2814 vss.n2808 0.011
R60326 vss.n2800 vss.n2797 0.011
R60327 vss.n2800 vss.n2799 0.011
R60328 vss.n2790 vss.n2787 0.011
R60329 vss.n2790 vss.n2789 0.011
R60330 vss.n2780 vss.n2777 0.011
R60331 vss.n2780 vss.n2779 0.011
R60332 vss.n2772 vss.n2765 0.011
R60333 vss.n2772 vss.n2766 0.011
R60334 vss.n2758 vss.n2755 0.011
R60335 vss.n2758 vss.n2757 0.011
R60336 vss.n2748 vss.n2745 0.011
R60337 vss.n2748 vss.n2747 0.011
R60338 vss.n2738 vss.n2735 0.011
R60339 vss.n2738 vss.n2737 0.011
R60340 vss.n2730 vss.n2723 0.011
R60341 vss.n2730 vss.n2724 0.011
R60342 vss.n2716 vss.n2713 0.011
R60343 vss.n2716 vss.n2715 0.011
R60344 vss.n2706 vss.n2703 0.011
R60345 vss.n2706 vss.n2705 0.011
R60346 vss.n2696 vss.n2693 0.011
R60347 vss.n2696 vss.n2695 0.011
R60348 vss.n2688 vss.n2681 0.011
R60349 vss.n2688 vss.n2682 0.011
R60350 vss.n2674 vss.n2671 0.011
R60351 vss.n2674 vss.n2673 0.011
R60352 vss.n2664 vss.n2661 0.011
R60353 vss.n2664 vss.n2663 0.011
R60354 vss.n2654 vss.n2651 0.011
R60355 vss.n2654 vss.n2653 0.011
R60356 vss.n2646 vss.n2639 0.011
R60357 vss.n2646 vss.n2640 0.011
R60358 vss.n2632 vss.n2629 0.011
R60359 vss.n2632 vss.n2631 0.011
R60360 vss.n2622 vss.n2619 0.011
R60361 vss.n2622 vss.n2621 0.011
R60362 vss.n2612 vss.n2609 0.011
R60363 vss.n2612 vss.n2611 0.011
R60364 vss.n2604 vss.n2597 0.011
R60365 vss.n2604 vss.n2598 0.011
R60366 vss.n2590 vss.n2587 0.011
R60367 vss.n2590 vss.n2589 0.011
R60368 vss.n2580 vss.n2577 0.011
R60369 vss.n2580 vss.n2579 0.011
R60370 vss.n2570 vss.n2567 0.011
R60371 vss.n2570 vss.n2569 0.011
R60372 vss.n2562 vss.n2555 0.011
R60373 vss.n2562 vss.n2556 0.011
R60374 vss.n2548 vss.n2545 0.011
R60375 vss.n2548 vss.n2547 0.011
R60376 vss.n2538 vss.n2535 0.011
R60377 vss.n2538 vss.n2537 0.011
R60378 vss.n2528 vss.n2525 0.011
R60379 vss.n2528 vss.n2527 0.011
R60380 vss.n2520 vss.n2513 0.011
R60381 vss.n2520 vss.n2514 0.011
R60382 vss.n2506 vss.n2503 0.011
R60383 vss.n2506 vss.n2505 0.011
R60384 vss.n2496 vss.n2493 0.011
R60385 vss.n2496 vss.n2495 0.011
R60386 vss.n2486 vss.n2483 0.011
R60387 vss.n2486 vss.n2485 0.011
R60388 vss.n2478 vss.n2471 0.011
R60389 vss.n2478 vss.n2472 0.011
R60390 vss.n39 vss.n36 0.011
R60391 vss.n39 vss.n38 0.011
R60392 vss.n29 vss.n26 0.011
R60393 vss.n29 vss.n28 0.011
R60394 vss.n19 vss.n16 0.011
R60395 vss.n19 vss.n18 0.011
R60396 vss.n11 vss.n4 0.011
R60397 vss.n11 vss.n5 0.011
R60398 vss.n81 vss.n78 0.011
R60399 vss.n81 vss.n80 0.011
R60400 vss.n71 vss.n68 0.011
R60401 vss.n71 vss.n70 0.011
R60402 vss.n61 vss.n58 0.011
R60403 vss.n61 vss.n60 0.011
R60404 vss.n53 vss.n46 0.011
R60405 vss.n53 vss.n47 0.011
R60406 vss.n123 vss.n120 0.011
R60407 vss.n123 vss.n122 0.011
R60408 vss.n113 vss.n110 0.011
R60409 vss.n113 vss.n112 0.011
R60410 vss.n103 vss.n100 0.011
R60411 vss.n103 vss.n102 0.011
R60412 vss.n95 vss.n88 0.011
R60413 vss.n95 vss.n89 0.011
R60414 vss.n165 vss.n162 0.011
R60415 vss.n165 vss.n164 0.011
R60416 vss.n155 vss.n152 0.011
R60417 vss.n155 vss.n154 0.011
R60418 vss.n145 vss.n142 0.011
R60419 vss.n145 vss.n144 0.011
R60420 vss.n137 vss.n130 0.011
R60421 vss.n137 vss.n131 0.011
R60422 vss.n207 vss.n204 0.011
R60423 vss.n207 vss.n206 0.011
R60424 vss.n197 vss.n194 0.011
R60425 vss.n197 vss.n196 0.011
R60426 vss.n187 vss.n184 0.011
R60427 vss.n187 vss.n186 0.011
R60428 vss.n179 vss.n172 0.011
R60429 vss.n179 vss.n173 0.011
R60430 vss.n249 vss.n246 0.011
R60431 vss.n249 vss.n248 0.011
R60432 vss.n239 vss.n236 0.011
R60433 vss.n239 vss.n238 0.011
R60434 vss.n229 vss.n226 0.011
R60435 vss.n229 vss.n228 0.011
R60436 vss.n221 vss.n214 0.011
R60437 vss.n221 vss.n215 0.011
R60438 vss.n291 vss.n288 0.011
R60439 vss.n291 vss.n290 0.011
R60440 vss.n281 vss.n278 0.011
R60441 vss.n281 vss.n280 0.011
R60442 vss.n271 vss.n268 0.011
R60443 vss.n271 vss.n270 0.011
R60444 vss.n263 vss.n256 0.011
R60445 vss.n263 vss.n257 0.011
R60446 vss.n333 vss.n330 0.011
R60447 vss.n333 vss.n332 0.011
R60448 vss.n323 vss.n320 0.011
R60449 vss.n323 vss.n322 0.011
R60450 vss.n313 vss.n310 0.011
R60451 vss.n313 vss.n312 0.011
R60452 vss.n305 vss.n298 0.011
R60453 vss.n305 vss.n299 0.011
R60454 vss.n375 vss.n372 0.011
R60455 vss.n375 vss.n374 0.011
R60456 vss.n365 vss.n362 0.011
R60457 vss.n365 vss.n364 0.011
R60458 vss.n355 vss.n352 0.011
R60459 vss.n355 vss.n354 0.011
R60460 vss.n347 vss.n340 0.011
R60461 vss.n347 vss.n341 0.011
R60462 vss.n417 vss.n414 0.011
R60463 vss.n417 vss.n416 0.011
R60464 vss.n407 vss.n404 0.011
R60465 vss.n407 vss.n406 0.011
R60466 vss.n397 vss.n394 0.011
R60467 vss.n397 vss.n396 0.011
R60468 vss.n389 vss.n382 0.011
R60469 vss.n389 vss.n383 0.011
R60470 vss.n459 vss.n456 0.011
R60471 vss.n459 vss.n458 0.011
R60472 vss.n449 vss.n446 0.011
R60473 vss.n449 vss.n448 0.011
R60474 vss.n439 vss.n436 0.011
R60475 vss.n439 vss.n438 0.011
R60476 vss.n431 vss.n424 0.011
R60477 vss.n431 vss.n425 0.011
R60478 vss.n501 vss.n498 0.011
R60479 vss.n501 vss.n500 0.011
R60480 vss.n491 vss.n488 0.011
R60481 vss.n491 vss.n490 0.011
R60482 vss.n481 vss.n478 0.011
R60483 vss.n481 vss.n480 0.011
R60484 vss.n473 vss.n466 0.011
R60485 vss.n473 vss.n467 0.011
R60486 vss.n543 vss.n540 0.011
R60487 vss.n543 vss.n542 0.011
R60488 vss.n533 vss.n530 0.011
R60489 vss.n533 vss.n532 0.011
R60490 vss.n523 vss.n520 0.011
R60491 vss.n523 vss.n522 0.011
R60492 vss.n515 vss.n508 0.011
R60493 vss.n515 vss.n509 0.011
R60494 vss.n585 vss.n582 0.011
R60495 vss.n585 vss.n584 0.011
R60496 vss.n575 vss.n572 0.011
R60497 vss.n575 vss.n574 0.011
R60498 vss.n565 vss.n562 0.011
R60499 vss.n565 vss.n564 0.011
R60500 vss.n557 vss.n550 0.011
R60501 vss.n557 vss.n551 0.011
R60502 vss.n627 vss.n624 0.011
R60503 vss.n627 vss.n626 0.011
R60504 vss.n617 vss.n614 0.011
R60505 vss.n617 vss.n616 0.011
R60506 vss.n607 vss.n604 0.011
R60507 vss.n607 vss.n606 0.011
R60508 vss.n599 vss.n592 0.011
R60509 vss.n599 vss.n593 0.011
R60510 vss.n669 vss.n666 0.011
R60511 vss.n669 vss.n668 0.011
R60512 vss.n659 vss.n656 0.011
R60513 vss.n659 vss.n658 0.011
R60514 vss.n649 vss.n646 0.011
R60515 vss.n649 vss.n648 0.011
R60516 vss.n641 vss.n634 0.011
R60517 vss.n641 vss.n635 0.011
R60518 vss.n711 vss.n708 0.011
R60519 vss.n711 vss.n710 0.011
R60520 vss.n701 vss.n698 0.011
R60521 vss.n701 vss.n700 0.011
R60522 vss.n691 vss.n688 0.011
R60523 vss.n691 vss.n690 0.011
R60524 vss.n683 vss.n676 0.011
R60525 vss.n683 vss.n677 0.011
R60526 vss.n753 vss.n750 0.011
R60527 vss.n753 vss.n752 0.011
R60528 vss.n743 vss.n740 0.011
R60529 vss.n743 vss.n742 0.011
R60530 vss.n733 vss.n730 0.011
R60531 vss.n733 vss.n732 0.011
R60532 vss.n725 vss.n718 0.011
R60533 vss.n725 vss.n719 0.011
R60534 vss.n795 vss.n792 0.011
R60535 vss.n795 vss.n794 0.011
R60536 vss.n785 vss.n782 0.011
R60537 vss.n785 vss.n784 0.011
R60538 vss.n775 vss.n772 0.011
R60539 vss.n775 vss.n774 0.011
R60540 vss.n767 vss.n760 0.011
R60541 vss.n767 vss.n761 0.011
R60542 vss.n837 vss.n834 0.011
R60543 vss.n837 vss.n836 0.011
R60544 vss.n827 vss.n824 0.011
R60545 vss.n827 vss.n826 0.011
R60546 vss.n817 vss.n814 0.011
R60547 vss.n817 vss.n816 0.011
R60548 vss.n809 vss.n802 0.011
R60549 vss.n809 vss.n803 0.011
R60550 vss.n879 vss.n876 0.011
R60551 vss.n879 vss.n878 0.011
R60552 vss.n869 vss.n866 0.011
R60553 vss.n869 vss.n868 0.011
R60554 vss.n859 vss.n856 0.011
R60555 vss.n859 vss.n858 0.011
R60556 vss.n851 vss.n844 0.011
R60557 vss.n851 vss.n845 0.011
R60558 vss.n921 vss.n918 0.011
R60559 vss.n921 vss.n920 0.011
R60560 vss.n911 vss.n908 0.011
R60561 vss.n911 vss.n910 0.011
R60562 vss.n901 vss.n898 0.011
R60563 vss.n901 vss.n900 0.011
R60564 vss.n893 vss.n886 0.011
R60565 vss.n893 vss.n887 0.011
R60566 vss.n963 vss.n960 0.011
R60567 vss.n963 vss.n962 0.011
R60568 vss.n953 vss.n950 0.011
R60569 vss.n953 vss.n952 0.011
R60570 vss.n943 vss.n940 0.011
R60571 vss.n943 vss.n942 0.011
R60572 vss.n935 vss.n928 0.011
R60573 vss.n935 vss.n929 0.011
R60574 vss.n1005 vss.n1002 0.011
R60575 vss.n1005 vss.n1004 0.011
R60576 vss.n995 vss.n992 0.011
R60577 vss.n995 vss.n994 0.011
R60578 vss.n985 vss.n982 0.011
R60579 vss.n985 vss.n984 0.011
R60580 vss.n977 vss.n970 0.011
R60581 vss.n977 vss.n971 0.011
R60582 vss.n1047 vss.n1044 0.011
R60583 vss.n1047 vss.n1046 0.011
R60584 vss.n1037 vss.n1034 0.011
R60585 vss.n1037 vss.n1036 0.011
R60586 vss.n1027 vss.n1024 0.011
R60587 vss.n1027 vss.n1026 0.011
R60588 vss.n1019 vss.n1012 0.011
R60589 vss.n1019 vss.n1013 0.011
R60590 vss.n1089 vss.n1086 0.011
R60591 vss.n1089 vss.n1088 0.011
R60592 vss.n1079 vss.n1076 0.011
R60593 vss.n1079 vss.n1078 0.011
R60594 vss.n1069 vss.n1066 0.011
R60595 vss.n1069 vss.n1068 0.011
R60596 vss.n1061 vss.n1054 0.011
R60597 vss.n1061 vss.n1055 0.011
R60598 vss.n1131 vss.n1128 0.011
R60599 vss.n1131 vss.n1130 0.011
R60600 vss.n1121 vss.n1118 0.011
R60601 vss.n1121 vss.n1120 0.011
R60602 vss.n1111 vss.n1108 0.011
R60603 vss.n1111 vss.n1110 0.011
R60604 vss.n1103 vss.n1096 0.011
R60605 vss.n1103 vss.n1097 0.011
R60606 vss.n1173 vss.n1170 0.011
R60607 vss.n1173 vss.n1172 0.011
R60608 vss.n1163 vss.n1160 0.011
R60609 vss.n1163 vss.n1162 0.011
R60610 vss.n1153 vss.n1150 0.011
R60611 vss.n1153 vss.n1152 0.011
R60612 vss.n1145 vss.n1138 0.011
R60613 vss.n1145 vss.n1139 0.011
R60614 vss.n1215 vss.n1212 0.011
R60615 vss.n1215 vss.n1214 0.011
R60616 vss.n1205 vss.n1202 0.011
R60617 vss.n1205 vss.n1204 0.011
R60618 vss.n1195 vss.n1192 0.011
R60619 vss.n1195 vss.n1194 0.011
R60620 vss.n1187 vss.n1180 0.011
R60621 vss.n1187 vss.n1181 0.011
R60622 vss.n1257 vss.n1254 0.011
R60623 vss.n1257 vss.n1256 0.011
R60624 vss.n1247 vss.n1244 0.011
R60625 vss.n1247 vss.n1246 0.011
R60626 vss.n1237 vss.n1234 0.011
R60627 vss.n1237 vss.n1236 0.011
R60628 vss.n1229 vss.n1222 0.011
R60629 vss.n1229 vss.n1223 0.011
R60630 vss.n1299 vss.n1296 0.011
R60631 vss.n1299 vss.n1298 0.011
R60632 vss.n1289 vss.n1286 0.011
R60633 vss.n1289 vss.n1288 0.011
R60634 vss.n1279 vss.n1276 0.011
R60635 vss.n1279 vss.n1278 0.011
R60636 vss.n1271 vss.n1264 0.011
R60637 vss.n1271 vss.n1265 0.011
R60638 vss.n1341 vss.n1338 0.011
R60639 vss.n1341 vss.n1340 0.011
R60640 vss.n1331 vss.n1328 0.011
R60641 vss.n1331 vss.n1330 0.011
R60642 vss.n1321 vss.n1318 0.011
R60643 vss.n1321 vss.n1320 0.011
R60644 vss.n1313 vss.n1306 0.011
R60645 vss.n1313 vss.n1307 0.011
R60646 vss.n1383 vss.n1380 0.011
R60647 vss.n1383 vss.n1382 0.011
R60648 vss.n1373 vss.n1370 0.011
R60649 vss.n1373 vss.n1372 0.011
R60650 vss.n1363 vss.n1360 0.011
R60651 vss.n1363 vss.n1362 0.011
R60652 vss.n1355 vss.n1348 0.011
R60653 vss.n1355 vss.n1349 0.011
R60654 vss.n1425 vss.n1422 0.011
R60655 vss.n1425 vss.n1424 0.011
R60656 vss.n1415 vss.n1412 0.011
R60657 vss.n1415 vss.n1414 0.011
R60658 vss.n1405 vss.n1402 0.011
R60659 vss.n1405 vss.n1404 0.011
R60660 vss.n1397 vss.n1390 0.011
R60661 vss.n1397 vss.n1391 0.011
R60662 vss.n1467 vss.n1464 0.011
R60663 vss.n1467 vss.n1466 0.011
R60664 vss.n1457 vss.n1454 0.011
R60665 vss.n1457 vss.n1456 0.011
R60666 vss.n1447 vss.n1444 0.011
R60667 vss.n1447 vss.n1446 0.011
R60668 vss.n1439 vss.n1432 0.011
R60669 vss.n1439 vss.n1433 0.011
R60670 vss.n1509 vss.n1506 0.011
R60671 vss.n1509 vss.n1508 0.011
R60672 vss.n1499 vss.n1496 0.011
R60673 vss.n1499 vss.n1498 0.011
R60674 vss.n1489 vss.n1486 0.011
R60675 vss.n1489 vss.n1488 0.011
R60676 vss.n1481 vss.n1474 0.011
R60677 vss.n1481 vss.n1475 0.011
R60678 vss.n1551 vss.n1548 0.011
R60679 vss.n1551 vss.n1550 0.011
R60680 vss.n1541 vss.n1538 0.011
R60681 vss.n1541 vss.n1540 0.011
R60682 vss.n1531 vss.n1528 0.011
R60683 vss.n1531 vss.n1530 0.011
R60684 vss.n1523 vss.n1516 0.011
R60685 vss.n1523 vss.n1517 0.011
R60686 vss.n1593 vss.n1590 0.011
R60687 vss.n1593 vss.n1592 0.011
R60688 vss.n1583 vss.n1580 0.011
R60689 vss.n1583 vss.n1582 0.011
R60690 vss.n1573 vss.n1570 0.011
R60691 vss.n1573 vss.n1572 0.011
R60692 vss.n1565 vss.n1558 0.011
R60693 vss.n1565 vss.n1559 0.011
R60694 vss.n1635 vss.n1632 0.011
R60695 vss.n1635 vss.n1634 0.011
R60696 vss.n1625 vss.n1622 0.011
R60697 vss.n1625 vss.n1624 0.011
R60698 vss.n1615 vss.n1612 0.011
R60699 vss.n1615 vss.n1614 0.011
R60700 vss.n1607 vss.n1600 0.011
R60701 vss.n1607 vss.n1601 0.011
R60702 vss.n1677 vss.n1674 0.011
R60703 vss.n1677 vss.n1676 0.011
R60704 vss.n1667 vss.n1664 0.011
R60705 vss.n1667 vss.n1666 0.011
R60706 vss.n1657 vss.n1654 0.011
R60707 vss.n1657 vss.n1656 0.011
R60708 vss.n1649 vss.n1642 0.011
R60709 vss.n1649 vss.n1643 0.011
R60710 vss.n1719 vss.n1716 0.011
R60711 vss.n1719 vss.n1718 0.011
R60712 vss.n1709 vss.n1706 0.011
R60713 vss.n1709 vss.n1708 0.011
R60714 vss.n1699 vss.n1696 0.011
R60715 vss.n1699 vss.n1698 0.011
R60716 vss.n1691 vss.n1684 0.011
R60717 vss.n1691 vss.n1685 0.011
R60718 vss.n1761 vss.n1758 0.011
R60719 vss.n1761 vss.n1760 0.011
R60720 vss.n1751 vss.n1748 0.011
R60721 vss.n1751 vss.n1750 0.011
R60722 vss.n1741 vss.n1738 0.011
R60723 vss.n1741 vss.n1740 0.011
R60724 vss.n1733 vss.n1726 0.011
R60725 vss.n1733 vss.n1727 0.011
R60726 vss.n1803 vss.n1800 0.011
R60727 vss.n1803 vss.n1802 0.011
R60728 vss.n1793 vss.n1790 0.011
R60729 vss.n1793 vss.n1792 0.011
R60730 vss.n1783 vss.n1780 0.011
R60731 vss.n1783 vss.n1782 0.011
R60732 vss.n1775 vss.n1768 0.011
R60733 vss.n1775 vss.n1769 0.011
R60734 vss.n1845 vss.n1842 0.011
R60735 vss.n1845 vss.n1844 0.011
R60736 vss.n1835 vss.n1832 0.011
R60737 vss.n1835 vss.n1834 0.011
R60738 vss.n1825 vss.n1822 0.011
R60739 vss.n1825 vss.n1824 0.011
R60740 vss.n1817 vss.n1810 0.011
R60741 vss.n1817 vss.n1811 0.011
R60742 vss.n1887 vss.n1884 0.011
R60743 vss.n1887 vss.n1886 0.011
R60744 vss.n1877 vss.n1874 0.011
R60745 vss.n1877 vss.n1876 0.011
R60746 vss.n1867 vss.n1864 0.011
R60747 vss.n1867 vss.n1866 0.011
R60748 vss.n1859 vss.n1852 0.011
R60749 vss.n1859 vss.n1853 0.011
R60750 vss.n1929 vss.n1926 0.011
R60751 vss.n1929 vss.n1928 0.011
R60752 vss.n1919 vss.n1916 0.011
R60753 vss.n1919 vss.n1918 0.011
R60754 vss.n1909 vss.n1906 0.011
R60755 vss.n1909 vss.n1908 0.011
R60756 vss.n1901 vss.n1894 0.011
R60757 vss.n1901 vss.n1895 0.011
R60758 vss.n1971 vss.n1968 0.011
R60759 vss.n1971 vss.n1970 0.011
R60760 vss.n1961 vss.n1958 0.011
R60761 vss.n1961 vss.n1960 0.011
R60762 vss.n1951 vss.n1948 0.011
R60763 vss.n1951 vss.n1950 0.011
R60764 vss.n1943 vss.n1936 0.011
R60765 vss.n1943 vss.n1937 0.011
R60766 vss.n2013 vss.n2010 0.011
R60767 vss.n2013 vss.n2012 0.011
R60768 vss.n2003 vss.n2000 0.011
R60769 vss.n2003 vss.n2002 0.011
R60770 vss.n1993 vss.n1990 0.011
R60771 vss.n1993 vss.n1992 0.011
R60772 vss.n1985 vss.n1978 0.011
R60773 vss.n1985 vss.n1979 0.011
R60774 vss.n2055 vss.n2052 0.011
R60775 vss.n2055 vss.n2054 0.011
R60776 vss.n2045 vss.n2042 0.011
R60777 vss.n2045 vss.n2044 0.011
R60778 vss.n2035 vss.n2032 0.011
R60779 vss.n2035 vss.n2034 0.011
R60780 vss.n2027 vss.n2020 0.011
R60781 vss.n2027 vss.n2021 0.011
R60782 vss.n2097 vss.n2094 0.011
R60783 vss.n2097 vss.n2096 0.011
R60784 vss.n2087 vss.n2084 0.011
R60785 vss.n2087 vss.n2086 0.011
R60786 vss.n2077 vss.n2074 0.011
R60787 vss.n2077 vss.n2076 0.011
R60788 vss.n2069 vss.n2062 0.011
R60789 vss.n2069 vss.n2063 0.011
R60790 vss.n2139 vss.n2136 0.011
R60791 vss.n2139 vss.n2138 0.011
R60792 vss.n2129 vss.n2126 0.011
R60793 vss.n2129 vss.n2128 0.011
R60794 vss.n2119 vss.n2116 0.011
R60795 vss.n2119 vss.n2118 0.011
R60796 vss.n2111 vss.n2104 0.011
R60797 vss.n2111 vss.n2105 0.011
R60798 vss.n2181 vss.n2178 0.011
R60799 vss.n2181 vss.n2180 0.011
R60800 vss.n2171 vss.n2168 0.011
R60801 vss.n2171 vss.n2170 0.011
R60802 vss.n2161 vss.n2158 0.011
R60803 vss.n2161 vss.n2160 0.011
R60804 vss.n2153 vss.n2146 0.011
R60805 vss.n2153 vss.n2147 0.011
R60806 vss.n2223 vss.n2220 0.011
R60807 vss.n2223 vss.n2222 0.011
R60808 vss.n2213 vss.n2210 0.011
R60809 vss.n2213 vss.n2212 0.011
R60810 vss.n2203 vss.n2200 0.011
R60811 vss.n2203 vss.n2202 0.011
R60812 vss.n2195 vss.n2188 0.011
R60813 vss.n2195 vss.n2189 0.011
R60814 vss.n2265 vss.n2262 0.011
R60815 vss.n2265 vss.n2264 0.011
R60816 vss.n2255 vss.n2252 0.011
R60817 vss.n2255 vss.n2254 0.011
R60818 vss.n2245 vss.n2242 0.011
R60819 vss.n2245 vss.n2244 0.011
R60820 vss.n2237 vss.n2230 0.011
R60821 vss.n2237 vss.n2231 0.011
R60822 vss.n2307 vss.n2304 0.011
R60823 vss.n2307 vss.n2306 0.011
R60824 vss.n2297 vss.n2294 0.011
R60825 vss.n2297 vss.n2296 0.011
R60826 vss.n2287 vss.n2284 0.011
R60827 vss.n2287 vss.n2286 0.011
R60828 vss.n2279 vss.n2272 0.011
R60829 vss.n2279 vss.n2273 0.011
R60830 vss.n2349 vss.n2346 0.011
R60831 vss.n2349 vss.n2348 0.011
R60832 vss.n2339 vss.n2336 0.011
R60833 vss.n2339 vss.n2338 0.011
R60834 vss.n2329 vss.n2326 0.011
R60835 vss.n2329 vss.n2328 0.011
R60836 vss.n2321 vss.n2314 0.011
R60837 vss.n2321 vss.n2315 0.011
R60838 vss.n2391 vss.n2388 0.011
R60839 vss.n2391 vss.n2390 0.011
R60840 vss.n2381 vss.n2378 0.011
R60841 vss.n2381 vss.n2380 0.011
R60842 vss.n2371 vss.n2368 0.011
R60843 vss.n2371 vss.n2370 0.011
R60844 vss.n2363 vss.n2356 0.011
R60845 vss.n2363 vss.n2357 0.011
R60846 vss.n3183 vss.n3182 0.003
R60847 vss.n2396 vss.n2395 0.003
R60848 vss.n3188 vss.n3187 0.002
R60849 vss.n3191 vss.n3190 0.002
R60850 vss.n3196 vss.n3195 0.002
R60851 vss.n2401 vss.n2400 0.002
R60852 vss.n2404 vss.n2403 0.002
R60853 vss.n2409 vss.n2408 0.002
R60854 vss.n3151 vss.n3150 0.002
R60855 vss.n3109 vss.n3108 0.002
R60856 vss.n3067 vss.n3066 0.002
R60857 vss.n3025 vss.n3024 0.002
R60858 vss.n2983 vss.n2982 0.002
R60859 vss.n2941 vss.n2940 0.002
R60860 vss.n2899 vss.n2898 0.002
R60861 vss.n2857 vss.n2856 0.002
R60862 vss.n2815 vss.n2814 0.002
R60863 vss.n2773 vss.n2772 0.002
R60864 vss.n2731 vss.n2730 0.002
R60865 vss.n2689 vss.n2688 0.002
R60866 vss.n2647 vss.n2646 0.002
R60867 vss.n2605 vss.n2604 0.002
R60868 vss.n2563 vss.n2562 0.002
R60869 vss.n2521 vss.n2520 0.002
R60870 vss.n2479 vss.n2478 0.002
R60871 vss.n12 vss.n11 0.002
R60872 vss.n54 vss.n53 0.002
R60873 vss.n96 vss.n95 0.002
R60874 vss.n138 vss.n137 0.002
R60875 vss.n180 vss.n179 0.002
R60876 vss.n222 vss.n221 0.002
R60877 vss.n264 vss.n263 0.002
R60878 vss.n306 vss.n305 0.002
R60879 vss.n348 vss.n347 0.002
R60880 vss.n390 vss.n389 0.002
R60881 vss.n432 vss.n431 0.002
R60882 vss.n474 vss.n473 0.002
R60883 vss.n516 vss.n515 0.002
R60884 vss.n558 vss.n557 0.002
R60885 vss.n600 vss.n599 0.002
R60886 vss.n642 vss.n641 0.002
R60887 vss.n684 vss.n683 0.002
R60888 vss.n726 vss.n725 0.002
R60889 vss.n768 vss.n767 0.002
R60890 vss.n810 vss.n809 0.002
R60891 vss.n852 vss.n851 0.002
R60892 vss.n894 vss.n893 0.002
R60893 vss.n936 vss.n935 0.002
R60894 vss.n978 vss.n977 0.002
R60895 vss.n1020 vss.n1019 0.002
R60896 vss.n1062 vss.n1061 0.002
R60897 vss.n1104 vss.n1103 0.002
R60898 vss.n1146 vss.n1145 0.002
R60899 vss.n1188 vss.n1187 0.002
R60900 vss.n1230 vss.n1229 0.002
R60901 vss.n1272 vss.n1271 0.002
R60902 vss.n1314 vss.n1313 0.002
R60903 vss.n1356 vss.n1355 0.002
R60904 vss.n1398 vss.n1397 0.002
R60905 vss.n1440 vss.n1439 0.002
R60906 vss.n1482 vss.n1481 0.002
R60907 vss.n1524 vss.n1523 0.002
R60908 vss.n1566 vss.n1565 0.002
R60909 vss.n1608 vss.n1607 0.002
R60910 vss.n1650 vss.n1649 0.002
R60911 vss.n1692 vss.n1691 0.002
R60912 vss.n1734 vss.n1733 0.002
R60913 vss.n1776 vss.n1775 0.002
R60914 vss.n1818 vss.n1817 0.002
R60915 vss.n1860 vss.n1859 0.002
R60916 vss.n1902 vss.n1901 0.002
R60917 vss.n1944 vss.n1943 0.002
R60918 vss.n1986 vss.n1985 0.002
R60919 vss.n2028 vss.n2027 0.002
R60920 vss.n2070 vss.n2069 0.002
R60921 vss.n2112 vss.n2111 0.002
R60922 vss.n2154 vss.n2153 0.002
R60923 vss.n2196 vss.n2195 0.002
R60924 vss.n2238 vss.n2237 0.002
R60925 vss.n2280 vss.n2279 0.002
R60926 vss.n2322 vss.n2321 0.002
R60927 vss.n2364 vss.n2363 0.002
R60928 vss.n2411 vss.n2410 0.002
R60929 vss.n2412 vss.n2411 0.002
R60930 vss.n2413 vss.n2412 0.002
R60931 vss.n2414 vss.n2413 0.002
R60932 vss.n2415 vss.n2414 0.002
R60933 vss.n2416 vss.n2415 0.002
R60934 vss.n2417 vss.n2416 0.002
R60935 vss.n2418 vss.n2417 0.002
R60936 vss.n2419 vss.n2418 0.002
R60937 vss.n2420 vss.n2419 0.002
R60938 vss.n2421 vss.n2420 0.002
R60939 vss.n2422 vss.n2421 0.002
R60940 vss.n2423 vss.n2422 0.002
R60941 vss.n2424 vss.n2423 0.002
R60942 vss.n2425 vss.n2424 0.002
R60943 vss.n2426 vss.n2425 0.002
R60944 vss.n2427 vss.n2426 0.002
R60945 vss.n2428 vss.n2427 0.002
R60946 vss.n2429 vss.n2428 0.002
R60947 vss.n2430 vss.n2429 0.002
R60948 vss.n2431 vss.n2430 0.002
R60949 vss.n2432 vss.n2431 0.002
R60950 vss.n2433 vss.n2432 0.002
R60951 vss.n2434 vss.n2433 0.002
R60952 vss.n2435 vss.n2434 0.002
R60953 vss.n2436 vss.n2435 0.002
R60954 vss.n2437 vss.n2436 0.002
R60955 vss.n2438 vss.n2437 0.002
R60956 vss.n2439 vss.n2438 0.002
R60957 vss.n2440 vss.n2439 0.002
R60958 vss.n2441 vss.n2440 0.002
R60959 vss.n2442 vss.n2441 0.002
R60960 vss.n2443 vss.n2442 0.002
R60961 vss.n2444 vss.n2443 0.002
R60962 vss.n2445 vss.n2444 0.002
R60963 vss.n2446 vss.n2445 0.002
R60964 vss.n2447 vss.n2446 0.002
R60965 vss.n2448 vss.n2447 0.002
R60966 vss.n2449 vss.n2448 0.002
R60967 vss.n2450 vss.n2449 0.002
R60968 vss.n2451 vss.n2450 0.002
R60969 vss.n2452 vss.n2451 0.002
R60970 vss.n2453 vss.n2452 0.002
R60971 vss.n2454 vss.n2453 0.002
R60972 vss.n2455 vss.n2454 0.002
R60973 vss.n2456 vss.n2455 0.002
R60974 vss.n2457 vss.n2456 0.002
R60975 vss.n2458 vss.n2457 0.002
R60976 vss.n2459 vss.n2458 0.002
R60977 vss.n2460 vss.n2459 0.002
R60978 vss.n2461 vss.n2460 0.002
R60979 vss.n2462 vss.n2461 0.002
R60980 vss.n2463 vss.n2462 0.002
R60981 vss.n2464 vss.n2463 0.002
R60982 vss.n2465 vss.n2464 0.002
R60983 vss.n2466 vss.n2465 0.002
R60984 vss.n3213 vss.n3212 0.002
R60985 vss.n3212 vss.n3211 0.002
R60986 vss.n3211 vss.n3210 0.002
R60987 vss.n3210 vss.n3209 0.002
R60988 vss.n3209 vss.n3208 0.002
R60989 vss.n3208 vss.n3207 0.002
R60990 vss.n3207 vss.n3206 0.002
R60991 vss.n3206 vss.n3205 0.002
R60992 vss.n3205 vss.n3204 0.002
R60993 vss.n3204 vss.n3203 0.002
R60994 vss.n3203 vss.n3202 0.002
R60995 vss.n3202 vss.n3201 0.002
R60996 vss.n3201 vss.n3200 0.002
R60997 vss.n3200 vss.n3199 0.002
R60998 vss.n3199 vss.n3198 0.002
R60999 vss.n3198 vss.n3197 0.002
R61000 vss.n3159 vss.n3158 0.002
R61001 vss.n3169 vss.n3168 0.002
R61002 vss.n3179 vss.n3178 0.002
R61003 vss.n3117 vss.n3116 0.002
R61004 vss.n3127 vss.n3126 0.002
R61005 vss.n3137 vss.n3136 0.002
R61006 vss.n3075 vss.n3074 0.002
R61007 vss.n3085 vss.n3084 0.002
R61008 vss.n3095 vss.n3094 0.002
R61009 vss.n3033 vss.n3032 0.002
R61010 vss.n3043 vss.n3042 0.002
R61011 vss.n3053 vss.n3052 0.002
R61012 vss.n2991 vss.n2990 0.002
R61013 vss.n3001 vss.n3000 0.002
R61014 vss.n3011 vss.n3010 0.002
R61015 vss.n2949 vss.n2948 0.002
R61016 vss.n2959 vss.n2958 0.002
R61017 vss.n2969 vss.n2968 0.002
R61018 vss.n2907 vss.n2906 0.002
R61019 vss.n2917 vss.n2916 0.002
R61020 vss.n2927 vss.n2926 0.002
R61021 vss.n2865 vss.n2864 0.002
R61022 vss.n2875 vss.n2874 0.002
R61023 vss.n2885 vss.n2884 0.002
R61024 vss.n2823 vss.n2822 0.002
R61025 vss.n2833 vss.n2832 0.002
R61026 vss.n2843 vss.n2842 0.002
R61027 vss.n2781 vss.n2780 0.002
R61028 vss.n2791 vss.n2790 0.002
R61029 vss.n2801 vss.n2800 0.002
R61030 vss.n2739 vss.n2738 0.002
R61031 vss.n2749 vss.n2748 0.002
R61032 vss.n2759 vss.n2758 0.002
R61033 vss.n2697 vss.n2696 0.002
R61034 vss.n2707 vss.n2706 0.002
R61035 vss.n2717 vss.n2716 0.002
R61036 vss.n2655 vss.n2654 0.002
R61037 vss.n2665 vss.n2664 0.002
R61038 vss.n2675 vss.n2674 0.002
R61039 vss.n2613 vss.n2612 0.002
R61040 vss.n2623 vss.n2622 0.002
R61041 vss.n2633 vss.n2632 0.002
R61042 vss.n2571 vss.n2570 0.002
R61043 vss.n2581 vss.n2580 0.002
R61044 vss.n2591 vss.n2590 0.002
R61045 vss.n2529 vss.n2528 0.002
R61046 vss.n2539 vss.n2538 0.002
R61047 vss.n2549 vss.n2548 0.002
R61048 vss.n2487 vss.n2486 0.002
R61049 vss.n2497 vss.n2496 0.002
R61050 vss.n2507 vss.n2506 0.002
R61051 vss.n20 vss.n19 0.002
R61052 vss.n30 vss.n29 0.002
R61053 vss.n40 vss.n39 0.002
R61054 vss.n62 vss.n61 0.002
R61055 vss.n72 vss.n71 0.002
R61056 vss.n82 vss.n81 0.002
R61057 vss.n104 vss.n103 0.002
R61058 vss.n114 vss.n113 0.002
R61059 vss.n124 vss.n123 0.002
R61060 vss.n146 vss.n145 0.002
R61061 vss.n156 vss.n155 0.002
R61062 vss.n166 vss.n165 0.002
R61063 vss.n188 vss.n187 0.002
R61064 vss.n198 vss.n197 0.002
R61065 vss.n208 vss.n207 0.002
R61066 vss.n230 vss.n229 0.002
R61067 vss.n240 vss.n239 0.002
R61068 vss.n250 vss.n249 0.002
R61069 vss.n272 vss.n271 0.002
R61070 vss.n282 vss.n281 0.002
R61071 vss.n292 vss.n291 0.002
R61072 vss.n314 vss.n313 0.002
R61073 vss.n324 vss.n323 0.002
R61074 vss.n334 vss.n333 0.002
R61075 vss.n356 vss.n355 0.002
R61076 vss.n366 vss.n365 0.002
R61077 vss.n376 vss.n375 0.002
R61078 vss.n398 vss.n397 0.002
R61079 vss.n408 vss.n407 0.002
R61080 vss.n418 vss.n417 0.002
R61081 vss.n440 vss.n439 0.002
R61082 vss.n450 vss.n449 0.002
R61083 vss.n460 vss.n459 0.002
R61084 vss.n482 vss.n481 0.002
R61085 vss.n492 vss.n491 0.002
R61086 vss.n502 vss.n501 0.002
R61087 vss.n524 vss.n523 0.002
R61088 vss.n534 vss.n533 0.002
R61089 vss.n544 vss.n543 0.002
R61090 vss.n566 vss.n565 0.002
R61091 vss.n576 vss.n575 0.002
R61092 vss.n586 vss.n585 0.002
R61093 vss.n608 vss.n607 0.002
R61094 vss.n618 vss.n617 0.002
R61095 vss.n628 vss.n627 0.002
R61096 vss.n650 vss.n649 0.002
R61097 vss.n660 vss.n659 0.002
R61098 vss.n670 vss.n669 0.002
R61099 vss.n692 vss.n691 0.002
R61100 vss.n702 vss.n701 0.002
R61101 vss.n712 vss.n711 0.002
R61102 vss.n734 vss.n733 0.002
R61103 vss.n744 vss.n743 0.002
R61104 vss.n754 vss.n753 0.002
R61105 vss.n776 vss.n775 0.002
R61106 vss.n786 vss.n785 0.002
R61107 vss.n796 vss.n795 0.002
R61108 vss.n818 vss.n817 0.002
R61109 vss.n828 vss.n827 0.002
R61110 vss.n838 vss.n837 0.002
R61111 vss.n860 vss.n859 0.002
R61112 vss.n870 vss.n869 0.002
R61113 vss.n880 vss.n879 0.002
R61114 vss.n902 vss.n901 0.002
R61115 vss.n912 vss.n911 0.002
R61116 vss.n922 vss.n921 0.002
R61117 vss.n944 vss.n943 0.002
R61118 vss.n954 vss.n953 0.002
R61119 vss.n964 vss.n963 0.002
R61120 vss.n986 vss.n985 0.002
R61121 vss.n996 vss.n995 0.002
R61122 vss.n1006 vss.n1005 0.002
R61123 vss.n1028 vss.n1027 0.002
R61124 vss.n1038 vss.n1037 0.002
R61125 vss.n1048 vss.n1047 0.002
R61126 vss.n1070 vss.n1069 0.002
R61127 vss.n1080 vss.n1079 0.002
R61128 vss.n1090 vss.n1089 0.002
R61129 vss.n1112 vss.n1111 0.002
R61130 vss.n1122 vss.n1121 0.002
R61131 vss.n1132 vss.n1131 0.002
R61132 vss.n1154 vss.n1153 0.002
R61133 vss.n1164 vss.n1163 0.002
R61134 vss.n1174 vss.n1173 0.002
R61135 vss.n1196 vss.n1195 0.002
R61136 vss.n1206 vss.n1205 0.002
R61137 vss.n1216 vss.n1215 0.002
R61138 vss.n1238 vss.n1237 0.002
R61139 vss.n1248 vss.n1247 0.002
R61140 vss.n1258 vss.n1257 0.002
R61141 vss.n1280 vss.n1279 0.002
R61142 vss.n1290 vss.n1289 0.002
R61143 vss.n1300 vss.n1299 0.002
R61144 vss.n1322 vss.n1321 0.002
R61145 vss.n1332 vss.n1331 0.002
R61146 vss.n1342 vss.n1341 0.002
R61147 vss.n1364 vss.n1363 0.002
R61148 vss.n1374 vss.n1373 0.002
R61149 vss.n1384 vss.n1383 0.002
R61150 vss.n1406 vss.n1405 0.002
R61151 vss.n1416 vss.n1415 0.002
R61152 vss.n1426 vss.n1425 0.002
R61153 vss.n1448 vss.n1447 0.002
R61154 vss.n1458 vss.n1457 0.002
R61155 vss.n1468 vss.n1467 0.002
R61156 vss.n1490 vss.n1489 0.002
R61157 vss.n1500 vss.n1499 0.002
R61158 vss.n1510 vss.n1509 0.002
R61159 vss.n1532 vss.n1531 0.002
R61160 vss.n1542 vss.n1541 0.002
R61161 vss.n1552 vss.n1551 0.002
R61162 vss.n1574 vss.n1573 0.002
R61163 vss.n1584 vss.n1583 0.002
R61164 vss.n1594 vss.n1593 0.002
R61165 vss.n1616 vss.n1615 0.002
R61166 vss.n1626 vss.n1625 0.002
R61167 vss.n1636 vss.n1635 0.002
R61168 vss.n1658 vss.n1657 0.002
R61169 vss.n1668 vss.n1667 0.002
R61170 vss.n1678 vss.n1677 0.002
R61171 vss.n1700 vss.n1699 0.002
R61172 vss.n1710 vss.n1709 0.002
R61173 vss.n1720 vss.n1719 0.002
R61174 vss.n1742 vss.n1741 0.002
R61175 vss.n1752 vss.n1751 0.002
R61176 vss.n1762 vss.n1761 0.002
R61177 vss.n1784 vss.n1783 0.002
R61178 vss.n1794 vss.n1793 0.002
R61179 vss.n1804 vss.n1803 0.002
R61180 vss.n1826 vss.n1825 0.002
R61181 vss.n1836 vss.n1835 0.002
R61182 vss.n1846 vss.n1845 0.002
R61183 vss.n1868 vss.n1867 0.002
R61184 vss.n1878 vss.n1877 0.002
R61185 vss.n1888 vss.n1887 0.002
R61186 vss.n1910 vss.n1909 0.002
R61187 vss.n1920 vss.n1919 0.002
R61188 vss.n1930 vss.n1929 0.002
R61189 vss.n1952 vss.n1951 0.002
R61190 vss.n1962 vss.n1961 0.002
R61191 vss.n1972 vss.n1971 0.002
R61192 vss.n1994 vss.n1993 0.002
R61193 vss.n2004 vss.n2003 0.002
R61194 vss.n2014 vss.n2013 0.002
R61195 vss.n2036 vss.n2035 0.002
R61196 vss.n2046 vss.n2045 0.002
R61197 vss.n2056 vss.n2055 0.002
R61198 vss.n2078 vss.n2077 0.002
R61199 vss.n2088 vss.n2087 0.002
R61200 vss.n2098 vss.n2097 0.002
R61201 vss.n2120 vss.n2119 0.002
R61202 vss.n2130 vss.n2129 0.002
R61203 vss.n2140 vss.n2139 0.002
R61204 vss.n2162 vss.n2161 0.002
R61205 vss.n2172 vss.n2171 0.002
R61206 vss.n2182 vss.n2181 0.002
R61207 vss.n2204 vss.n2203 0.002
R61208 vss.n2214 vss.n2213 0.002
R61209 vss.n2224 vss.n2223 0.002
R61210 vss.n2246 vss.n2245 0.002
R61211 vss.n2256 vss.n2255 0.002
R61212 vss.n2266 vss.n2265 0.002
R61213 vss.n2288 vss.n2287 0.002
R61214 vss.n2298 vss.n2297 0.002
R61215 vss.n2308 vss.n2307 0.002
R61216 vss.n2330 vss.n2329 0.002
R61217 vss.n2340 vss.n2339 0.002
R61218 vss.n2350 vss.n2349 0.002
R61219 vss.n2372 vss.n2371 0.002
R61220 vss.n2382 vss.n2381 0.002
R61221 vss.n2392 vss.n2391 0.002
R61222 vss.n3193 vss.n3192 0.001
R61223 vss.n3185 vss.n3184 0.001
R61224 vss.n3146 vss.n3145 0.001
R61225 vss.n3148 vss.n3147 0.001
R61226 vss.n3163 vss.n3162 0.001
R61227 vss.n3161 vss.n3160 0.001
R61228 vss.n3104 vss.n3103 0.001
R61229 vss.n3106 vss.n3105 0.001
R61230 vss.n3121 vss.n3120 0.001
R61231 vss.n3119 vss.n3118 0.001
R61232 vss.n3062 vss.n3061 0.001
R61233 vss.n3064 vss.n3063 0.001
R61234 vss.n3079 vss.n3078 0.001
R61235 vss.n3077 vss.n3076 0.001
R61236 vss.n3020 vss.n3019 0.001
R61237 vss.n3022 vss.n3021 0.001
R61238 vss.n3037 vss.n3036 0.001
R61239 vss.n3035 vss.n3034 0.001
R61240 vss.n2978 vss.n2977 0.001
R61241 vss.n2980 vss.n2979 0.001
R61242 vss.n2995 vss.n2994 0.001
R61243 vss.n2993 vss.n2992 0.001
R61244 vss.n2936 vss.n2935 0.001
R61245 vss.n2938 vss.n2937 0.001
R61246 vss.n2953 vss.n2952 0.001
R61247 vss.n2951 vss.n2950 0.001
R61248 vss.n2894 vss.n2893 0.001
R61249 vss.n2896 vss.n2895 0.001
R61250 vss.n2911 vss.n2910 0.001
R61251 vss.n2909 vss.n2908 0.001
R61252 vss.n2852 vss.n2851 0.001
R61253 vss.n2854 vss.n2853 0.001
R61254 vss.n2869 vss.n2868 0.001
R61255 vss.n2867 vss.n2866 0.001
R61256 vss.n2810 vss.n2809 0.001
R61257 vss.n2812 vss.n2811 0.001
R61258 vss.n2827 vss.n2826 0.001
R61259 vss.n2825 vss.n2824 0.001
R61260 vss.n2768 vss.n2767 0.001
R61261 vss.n2770 vss.n2769 0.001
R61262 vss.n2785 vss.n2784 0.001
R61263 vss.n2783 vss.n2782 0.001
R61264 vss.n2726 vss.n2725 0.001
R61265 vss.n2728 vss.n2727 0.001
R61266 vss.n2743 vss.n2742 0.001
R61267 vss.n2741 vss.n2740 0.001
R61268 vss.n2684 vss.n2683 0.001
R61269 vss.n2686 vss.n2685 0.001
R61270 vss.n2701 vss.n2700 0.001
R61271 vss.n2699 vss.n2698 0.001
R61272 vss.n2642 vss.n2641 0.001
R61273 vss.n2644 vss.n2643 0.001
R61274 vss.n2659 vss.n2658 0.001
R61275 vss.n2657 vss.n2656 0.001
R61276 vss.n2600 vss.n2599 0.001
R61277 vss.n2602 vss.n2601 0.001
R61278 vss.n2617 vss.n2616 0.001
R61279 vss.n2615 vss.n2614 0.001
R61280 vss.n2558 vss.n2557 0.001
R61281 vss.n2560 vss.n2559 0.001
R61282 vss.n2575 vss.n2574 0.001
R61283 vss.n2573 vss.n2572 0.001
R61284 vss.n2516 vss.n2515 0.001
R61285 vss.n2518 vss.n2517 0.001
R61286 vss.n2533 vss.n2532 0.001
R61287 vss.n2531 vss.n2530 0.001
R61288 vss.n2474 vss.n2473 0.001
R61289 vss.n2476 vss.n2475 0.001
R61290 vss.n2491 vss.n2490 0.001
R61291 vss.n2489 vss.n2488 0.001
R61292 vss.n7 vss.n6 0.001
R61293 vss.n9 vss.n8 0.001
R61294 vss.n24 vss.n23 0.001
R61295 vss.n22 vss.n21 0.001
R61296 vss.n49 vss.n48 0.001
R61297 vss.n51 vss.n50 0.001
R61298 vss.n66 vss.n65 0.001
R61299 vss.n64 vss.n63 0.001
R61300 vss.n91 vss.n90 0.001
R61301 vss.n93 vss.n92 0.001
R61302 vss.n108 vss.n107 0.001
R61303 vss.n106 vss.n105 0.001
R61304 vss.n133 vss.n132 0.001
R61305 vss.n135 vss.n134 0.001
R61306 vss.n150 vss.n149 0.001
R61307 vss.n148 vss.n147 0.001
R61308 vss.n175 vss.n174 0.001
R61309 vss.n177 vss.n176 0.001
R61310 vss.n192 vss.n191 0.001
R61311 vss.n190 vss.n189 0.001
R61312 vss.n217 vss.n216 0.001
R61313 vss.n219 vss.n218 0.001
R61314 vss.n234 vss.n233 0.001
R61315 vss.n232 vss.n231 0.001
R61316 vss.n259 vss.n258 0.001
R61317 vss.n261 vss.n260 0.001
R61318 vss.n276 vss.n275 0.001
R61319 vss.n274 vss.n273 0.001
R61320 vss.n301 vss.n300 0.001
R61321 vss.n303 vss.n302 0.001
R61322 vss.n318 vss.n317 0.001
R61323 vss.n316 vss.n315 0.001
R61324 vss.n343 vss.n342 0.001
R61325 vss.n345 vss.n344 0.001
R61326 vss.n360 vss.n359 0.001
R61327 vss.n358 vss.n357 0.001
R61328 vss.n385 vss.n384 0.001
R61329 vss.n387 vss.n386 0.001
R61330 vss.n402 vss.n401 0.001
R61331 vss.n400 vss.n399 0.001
R61332 vss.n427 vss.n426 0.001
R61333 vss.n429 vss.n428 0.001
R61334 vss.n444 vss.n443 0.001
R61335 vss.n442 vss.n441 0.001
R61336 vss.n469 vss.n468 0.001
R61337 vss.n471 vss.n470 0.001
R61338 vss.n486 vss.n485 0.001
R61339 vss.n484 vss.n483 0.001
R61340 vss.n511 vss.n510 0.001
R61341 vss.n513 vss.n512 0.001
R61342 vss.n528 vss.n527 0.001
R61343 vss.n526 vss.n525 0.001
R61344 vss.n553 vss.n552 0.001
R61345 vss.n555 vss.n554 0.001
R61346 vss.n570 vss.n569 0.001
R61347 vss.n568 vss.n567 0.001
R61348 vss.n595 vss.n594 0.001
R61349 vss.n597 vss.n596 0.001
R61350 vss.n612 vss.n611 0.001
R61351 vss.n610 vss.n609 0.001
R61352 vss.n637 vss.n636 0.001
R61353 vss.n639 vss.n638 0.001
R61354 vss.n654 vss.n653 0.001
R61355 vss.n652 vss.n651 0.001
R61356 vss.n679 vss.n678 0.001
R61357 vss.n681 vss.n680 0.001
R61358 vss.n696 vss.n695 0.001
R61359 vss.n694 vss.n693 0.001
R61360 vss.n721 vss.n720 0.001
R61361 vss.n723 vss.n722 0.001
R61362 vss.n738 vss.n737 0.001
R61363 vss.n736 vss.n735 0.001
R61364 vss.n763 vss.n762 0.001
R61365 vss.n765 vss.n764 0.001
R61366 vss.n780 vss.n779 0.001
R61367 vss.n778 vss.n777 0.001
R61368 vss.n805 vss.n804 0.001
R61369 vss.n807 vss.n806 0.001
R61370 vss.n822 vss.n821 0.001
R61371 vss.n820 vss.n819 0.001
R61372 vss.n847 vss.n846 0.001
R61373 vss.n849 vss.n848 0.001
R61374 vss.n864 vss.n863 0.001
R61375 vss.n862 vss.n861 0.001
R61376 vss.n889 vss.n888 0.001
R61377 vss.n891 vss.n890 0.001
R61378 vss.n906 vss.n905 0.001
R61379 vss.n904 vss.n903 0.001
R61380 vss.n931 vss.n930 0.001
R61381 vss.n933 vss.n932 0.001
R61382 vss.n948 vss.n947 0.001
R61383 vss.n946 vss.n945 0.001
R61384 vss.n973 vss.n972 0.001
R61385 vss.n975 vss.n974 0.001
R61386 vss.n990 vss.n989 0.001
R61387 vss.n988 vss.n987 0.001
R61388 vss.n1015 vss.n1014 0.001
R61389 vss.n1017 vss.n1016 0.001
R61390 vss.n1032 vss.n1031 0.001
R61391 vss.n1030 vss.n1029 0.001
R61392 vss.n1057 vss.n1056 0.001
R61393 vss.n1059 vss.n1058 0.001
R61394 vss.n1074 vss.n1073 0.001
R61395 vss.n1072 vss.n1071 0.001
R61396 vss.n1099 vss.n1098 0.001
R61397 vss.n1101 vss.n1100 0.001
R61398 vss.n1116 vss.n1115 0.001
R61399 vss.n1114 vss.n1113 0.001
R61400 vss.n1141 vss.n1140 0.001
R61401 vss.n1143 vss.n1142 0.001
R61402 vss.n1158 vss.n1157 0.001
R61403 vss.n1156 vss.n1155 0.001
R61404 vss.n1183 vss.n1182 0.001
R61405 vss.n1185 vss.n1184 0.001
R61406 vss.n1200 vss.n1199 0.001
R61407 vss.n1198 vss.n1197 0.001
R61408 vss.n1225 vss.n1224 0.001
R61409 vss.n1227 vss.n1226 0.001
R61410 vss.n1242 vss.n1241 0.001
R61411 vss.n1240 vss.n1239 0.001
R61412 vss.n1267 vss.n1266 0.001
R61413 vss.n1269 vss.n1268 0.001
R61414 vss.n1284 vss.n1283 0.001
R61415 vss.n1282 vss.n1281 0.001
R61416 vss.n1309 vss.n1308 0.001
R61417 vss.n1311 vss.n1310 0.001
R61418 vss.n1326 vss.n1325 0.001
R61419 vss.n1324 vss.n1323 0.001
R61420 vss.n1351 vss.n1350 0.001
R61421 vss.n1353 vss.n1352 0.001
R61422 vss.n1368 vss.n1367 0.001
R61423 vss.n1366 vss.n1365 0.001
R61424 vss.n1393 vss.n1392 0.001
R61425 vss.n1395 vss.n1394 0.001
R61426 vss.n1410 vss.n1409 0.001
R61427 vss.n1408 vss.n1407 0.001
R61428 vss.n1435 vss.n1434 0.001
R61429 vss.n1437 vss.n1436 0.001
R61430 vss.n1452 vss.n1451 0.001
R61431 vss.n1450 vss.n1449 0.001
R61432 vss.n1477 vss.n1476 0.001
R61433 vss.n1479 vss.n1478 0.001
R61434 vss.n1494 vss.n1493 0.001
R61435 vss.n1492 vss.n1491 0.001
R61436 vss.n1519 vss.n1518 0.001
R61437 vss.n1521 vss.n1520 0.001
R61438 vss.n1536 vss.n1535 0.001
R61439 vss.n1534 vss.n1533 0.001
R61440 vss.n1561 vss.n1560 0.001
R61441 vss.n1563 vss.n1562 0.001
R61442 vss.n1578 vss.n1577 0.001
R61443 vss.n1576 vss.n1575 0.001
R61444 vss.n1603 vss.n1602 0.001
R61445 vss.n1605 vss.n1604 0.001
R61446 vss.n1620 vss.n1619 0.001
R61447 vss.n1618 vss.n1617 0.001
R61448 vss.n1645 vss.n1644 0.001
R61449 vss.n1647 vss.n1646 0.001
R61450 vss.n1662 vss.n1661 0.001
R61451 vss.n1660 vss.n1659 0.001
R61452 vss.n1687 vss.n1686 0.001
R61453 vss.n1689 vss.n1688 0.001
R61454 vss.n1704 vss.n1703 0.001
R61455 vss.n1702 vss.n1701 0.001
R61456 vss.n1729 vss.n1728 0.001
R61457 vss.n1731 vss.n1730 0.001
R61458 vss.n1746 vss.n1745 0.001
R61459 vss.n1744 vss.n1743 0.001
R61460 vss.n1771 vss.n1770 0.001
R61461 vss.n1773 vss.n1772 0.001
R61462 vss.n1788 vss.n1787 0.001
R61463 vss.n1786 vss.n1785 0.001
R61464 vss.n1813 vss.n1812 0.001
R61465 vss.n1815 vss.n1814 0.001
R61466 vss.n1830 vss.n1829 0.001
R61467 vss.n1828 vss.n1827 0.001
R61468 vss.n1855 vss.n1854 0.001
R61469 vss.n1857 vss.n1856 0.001
R61470 vss.n1872 vss.n1871 0.001
R61471 vss.n1870 vss.n1869 0.001
R61472 vss.n1897 vss.n1896 0.001
R61473 vss.n1899 vss.n1898 0.001
R61474 vss.n1914 vss.n1913 0.001
R61475 vss.n1912 vss.n1911 0.001
R61476 vss.n1939 vss.n1938 0.001
R61477 vss.n1941 vss.n1940 0.001
R61478 vss.n1956 vss.n1955 0.001
R61479 vss.n1954 vss.n1953 0.001
R61480 vss.n1981 vss.n1980 0.001
R61481 vss.n1983 vss.n1982 0.001
R61482 vss.n1998 vss.n1997 0.001
R61483 vss.n1996 vss.n1995 0.001
R61484 vss.n2023 vss.n2022 0.001
R61485 vss.n2025 vss.n2024 0.001
R61486 vss.n2040 vss.n2039 0.001
R61487 vss.n2038 vss.n2037 0.001
R61488 vss.n2065 vss.n2064 0.001
R61489 vss.n2067 vss.n2066 0.001
R61490 vss.n2082 vss.n2081 0.001
R61491 vss.n2080 vss.n2079 0.001
R61492 vss.n2107 vss.n2106 0.001
R61493 vss.n2109 vss.n2108 0.001
R61494 vss.n2124 vss.n2123 0.001
R61495 vss.n2122 vss.n2121 0.001
R61496 vss.n2149 vss.n2148 0.001
R61497 vss.n2151 vss.n2150 0.001
R61498 vss.n2166 vss.n2165 0.001
R61499 vss.n2164 vss.n2163 0.001
R61500 vss.n2191 vss.n2190 0.001
R61501 vss.n2193 vss.n2192 0.001
R61502 vss.n2208 vss.n2207 0.001
R61503 vss.n2206 vss.n2205 0.001
R61504 vss.n2233 vss.n2232 0.001
R61505 vss.n2235 vss.n2234 0.001
R61506 vss.n2250 vss.n2249 0.001
R61507 vss.n2248 vss.n2247 0.001
R61508 vss.n2275 vss.n2274 0.001
R61509 vss.n2277 vss.n2276 0.001
R61510 vss.n2292 vss.n2291 0.001
R61511 vss.n2290 vss.n2289 0.001
R61512 vss.n2317 vss.n2316 0.001
R61513 vss.n2319 vss.n2318 0.001
R61514 vss.n2334 vss.n2333 0.001
R61515 vss.n2332 vss.n2331 0.001
R61516 vss.n2359 vss.n2358 0.001
R61517 vss.n2361 vss.n2360 0.001
R61518 vss.n2376 vss.n2375 0.001
R61519 vss.n2374 vss.n2373 0.001
R61520 vss.n2406 vss.n2405 0.001
R61521 vss.n2398 vss.n2397 0.001
R61522 vss vss.n2466 0.001
R61523 vss vss.n3213 0.001
R61524 vss.n3151 vss.n3139 0.001
R61525 vss.n3180 vss.n3151 0.001
R61526 vss.n3109 vss.n3097 0.001
R61527 vss.n3138 vss.n3109 0.001
R61528 vss.n3067 vss.n3055 0.001
R61529 vss.n3096 vss.n3067 0.001
R61530 vss.n3025 vss.n3013 0.001
R61531 vss.n3054 vss.n3025 0.001
R61532 vss.n2983 vss.n2971 0.001
R61533 vss.n3012 vss.n2983 0.001
R61534 vss.n2941 vss.n2929 0.001
R61535 vss.n2970 vss.n2941 0.001
R61536 vss.n2899 vss.n2887 0.001
R61537 vss.n2928 vss.n2899 0.001
R61538 vss.n2857 vss.n2845 0.001
R61539 vss.n2886 vss.n2857 0.001
R61540 vss.n2815 vss.n2803 0.001
R61541 vss.n2844 vss.n2815 0.001
R61542 vss.n2773 vss.n2761 0.001
R61543 vss.n2802 vss.n2773 0.001
R61544 vss.n2731 vss.n2719 0.001
R61545 vss.n2760 vss.n2731 0.001
R61546 vss.n2689 vss.n2677 0.001
R61547 vss.n2718 vss.n2689 0.001
R61548 vss.n2647 vss.n2635 0.001
R61549 vss.n2676 vss.n2647 0.001
R61550 vss.n2605 vss.n2593 0.001
R61551 vss.n2634 vss.n2605 0.001
R61552 vss.n2563 vss.n2551 0.001
R61553 vss.n2592 vss.n2563 0.001
R61554 vss.n2521 vss.n2509 0.001
R61555 vss.n2550 vss.n2521 0.001
R61556 vss.n2479 vss.n2467 0.001
R61557 vss.n2508 vss.n2479 0.001
R61558 vss.n12 vss.n0 0.001
R61559 vss.n41 vss.n12 0.001
R61560 vss.n54 vss.n42 0.001
R61561 vss.n83 vss.n54 0.001
R61562 vss.n96 vss.n84 0.001
R61563 vss.n125 vss.n96 0.001
R61564 vss.n138 vss.n126 0.001
R61565 vss.n167 vss.n138 0.001
R61566 vss.n180 vss.n168 0.001
R61567 vss.n209 vss.n180 0.001
R61568 vss.n222 vss.n210 0.001
R61569 vss.n251 vss.n222 0.001
R61570 vss.n264 vss.n252 0.001
R61571 vss.n293 vss.n264 0.001
R61572 vss.n306 vss.n294 0.001
R61573 vss.n335 vss.n306 0.001
R61574 vss.n348 vss.n336 0.001
R61575 vss.n377 vss.n348 0.001
R61576 vss.n390 vss.n378 0.001
R61577 vss.n419 vss.n390 0.001
R61578 vss.n432 vss.n420 0.001
R61579 vss.n461 vss.n432 0.001
R61580 vss.n474 vss.n462 0.001
R61581 vss.n503 vss.n474 0.001
R61582 vss.n516 vss.n504 0.001
R61583 vss.n545 vss.n516 0.001
R61584 vss.n558 vss.n546 0.001
R61585 vss.n587 vss.n558 0.001
R61586 vss.n600 vss.n588 0.001
R61587 vss.n629 vss.n600 0.001
R61588 vss.n642 vss.n630 0.001
R61589 vss.n671 vss.n642 0.001
R61590 vss.n684 vss.n672 0.001
R61591 vss.n713 vss.n684 0.001
R61592 vss.n726 vss.n714 0.001
R61593 vss.n755 vss.n726 0.001
R61594 vss.n768 vss.n756 0.001
R61595 vss.n797 vss.n768 0.001
R61596 vss.n810 vss.n798 0.001
R61597 vss.n839 vss.n810 0.001
R61598 vss.n852 vss.n840 0.001
R61599 vss.n881 vss.n852 0.001
R61600 vss.n894 vss.n882 0.001
R61601 vss.n923 vss.n894 0.001
R61602 vss.n936 vss.n924 0.001
R61603 vss.n965 vss.n936 0.001
R61604 vss.n978 vss.n966 0.001
R61605 vss.n1007 vss.n978 0.001
R61606 vss.n1020 vss.n1008 0.001
R61607 vss.n1049 vss.n1020 0.001
R61608 vss.n1062 vss.n1050 0.001
R61609 vss.n1091 vss.n1062 0.001
R61610 vss.n1104 vss.n1092 0.001
R61611 vss.n1133 vss.n1104 0.001
R61612 vss.n1146 vss.n1134 0.001
R61613 vss.n1175 vss.n1146 0.001
R61614 vss.n1188 vss.n1176 0.001
R61615 vss.n1217 vss.n1188 0.001
R61616 vss.n1230 vss.n1218 0.001
R61617 vss.n1259 vss.n1230 0.001
R61618 vss.n1272 vss.n1260 0.001
R61619 vss.n1301 vss.n1272 0.001
R61620 vss.n1314 vss.n1302 0.001
R61621 vss.n1343 vss.n1314 0.001
R61622 vss.n1356 vss.n1344 0.001
R61623 vss.n1385 vss.n1356 0.001
R61624 vss.n1398 vss.n1386 0.001
R61625 vss.n1427 vss.n1398 0.001
R61626 vss.n1440 vss.n1428 0.001
R61627 vss.n1469 vss.n1440 0.001
R61628 vss.n1482 vss.n1470 0.001
R61629 vss.n1511 vss.n1482 0.001
R61630 vss.n1524 vss.n1512 0.001
R61631 vss.n1553 vss.n1524 0.001
R61632 vss.n1566 vss.n1554 0.001
R61633 vss.n1595 vss.n1566 0.001
R61634 vss.n1608 vss.n1596 0.001
R61635 vss.n1637 vss.n1608 0.001
R61636 vss.n1650 vss.n1638 0.001
R61637 vss.n1679 vss.n1650 0.001
R61638 vss.n1692 vss.n1680 0.001
R61639 vss.n1721 vss.n1692 0.001
R61640 vss.n1734 vss.n1722 0.001
R61641 vss.n1763 vss.n1734 0.001
R61642 vss.n1776 vss.n1764 0.001
R61643 vss.n1805 vss.n1776 0.001
R61644 vss.n1818 vss.n1806 0.001
R61645 vss.n1847 vss.n1818 0.001
R61646 vss.n1860 vss.n1848 0.001
R61647 vss.n1889 vss.n1860 0.001
R61648 vss.n1902 vss.n1890 0.001
R61649 vss.n1931 vss.n1902 0.001
R61650 vss.n1944 vss.n1932 0.001
R61651 vss.n1973 vss.n1944 0.001
R61652 vss.n1986 vss.n1974 0.001
R61653 vss.n2015 vss.n1986 0.001
R61654 vss.n2028 vss.n2016 0.001
R61655 vss.n2057 vss.n2028 0.001
R61656 vss.n2070 vss.n2058 0.001
R61657 vss.n2099 vss.n2070 0.001
R61658 vss.n2112 vss.n2100 0.001
R61659 vss.n2141 vss.n2112 0.001
R61660 vss.n2154 vss.n2142 0.001
R61661 vss.n2183 vss.n2154 0.001
R61662 vss.n2196 vss.n2184 0.001
R61663 vss.n2225 vss.n2196 0.001
R61664 vss.n2238 vss.n2226 0.001
R61665 vss.n2267 vss.n2238 0.001
R61666 vss.n2280 vss.n2268 0.001
R61667 vss.n2309 vss.n2280 0.001
R61668 vss.n2322 vss.n2310 0.001
R61669 vss.n2351 vss.n2322 0.001
R61670 vss.n2364 vss.n2352 0.001
R61671 vss.n2393 vss.n2364 0.001
R61672 vss.n3187 vss.n3186 0.001
R61673 vss.n3190 vss.n3189 0.001
R61674 vss.n2400 vss.n2399 0.001
R61675 vss.n2403 vss.n2402 0.001
R61676 vss.n3195 vss.n3194 0.001
R61677 vss.n3182 vss.n3181 0.001
R61678 vss.n2408 vss.n2407 0.001
R61679 vss.n2395 vss.n2394 0.001
C4 vp_n vss 781.08fF
C5 out_p vss 1431.15fF
C6 vp_p vss 1012.73fF
C7 vdd vss 6229.81fF
C8 vp_n.n0 vss 10.84fF $ **FLOATING
C9 vp_n.n1550 vss 1.43fF $ **FLOATING
C10 vp_n.n1551 vss 15.03fF $ **FLOATING
C11 vp_n.n3151 vss 1.45fF $ **FLOATING
C12 vp_n.n3152 vss 17.74fF $ **FLOATING
C13 vp_n.n3153 vss 10.13fF $ **FLOATING
C14 vp_n.n3203 vss 1.43fF $ **FLOATING
C15 vp_n.n3204 vss 15.03fF $ **FLOATING
C16 vp_n.n4804 vss 1.45fF $ **FLOATING
C17 vp_n.n4805 vss 14.22fF $ **FLOATING
C18 vdd.n145 vss 5.17fF $ **FLOATING
C19 vdd.n146 vss 5.17fF $ **FLOATING
C20 vdd.n150 vss 7.24fF $ **FLOATING
C21 vdd.n151 vss 7.48fF $ **FLOATING
C22 vdd.n152 vss 7.48fF $ **FLOATING
C23 vdd.n153 vss 7.48fF $ **FLOATING
C24 vdd.n154 vss 7.48fF $ **FLOATING
C25 vdd.n155 vss 7.48fF $ **FLOATING
C26 vdd.n156 vss 7.48fF $ **FLOATING
C27 vdd.n157 vss 7.48fF $ **FLOATING
C28 vdd.n158 vss 7.48fF $ **FLOATING
C29 vdd.n159 vss 7.48fF $ **FLOATING
C30 vdd.n160 vss 7.48fF $ **FLOATING
C31 vdd.n161 vss 7.48fF $ **FLOATING
C32 vdd.n162 vss 7.48fF $ **FLOATING
C33 vdd.n163 vss 7.48fF $ **FLOATING
C34 vdd.n164 vss 7.48fF $ **FLOATING
C35 vdd.n165 vss 7.48fF $ **FLOATING
C36 vdd.n166 vss 7.48fF $ **FLOATING
C37 vdd.n167 vss 7.48fF $ **FLOATING
C38 vdd.n168 vss 7.48fF $ **FLOATING
C39 vdd.n176 vss 5.17fF $ **FLOATING
C40 vdd.n177 vss 5.17fF $ **FLOATING
C41 vdd.n179 vss 7.28fF $ **FLOATING
C42 vdd.n325 vss 5.17fF $ **FLOATING
C43 vdd.n326 vss 5.17fF $ **FLOATING
C44 vdd.n330 vss 7.24fF $ **FLOATING
C45 vdd.n331 vss 7.48fF $ **FLOATING
C46 vdd.n332 vss 7.48fF $ **FLOATING
C47 vdd.n333 vss 7.48fF $ **FLOATING
C48 vdd.n334 vss 7.48fF $ **FLOATING
C49 vdd.n335 vss 7.48fF $ **FLOATING
C50 vdd.n336 vss 7.48fF $ **FLOATING
C51 vdd.n337 vss 7.48fF $ **FLOATING
C52 vdd.n338 vss 7.48fF $ **FLOATING
C53 vdd.n339 vss 7.48fF $ **FLOATING
C54 vdd.n340 vss 7.48fF $ **FLOATING
C55 vdd.n341 vss 7.48fF $ **FLOATING
C56 vdd.n342 vss 7.48fF $ **FLOATING
C57 vdd.n343 vss 7.48fF $ **FLOATING
C58 vdd.n344 vss 7.48fF $ **FLOATING
C59 vdd.n345 vss 7.48fF $ **FLOATING
C60 vdd.n346 vss 7.48fF $ **FLOATING
C61 vdd.n347 vss 7.48fF $ **FLOATING
C62 vdd.n348 vss 7.48fF $ **FLOATING
C63 vdd.n356 vss 5.17fF $ **FLOATING
C64 vdd.n357 vss 5.17fF $ **FLOATING
C65 vdd.n359 vss 7.28fF $ **FLOATING
C66 vdd.n505 vss 5.17fF $ **FLOATING
C67 vdd.n506 vss 5.17fF $ **FLOATING
C68 vdd.n510 vss 7.24fF $ **FLOATING
C69 vdd.n511 vss 7.48fF $ **FLOATING
C70 vdd.n512 vss 7.48fF $ **FLOATING
C71 vdd.n513 vss 7.48fF $ **FLOATING
C72 vdd.n514 vss 7.48fF $ **FLOATING
C73 vdd.n515 vss 7.48fF $ **FLOATING
C74 vdd.n516 vss 7.48fF $ **FLOATING
C75 vdd.n517 vss 7.48fF $ **FLOATING
C76 vdd.n518 vss 7.48fF $ **FLOATING
C77 vdd.n519 vss 7.48fF $ **FLOATING
C78 vdd.n520 vss 7.48fF $ **FLOATING
C79 vdd.n521 vss 7.48fF $ **FLOATING
C80 vdd.n522 vss 7.48fF $ **FLOATING
C81 vdd.n523 vss 7.48fF $ **FLOATING
C82 vdd.n524 vss 7.48fF $ **FLOATING
C83 vdd.n525 vss 7.48fF $ **FLOATING
C84 vdd.n526 vss 7.48fF $ **FLOATING
C85 vdd.n527 vss 7.48fF $ **FLOATING
C86 vdd.n528 vss 7.48fF $ **FLOATING
C87 vdd.n536 vss 5.17fF $ **FLOATING
C88 vdd.n537 vss 5.17fF $ **FLOATING
C89 vdd.n539 vss 7.28fF $ **FLOATING
C90 vdd.n685 vss 5.17fF $ **FLOATING
C91 vdd.n686 vss 5.17fF $ **FLOATING
C92 vdd.n690 vss 7.24fF $ **FLOATING
C93 vdd.n691 vss 7.48fF $ **FLOATING
C94 vdd.n692 vss 7.48fF $ **FLOATING
C95 vdd.n693 vss 7.48fF $ **FLOATING
C96 vdd.n694 vss 7.48fF $ **FLOATING
C97 vdd.n695 vss 7.48fF $ **FLOATING
C98 vdd.n696 vss 7.48fF $ **FLOATING
C99 vdd.n697 vss 7.48fF $ **FLOATING
C100 vdd.n698 vss 7.48fF $ **FLOATING
C101 vdd.n699 vss 7.48fF $ **FLOATING
C102 vdd.n700 vss 7.48fF $ **FLOATING
C103 vdd.n701 vss 7.48fF $ **FLOATING
C104 vdd.n702 vss 7.48fF $ **FLOATING
C105 vdd.n703 vss 7.48fF $ **FLOATING
C106 vdd.n704 vss 7.48fF $ **FLOATING
C107 vdd.n705 vss 7.48fF $ **FLOATING
C108 vdd.n706 vss 7.48fF $ **FLOATING
C109 vdd.n707 vss 7.48fF $ **FLOATING
C110 vdd.n708 vss 7.48fF $ **FLOATING
C111 vdd.n716 vss 5.17fF $ **FLOATING
C112 vdd.n717 vss 5.17fF $ **FLOATING
C113 vdd.n719 vss 7.28fF $ **FLOATING
C114 vdd.n865 vss 5.17fF $ **FLOATING
C115 vdd.n866 vss 5.17fF $ **FLOATING
C116 vdd.n870 vss 7.24fF $ **FLOATING
C117 vdd.n871 vss 7.48fF $ **FLOATING
C118 vdd.n872 vss 7.48fF $ **FLOATING
C119 vdd.n873 vss 7.48fF $ **FLOATING
C120 vdd.n874 vss 7.48fF $ **FLOATING
C121 vdd.n875 vss 7.48fF $ **FLOATING
C122 vdd.n876 vss 7.48fF $ **FLOATING
C123 vdd.n877 vss 7.48fF $ **FLOATING
C124 vdd.n878 vss 7.48fF $ **FLOATING
C125 vdd.n879 vss 7.48fF $ **FLOATING
C126 vdd.n880 vss 7.48fF $ **FLOATING
C127 vdd.n881 vss 7.48fF $ **FLOATING
C128 vdd.n882 vss 7.48fF $ **FLOATING
C129 vdd.n883 vss 7.48fF $ **FLOATING
C130 vdd.n884 vss 7.48fF $ **FLOATING
C131 vdd.n885 vss 7.48fF $ **FLOATING
C132 vdd.n886 vss 7.48fF $ **FLOATING
C133 vdd.n887 vss 7.48fF $ **FLOATING
C134 vdd.n888 vss 7.48fF $ **FLOATING
C135 vdd.n896 vss 5.17fF $ **FLOATING
C136 vdd.n897 vss 5.17fF $ **FLOATING
C137 vdd.n899 vss 7.28fF $ **FLOATING
C138 vdd.n1045 vss 5.17fF $ **FLOATING
C139 vdd.n1046 vss 5.17fF $ **FLOATING
C140 vdd.n1050 vss 7.24fF $ **FLOATING
C141 vdd.n1051 vss 7.48fF $ **FLOATING
C142 vdd.n1052 vss 7.48fF $ **FLOATING
C143 vdd.n1053 vss 7.48fF $ **FLOATING
C144 vdd.n1054 vss 7.48fF $ **FLOATING
C145 vdd.n1055 vss 7.48fF $ **FLOATING
C146 vdd.n1056 vss 7.48fF $ **FLOATING
C147 vdd.n1057 vss 7.48fF $ **FLOATING
C148 vdd.n1058 vss 7.48fF $ **FLOATING
C149 vdd.n1059 vss 7.48fF $ **FLOATING
C150 vdd.n1060 vss 7.48fF $ **FLOATING
C151 vdd.n1061 vss 7.48fF $ **FLOATING
C152 vdd.n1062 vss 7.48fF $ **FLOATING
C153 vdd.n1063 vss 7.48fF $ **FLOATING
C154 vdd.n1064 vss 7.48fF $ **FLOATING
C155 vdd.n1065 vss 7.48fF $ **FLOATING
C156 vdd.n1066 vss 7.48fF $ **FLOATING
C157 vdd.n1067 vss 7.48fF $ **FLOATING
C158 vdd.n1068 vss 7.48fF $ **FLOATING
C159 vdd.n1076 vss 5.17fF $ **FLOATING
C160 vdd.n1077 vss 5.17fF $ **FLOATING
C161 vdd.n1079 vss 7.28fF $ **FLOATING
C162 vdd.n1225 vss 5.17fF $ **FLOATING
C163 vdd.n1226 vss 5.17fF $ **FLOATING
C164 vdd.n1230 vss 7.24fF $ **FLOATING
C165 vdd.n1231 vss 7.48fF $ **FLOATING
C166 vdd.n1232 vss 7.48fF $ **FLOATING
C167 vdd.n1233 vss 7.48fF $ **FLOATING
C168 vdd.n1234 vss 7.48fF $ **FLOATING
C169 vdd.n1235 vss 7.48fF $ **FLOATING
C170 vdd.n1236 vss 7.48fF $ **FLOATING
C171 vdd.n1237 vss 7.48fF $ **FLOATING
C172 vdd.n1238 vss 7.48fF $ **FLOATING
C173 vdd.n1239 vss 7.48fF $ **FLOATING
C174 vdd.n1240 vss 7.48fF $ **FLOATING
C175 vdd.n1241 vss 7.48fF $ **FLOATING
C176 vdd.n1242 vss 7.48fF $ **FLOATING
C177 vdd.n1243 vss 7.48fF $ **FLOATING
C178 vdd.n1244 vss 7.48fF $ **FLOATING
C179 vdd.n1245 vss 7.48fF $ **FLOATING
C180 vdd.n1246 vss 7.48fF $ **FLOATING
C181 vdd.n1247 vss 7.48fF $ **FLOATING
C182 vdd.n1248 vss 7.48fF $ **FLOATING
C183 vdd.n1256 vss 5.17fF $ **FLOATING
C184 vdd.n1257 vss 5.17fF $ **FLOATING
C185 vdd.n1259 vss 7.28fF $ **FLOATING
C186 vdd.n1405 vss 5.17fF $ **FLOATING
C187 vdd.n1406 vss 5.17fF $ **FLOATING
C188 vdd.n1410 vss 7.24fF $ **FLOATING
C189 vdd.n1411 vss 7.48fF $ **FLOATING
C190 vdd.n1412 vss 7.48fF $ **FLOATING
C191 vdd.n1413 vss 7.48fF $ **FLOATING
C192 vdd.n1414 vss 7.48fF $ **FLOATING
C193 vdd.n1415 vss 7.48fF $ **FLOATING
C194 vdd.n1416 vss 7.48fF $ **FLOATING
C195 vdd.n1417 vss 7.48fF $ **FLOATING
C196 vdd.n1418 vss 7.48fF $ **FLOATING
C197 vdd.n1419 vss 7.48fF $ **FLOATING
C198 vdd.n1420 vss 7.48fF $ **FLOATING
C199 vdd.n1421 vss 7.48fF $ **FLOATING
C200 vdd.n1422 vss 7.48fF $ **FLOATING
C201 vdd.n1423 vss 7.48fF $ **FLOATING
C202 vdd.n1424 vss 7.48fF $ **FLOATING
C203 vdd.n1425 vss 7.48fF $ **FLOATING
C204 vdd.n1426 vss 7.48fF $ **FLOATING
C205 vdd.n1427 vss 7.48fF $ **FLOATING
C206 vdd.n1428 vss 7.48fF $ **FLOATING
C207 vdd.n1436 vss 5.17fF $ **FLOATING
C208 vdd.n1437 vss 5.17fF $ **FLOATING
C209 vdd.n1439 vss 7.28fF $ **FLOATING
C210 vdd.n1585 vss 5.17fF $ **FLOATING
C211 vdd.n1586 vss 5.17fF $ **FLOATING
C212 vdd.n1590 vss 7.24fF $ **FLOATING
C213 vdd.n1591 vss 7.48fF $ **FLOATING
C214 vdd.n1592 vss 7.48fF $ **FLOATING
C215 vdd.n1593 vss 7.48fF $ **FLOATING
C216 vdd.n1594 vss 7.48fF $ **FLOATING
C217 vdd.n1595 vss 7.48fF $ **FLOATING
C218 vdd.n1596 vss 7.48fF $ **FLOATING
C219 vdd.n1597 vss 7.48fF $ **FLOATING
C220 vdd.n1598 vss 7.48fF $ **FLOATING
C221 vdd.n1599 vss 7.48fF $ **FLOATING
C222 vdd.n1600 vss 7.48fF $ **FLOATING
C223 vdd.n1601 vss 7.48fF $ **FLOATING
C224 vdd.n1602 vss 7.48fF $ **FLOATING
C225 vdd.n1603 vss 7.48fF $ **FLOATING
C226 vdd.n1604 vss 7.48fF $ **FLOATING
C227 vdd.n1605 vss 7.48fF $ **FLOATING
C228 vdd.n1606 vss 7.48fF $ **FLOATING
C229 vdd.n1607 vss 7.48fF $ **FLOATING
C230 vdd.n1608 vss 7.48fF $ **FLOATING
C231 vdd.n1616 vss 5.17fF $ **FLOATING
C232 vdd.n1617 vss 5.17fF $ **FLOATING
C233 vdd.n1619 vss 7.28fF $ **FLOATING
C234 vdd.n1765 vss 5.17fF $ **FLOATING
C235 vdd.n1766 vss 5.17fF $ **FLOATING
C236 vdd.n1770 vss 7.24fF $ **FLOATING
C237 vdd.n1771 vss 7.48fF $ **FLOATING
C238 vdd.n1772 vss 7.48fF $ **FLOATING
C239 vdd.n1773 vss 7.48fF $ **FLOATING
C240 vdd.n1774 vss 7.48fF $ **FLOATING
C241 vdd.n1775 vss 7.48fF $ **FLOATING
C242 vdd.n1776 vss 7.48fF $ **FLOATING
C243 vdd.n1777 vss 7.48fF $ **FLOATING
C244 vdd.n1778 vss 7.48fF $ **FLOATING
C245 vdd.n1779 vss 7.48fF $ **FLOATING
C246 vdd.n1780 vss 7.48fF $ **FLOATING
C247 vdd.n1781 vss 7.48fF $ **FLOATING
C248 vdd.n1782 vss 7.48fF $ **FLOATING
C249 vdd.n1783 vss 7.48fF $ **FLOATING
C250 vdd.n1784 vss 7.48fF $ **FLOATING
C251 vdd.n1785 vss 7.48fF $ **FLOATING
C252 vdd.n1786 vss 7.48fF $ **FLOATING
C253 vdd.n1787 vss 7.48fF $ **FLOATING
C254 vdd.n1788 vss 7.48fF $ **FLOATING
C255 vdd.n1796 vss 5.17fF $ **FLOATING
C256 vdd.n1797 vss 5.17fF $ **FLOATING
C257 vdd.n1799 vss 7.28fF $ **FLOATING
C258 vdd.n1945 vss 5.17fF $ **FLOATING
C259 vdd.n1946 vss 5.17fF $ **FLOATING
C260 vdd.n1950 vss 7.24fF $ **FLOATING
C261 vdd.n1951 vss 7.48fF $ **FLOATING
C262 vdd.n1952 vss 7.48fF $ **FLOATING
C263 vdd.n1953 vss 7.48fF $ **FLOATING
C264 vdd.n1954 vss 7.48fF $ **FLOATING
C265 vdd.n1955 vss 7.48fF $ **FLOATING
C266 vdd.n1956 vss 7.48fF $ **FLOATING
C267 vdd.n1957 vss 7.48fF $ **FLOATING
C268 vdd.n1958 vss 7.48fF $ **FLOATING
C269 vdd.n1959 vss 7.48fF $ **FLOATING
C270 vdd.n1960 vss 7.48fF $ **FLOATING
C271 vdd.n1961 vss 7.48fF $ **FLOATING
C272 vdd.n1962 vss 7.48fF $ **FLOATING
C273 vdd.n1963 vss 7.48fF $ **FLOATING
C274 vdd.n1964 vss 7.48fF $ **FLOATING
C275 vdd.n1965 vss 7.48fF $ **FLOATING
C276 vdd.n1966 vss 7.48fF $ **FLOATING
C277 vdd.n1967 vss 7.48fF $ **FLOATING
C278 vdd.n1968 vss 7.48fF $ **FLOATING
C279 vdd.n1976 vss 5.17fF $ **FLOATING
C280 vdd.n1977 vss 5.17fF $ **FLOATING
C281 vdd.n1979 vss 7.28fF $ **FLOATING
C282 vdd.n2125 vss 5.17fF $ **FLOATING
C283 vdd.n2126 vss 5.17fF $ **FLOATING
C284 vdd.n2130 vss 7.24fF $ **FLOATING
C285 vdd.n2131 vss 7.48fF $ **FLOATING
C286 vdd.n2132 vss 7.48fF $ **FLOATING
C287 vdd.n2133 vss 7.48fF $ **FLOATING
C288 vdd.n2134 vss 7.48fF $ **FLOATING
C289 vdd.n2135 vss 7.48fF $ **FLOATING
C290 vdd.n2136 vss 7.48fF $ **FLOATING
C291 vdd.n2137 vss 7.48fF $ **FLOATING
C292 vdd.n2138 vss 7.48fF $ **FLOATING
C293 vdd.n2139 vss 7.48fF $ **FLOATING
C294 vdd.n2140 vss 7.48fF $ **FLOATING
C295 vdd.n2141 vss 7.48fF $ **FLOATING
C296 vdd.n2142 vss 7.48fF $ **FLOATING
C297 vdd.n2143 vss 7.48fF $ **FLOATING
C298 vdd.n2144 vss 7.48fF $ **FLOATING
C299 vdd.n2145 vss 7.48fF $ **FLOATING
C300 vdd.n2146 vss 7.48fF $ **FLOATING
C301 vdd.n2147 vss 7.48fF $ **FLOATING
C302 vdd.n2148 vss 7.48fF $ **FLOATING
C303 vdd.n2156 vss 5.17fF $ **FLOATING
C304 vdd.n2157 vss 5.17fF $ **FLOATING
C305 vdd.n2159 vss 7.28fF $ **FLOATING
C306 vdd.n2305 vss 5.17fF $ **FLOATING
C307 vdd.n2306 vss 5.17fF $ **FLOATING
C308 vdd.n2310 vss 7.24fF $ **FLOATING
C309 vdd.n2311 vss 7.48fF $ **FLOATING
C310 vdd.n2312 vss 7.48fF $ **FLOATING
C311 vdd.n2313 vss 7.48fF $ **FLOATING
C312 vdd.n2314 vss 7.48fF $ **FLOATING
C313 vdd.n2315 vss 7.48fF $ **FLOATING
C314 vdd.n2316 vss 7.48fF $ **FLOATING
C315 vdd.n2317 vss 7.48fF $ **FLOATING
C316 vdd.n2318 vss 7.48fF $ **FLOATING
C317 vdd.n2319 vss 7.48fF $ **FLOATING
C318 vdd.n2320 vss 7.48fF $ **FLOATING
C319 vdd.n2321 vss 7.48fF $ **FLOATING
C320 vdd.n2322 vss 7.48fF $ **FLOATING
C321 vdd.n2323 vss 7.48fF $ **FLOATING
C322 vdd.n2324 vss 7.48fF $ **FLOATING
C323 vdd.n2325 vss 7.48fF $ **FLOATING
C324 vdd.n2326 vss 7.48fF $ **FLOATING
C325 vdd.n2327 vss 7.48fF $ **FLOATING
C326 vdd.n2328 vss 7.48fF $ **FLOATING
C327 vdd.n2336 vss 5.17fF $ **FLOATING
C328 vdd.n2337 vss 5.17fF $ **FLOATING
C329 vdd.n2339 vss 7.28fF $ **FLOATING
C330 vdd.n2485 vss 5.17fF $ **FLOATING
C331 vdd.n2486 vss 5.17fF $ **FLOATING
C332 vdd.n2490 vss 7.24fF $ **FLOATING
C333 vdd.n2491 vss 7.48fF $ **FLOATING
C334 vdd.n2492 vss 7.48fF $ **FLOATING
C335 vdd.n2493 vss 7.48fF $ **FLOATING
C336 vdd.n2494 vss 7.48fF $ **FLOATING
C337 vdd.n2495 vss 7.48fF $ **FLOATING
C338 vdd.n2496 vss 7.48fF $ **FLOATING
C339 vdd.n2497 vss 7.48fF $ **FLOATING
C340 vdd.n2498 vss 7.48fF $ **FLOATING
C341 vdd.n2499 vss 7.48fF $ **FLOATING
C342 vdd.n2500 vss 7.48fF $ **FLOATING
C343 vdd.n2501 vss 7.48fF $ **FLOATING
C344 vdd.n2502 vss 7.48fF $ **FLOATING
C345 vdd.n2503 vss 7.48fF $ **FLOATING
C346 vdd.n2504 vss 7.48fF $ **FLOATING
C347 vdd.n2505 vss 7.48fF $ **FLOATING
C348 vdd.n2506 vss 7.48fF $ **FLOATING
C349 vdd.n2507 vss 7.48fF $ **FLOATING
C350 vdd.n2508 vss 7.48fF $ **FLOATING
C351 vdd.n2516 vss 5.17fF $ **FLOATING
C352 vdd.n2517 vss 5.17fF $ **FLOATING
C353 vdd.n2519 vss 7.28fF $ **FLOATING
C354 vdd.n2665 vss 5.17fF $ **FLOATING
C355 vdd.n2666 vss 5.17fF $ **FLOATING
C356 vdd.n2670 vss 7.24fF $ **FLOATING
C357 vdd.n2671 vss 7.48fF $ **FLOATING
C358 vdd.n2672 vss 7.48fF $ **FLOATING
C359 vdd.n2673 vss 7.48fF $ **FLOATING
C360 vdd.n2674 vss 7.48fF $ **FLOATING
C361 vdd.n2675 vss 7.48fF $ **FLOATING
C362 vdd.n2676 vss 7.48fF $ **FLOATING
C363 vdd.n2677 vss 7.48fF $ **FLOATING
C364 vdd.n2678 vss 7.48fF $ **FLOATING
C365 vdd.n2679 vss 7.48fF $ **FLOATING
C366 vdd.n2680 vss 7.48fF $ **FLOATING
C367 vdd.n2681 vss 7.48fF $ **FLOATING
C368 vdd.n2682 vss 7.48fF $ **FLOATING
C369 vdd.n2683 vss 7.48fF $ **FLOATING
C370 vdd.n2684 vss 7.48fF $ **FLOATING
C371 vdd.n2685 vss 7.48fF $ **FLOATING
C372 vdd.n2686 vss 7.48fF $ **FLOATING
C373 vdd.n2687 vss 7.48fF $ **FLOATING
C374 vdd.n2688 vss 7.48fF $ **FLOATING
C375 vdd.n2696 vss 5.17fF $ **FLOATING
C376 vdd.n2697 vss 5.17fF $ **FLOATING
C377 vdd.n2699 vss 7.28fF $ **FLOATING
C378 vdd.n2845 vss 5.17fF $ **FLOATING
C379 vdd.n2846 vss 5.17fF $ **FLOATING
C380 vdd.n2850 vss 7.24fF $ **FLOATING
C381 vdd.n2851 vss 7.48fF $ **FLOATING
C382 vdd.n2852 vss 7.48fF $ **FLOATING
C383 vdd.n2853 vss 7.48fF $ **FLOATING
C384 vdd.n2854 vss 7.48fF $ **FLOATING
C385 vdd.n2855 vss 7.48fF $ **FLOATING
C386 vdd.n2856 vss 7.48fF $ **FLOATING
C387 vdd.n2857 vss 7.48fF $ **FLOATING
C388 vdd.n2858 vss 7.48fF $ **FLOATING
C389 vdd.n2859 vss 7.48fF $ **FLOATING
C390 vdd.n2860 vss 7.48fF $ **FLOATING
C391 vdd.n2861 vss 7.48fF $ **FLOATING
C392 vdd.n2862 vss 7.48fF $ **FLOATING
C393 vdd.n2863 vss 7.48fF $ **FLOATING
C394 vdd.n2864 vss 7.48fF $ **FLOATING
C395 vdd.n2865 vss 7.48fF $ **FLOATING
C396 vdd.n2866 vss 7.48fF $ **FLOATING
C397 vdd.n2867 vss 7.48fF $ **FLOATING
C398 vdd.n2868 vss 7.48fF $ **FLOATING
C399 vdd.n2876 vss 5.17fF $ **FLOATING
C400 vdd.n2877 vss 5.17fF $ **FLOATING
C401 vdd.n2879 vss 7.28fF $ **FLOATING
C402 vdd.n3025 vss 5.17fF $ **FLOATING
C403 vdd.n3026 vss 5.17fF $ **FLOATING
C404 vdd.n3030 vss 7.24fF $ **FLOATING
C405 vdd.n3031 vss 7.48fF $ **FLOATING
C406 vdd.n3032 vss 7.48fF $ **FLOATING
C407 vdd.n3033 vss 7.48fF $ **FLOATING
C408 vdd.n3034 vss 7.48fF $ **FLOATING
C409 vdd.n3035 vss 7.48fF $ **FLOATING
C410 vdd.n3036 vss 7.48fF $ **FLOATING
C411 vdd.n3037 vss 7.48fF $ **FLOATING
C412 vdd.n3038 vss 7.48fF $ **FLOATING
C413 vdd.n3039 vss 7.48fF $ **FLOATING
C414 vdd.n3040 vss 7.48fF $ **FLOATING
C415 vdd.n3041 vss 7.48fF $ **FLOATING
C416 vdd.n3042 vss 7.48fF $ **FLOATING
C417 vdd.n3043 vss 7.48fF $ **FLOATING
C418 vdd.n3044 vss 7.48fF $ **FLOATING
C419 vdd.n3045 vss 7.48fF $ **FLOATING
C420 vdd.n3046 vss 7.48fF $ **FLOATING
C421 vdd.n3047 vss 7.48fF $ **FLOATING
C422 vdd.n3048 vss 7.48fF $ **FLOATING
C423 vdd.n3056 vss 5.17fF $ **FLOATING
C424 vdd.n3057 vss 5.17fF $ **FLOATING
C425 vdd.n3059 vss 7.28fF $ **FLOATING
C426 vdd.n3205 vss 5.17fF $ **FLOATING
C427 vdd.n3206 vss 5.17fF $ **FLOATING
C428 vdd.n3210 vss 7.24fF $ **FLOATING
C429 vdd.n3211 vss 7.48fF $ **FLOATING
C430 vdd.n3212 vss 7.48fF $ **FLOATING
C431 vdd.n3213 vss 7.48fF $ **FLOATING
C432 vdd.n3214 vss 7.48fF $ **FLOATING
C433 vdd.n3215 vss 7.48fF $ **FLOATING
C434 vdd.n3216 vss 7.48fF $ **FLOATING
C435 vdd.n3217 vss 7.48fF $ **FLOATING
C436 vdd.n3218 vss 7.48fF $ **FLOATING
C437 vdd.n3219 vss 7.48fF $ **FLOATING
C438 vdd.n3220 vss 7.48fF $ **FLOATING
C439 vdd.n3221 vss 7.48fF $ **FLOATING
C440 vdd.n3222 vss 7.48fF $ **FLOATING
C441 vdd.n3223 vss 7.48fF $ **FLOATING
C442 vdd.n3224 vss 7.48fF $ **FLOATING
C443 vdd.n3225 vss 7.48fF $ **FLOATING
C444 vdd.n3226 vss 7.48fF $ **FLOATING
C445 vdd.n3227 vss 7.48fF $ **FLOATING
C446 vdd.n3228 vss 7.48fF $ **FLOATING
C447 vdd.n3236 vss 5.17fF $ **FLOATING
C448 vdd.n3237 vss 5.17fF $ **FLOATING
C449 vdd.n3239 vss 7.28fF $ **FLOATING
C450 vdd.n3385 vss 5.17fF $ **FLOATING
C451 vdd.n3386 vss 5.17fF $ **FLOATING
C452 vdd.n3390 vss 7.24fF $ **FLOATING
C453 vdd.n3391 vss 7.48fF $ **FLOATING
C454 vdd.n3392 vss 7.48fF $ **FLOATING
C455 vdd.n3393 vss 7.48fF $ **FLOATING
C456 vdd.n3394 vss 7.48fF $ **FLOATING
C457 vdd.n3395 vss 7.48fF $ **FLOATING
C458 vdd.n3396 vss 7.48fF $ **FLOATING
C459 vdd.n3397 vss 7.48fF $ **FLOATING
C460 vdd.n3398 vss 7.48fF $ **FLOATING
C461 vdd.n3399 vss 7.48fF $ **FLOATING
C462 vdd.n3400 vss 7.48fF $ **FLOATING
C463 vdd.n3401 vss 7.48fF $ **FLOATING
C464 vdd.n3402 vss 7.48fF $ **FLOATING
C465 vdd.n3403 vss 7.48fF $ **FLOATING
C466 vdd.n3404 vss 7.48fF $ **FLOATING
C467 vdd.n3405 vss 7.48fF $ **FLOATING
C468 vdd.n3406 vss 7.48fF $ **FLOATING
C469 vdd.n3407 vss 7.48fF $ **FLOATING
C470 vdd.n3408 vss 7.48fF $ **FLOATING
C471 vdd.n3416 vss 5.17fF $ **FLOATING
C472 vdd.n3417 vss 5.17fF $ **FLOATING
C473 vdd.n3419 vss 7.28fF $ **FLOATING
C474 vdd.n3565 vss 5.17fF $ **FLOATING
C475 vdd.n3566 vss 5.17fF $ **FLOATING
C476 vdd.n3570 vss 7.24fF $ **FLOATING
C477 vdd.n3571 vss 7.48fF $ **FLOATING
C478 vdd.n3572 vss 7.48fF $ **FLOATING
C479 vdd.n3573 vss 7.48fF $ **FLOATING
C480 vdd.n3574 vss 7.48fF $ **FLOATING
C481 vdd.n3575 vss 7.48fF $ **FLOATING
C482 vdd.n3576 vss 7.48fF $ **FLOATING
C483 vdd.n3577 vss 7.48fF $ **FLOATING
C484 vdd.n3578 vss 7.48fF $ **FLOATING
C485 vdd.n3579 vss 7.48fF $ **FLOATING
C486 vdd.n3580 vss 7.48fF $ **FLOATING
C487 vdd.n3581 vss 7.48fF $ **FLOATING
C488 vdd.n3582 vss 7.48fF $ **FLOATING
C489 vdd.n3583 vss 7.48fF $ **FLOATING
C490 vdd.n3584 vss 7.48fF $ **FLOATING
C491 vdd.n3585 vss 7.48fF $ **FLOATING
C492 vdd.n3586 vss 7.48fF $ **FLOATING
C493 vdd.n3587 vss 7.48fF $ **FLOATING
C494 vdd.n3588 vss 7.48fF $ **FLOATING
C495 vdd.n3596 vss 5.17fF $ **FLOATING
C496 vdd.n3597 vss 5.17fF $ **FLOATING
C497 vdd.n3599 vss 7.28fF $ **FLOATING
C498 vdd.n3745 vss 5.17fF $ **FLOATING
C499 vdd.n3746 vss 5.17fF $ **FLOATING
C500 vdd.n3750 vss 7.24fF $ **FLOATING
C501 vdd.n3751 vss 7.48fF $ **FLOATING
C502 vdd.n3752 vss 7.48fF $ **FLOATING
C503 vdd.n3753 vss 7.48fF $ **FLOATING
C504 vdd.n3754 vss 7.48fF $ **FLOATING
C505 vdd.n3755 vss 7.48fF $ **FLOATING
C506 vdd.n3756 vss 7.48fF $ **FLOATING
C507 vdd.n3757 vss 7.48fF $ **FLOATING
C508 vdd.n3758 vss 7.48fF $ **FLOATING
C509 vdd.n3759 vss 7.48fF $ **FLOATING
C510 vdd.n3760 vss 7.48fF $ **FLOATING
C511 vdd.n3761 vss 7.48fF $ **FLOATING
C512 vdd.n3762 vss 7.48fF $ **FLOATING
C513 vdd.n3763 vss 7.48fF $ **FLOATING
C514 vdd.n3764 vss 7.48fF $ **FLOATING
C515 vdd.n3765 vss 7.48fF $ **FLOATING
C516 vdd.n3766 vss 7.48fF $ **FLOATING
C517 vdd.n3767 vss 7.48fF $ **FLOATING
C518 vdd.n3768 vss 7.48fF $ **FLOATING
C519 vdd.n3776 vss 5.17fF $ **FLOATING
C520 vdd.n3777 vss 5.17fF $ **FLOATING
C521 vdd.n3779 vss 7.28fF $ **FLOATING
C522 vdd.n3925 vss 5.17fF $ **FLOATING
C523 vdd.n3926 vss 5.17fF $ **FLOATING
C524 vdd.n3930 vss 7.24fF $ **FLOATING
C525 vdd.n3931 vss 7.48fF $ **FLOATING
C526 vdd.n3932 vss 7.48fF $ **FLOATING
C527 vdd.n3933 vss 7.48fF $ **FLOATING
C528 vdd.n3934 vss 7.48fF $ **FLOATING
C529 vdd.n3935 vss 7.48fF $ **FLOATING
C530 vdd.n3936 vss 7.48fF $ **FLOATING
C531 vdd.n3937 vss 7.48fF $ **FLOATING
C532 vdd.n3938 vss 7.48fF $ **FLOATING
C533 vdd.n3939 vss 7.48fF $ **FLOATING
C534 vdd.n3940 vss 7.48fF $ **FLOATING
C535 vdd.n3941 vss 7.48fF $ **FLOATING
C536 vdd.n3942 vss 7.48fF $ **FLOATING
C537 vdd.n3943 vss 7.48fF $ **FLOATING
C538 vdd.n3944 vss 7.48fF $ **FLOATING
C539 vdd.n3945 vss 7.48fF $ **FLOATING
C540 vdd.n3946 vss 7.48fF $ **FLOATING
C541 vdd.n3947 vss 7.48fF $ **FLOATING
C542 vdd.n3948 vss 7.48fF $ **FLOATING
C543 vdd.n3956 vss 5.17fF $ **FLOATING
C544 vdd.n3957 vss 5.17fF $ **FLOATING
C545 vdd.n3959 vss 7.28fF $ **FLOATING
C546 vdd.n4105 vss 5.17fF $ **FLOATING
C547 vdd.n4106 vss 5.17fF $ **FLOATING
C548 vdd.n4110 vss 7.24fF $ **FLOATING
C549 vdd.n4111 vss 7.48fF $ **FLOATING
C550 vdd.n4112 vss 7.48fF $ **FLOATING
C551 vdd.n4113 vss 7.48fF $ **FLOATING
C552 vdd.n4114 vss 7.48fF $ **FLOATING
C553 vdd.n4115 vss 7.48fF $ **FLOATING
C554 vdd.n4116 vss 7.48fF $ **FLOATING
C555 vdd.n4117 vss 7.48fF $ **FLOATING
C556 vdd.n4118 vss 7.48fF $ **FLOATING
C557 vdd.n4119 vss 7.48fF $ **FLOATING
C558 vdd.n4120 vss 7.48fF $ **FLOATING
C559 vdd.n4121 vss 7.48fF $ **FLOATING
C560 vdd.n4122 vss 7.48fF $ **FLOATING
C561 vdd.n4123 vss 7.48fF $ **FLOATING
C562 vdd.n4124 vss 7.48fF $ **FLOATING
C563 vdd.n4125 vss 7.48fF $ **FLOATING
C564 vdd.n4126 vss 7.48fF $ **FLOATING
C565 vdd.n4127 vss 7.48fF $ **FLOATING
C566 vdd.n4128 vss 7.48fF $ **FLOATING
C567 vdd.n4136 vss 5.17fF $ **FLOATING
C568 vdd.n4137 vss 5.17fF $ **FLOATING
C569 vdd.n4139 vss 7.28fF $ **FLOATING
C570 vdd.n4285 vss 5.17fF $ **FLOATING
C571 vdd.n4286 vss 5.17fF $ **FLOATING
C572 vdd.n4290 vss 7.24fF $ **FLOATING
C573 vdd.n4291 vss 7.48fF $ **FLOATING
C574 vdd.n4292 vss 7.48fF $ **FLOATING
C575 vdd.n4293 vss 7.48fF $ **FLOATING
C576 vdd.n4294 vss 7.48fF $ **FLOATING
C577 vdd.n4295 vss 7.48fF $ **FLOATING
C578 vdd.n4296 vss 7.48fF $ **FLOATING
C579 vdd.n4297 vss 7.48fF $ **FLOATING
C580 vdd.n4298 vss 7.48fF $ **FLOATING
C581 vdd.n4299 vss 7.48fF $ **FLOATING
C582 vdd.n4300 vss 7.48fF $ **FLOATING
C583 vdd.n4301 vss 7.48fF $ **FLOATING
C584 vdd.n4302 vss 7.48fF $ **FLOATING
C585 vdd.n4303 vss 7.48fF $ **FLOATING
C586 vdd.n4304 vss 7.48fF $ **FLOATING
C587 vdd.n4305 vss 7.48fF $ **FLOATING
C588 vdd.n4306 vss 7.48fF $ **FLOATING
C589 vdd.n4307 vss 7.48fF $ **FLOATING
C590 vdd.n4308 vss 7.48fF $ **FLOATING
C591 vdd.n4316 vss 5.17fF $ **FLOATING
C592 vdd.n4317 vss 5.17fF $ **FLOATING
C593 vdd.n4319 vss 7.28fF $ **FLOATING
C594 vdd.n4465 vss 5.17fF $ **FLOATING
C595 vdd.n4466 vss 5.17fF $ **FLOATING
C596 vdd.n4470 vss 7.24fF $ **FLOATING
C597 vdd.n4471 vss 7.48fF $ **FLOATING
C598 vdd.n4472 vss 7.48fF $ **FLOATING
C599 vdd.n4473 vss 7.48fF $ **FLOATING
C600 vdd.n4474 vss 7.48fF $ **FLOATING
C601 vdd.n4475 vss 7.48fF $ **FLOATING
C602 vdd.n4476 vss 7.48fF $ **FLOATING
C603 vdd.n4477 vss 7.48fF $ **FLOATING
C604 vdd.n4478 vss 7.48fF $ **FLOATING
C605 vdd.n4479 vss 7.48fF $ **FLOATING
C606 vdd.n4480 vss 7.48fF $ **FLOATING
C607 vdd.n4481 vss 7.48fF $ **FLOATING
C608 vdd.n4482 vss 7.48fF $ **FLOATING
C609 vdd.n4483 vss 7.48fF $ **FLOATING
C610 vdd.n4484 vss 7.48fF $ **FLOATING
C611 vdd.n4485 vss 7.48fF $ **FLOATING
C612 vdd.n4486 vss 7.48fF $ **FLOATING
C613 vdd.n4487 vss 7.48fF $ **FLOATING
C614 vdd.n4488 vss 7.48fF $ **FLOATING
C615 vdd.n4496 vss 5.17fF $ **FLOATING
C616 vdd.n4497 vss 5.17fF $ **FLOATING
C617 vdd.n4499 vss 7.28fF $ **FLOATING
C618 vdd.n4645 vss 5.17fF $ **FLOATING
C619 vdd.n4646 vss 5.17fF $ **FLOATING
C620 vdd.n4650 vss 7.24fF $ **FLOATING
C621 vdd.n4651 vss 7.48fF $ **FLOATING
C622 vdd.n4652 vss 7.48fF $ **FLOATING
C623 vdd.n4653 vss 7.48fF $ **FLOATING
C624 vdd.n4654 vss 7.48fF $ **FLOATING
C625 vdd.n4655 vss 7.48fF $ **FLOATING
C626 vdd.n4656 vss 7.48fF $ **FLOATING
C627 vdd.n4657 vss 7.48fF $ **FLOATING
C628 vdd.n4658 vss 7.48fF $ **FLOATING
C629 vdd.n4659 vss 7.48fF $ **FLOATING
C630 vdd.n4660 vss 7.48fF $ **FLOATING
C631 vdd.n4661 vss 7.48fF $ **FLOATING
C632 vdd.n4662 vss 7.48fF $ **FLOATING
C633 vdd.n4663 vss 7.48fF $ **FLOATING
C634 vdd.n4664 vss 7.48fF $ **FLOATING
C635 vdd.n4665 vss 7.48fF $ **FLOATING
C636 vdd.n4666 vss 7.48fF $ **FLOATING
C637 vdd.n4667 vss 7.48fF $ **FLOATING
C638 vdd.n4668 vss 7.48fF $ **FLOATING
C639 vdd.n4676 vss 5.17fF $ **FLOATING
C640 vdd.n4677 vss 5.17fF $ **FLOATING
C641 vdd.n4679 vss 7.28fF $ **FLOATING
C642 vdd.n4825 vss 5.17fF $ **FLOATING
C643 vdd.n4826 vss 5.17fF $ **FLOATING
C644 vdd.n4830 vss 7.24fF $ **FLOATING
C645 vdd.n4831 vss 7.48fF $ **FLOATING
C646 vdd.n4832 vss 7.48fF $ **FLOATING
C647 vdd.n4833 vss 7.48fF $ **FLOATING
C648 vdd.n4834 vss 7.48fF $ **FLOATING
C649 vdd.n4835 vss 7.48fF $ **FLOATING
C650 vdd.n4836 vss 7.48fF $ **FLOATING
C651 vdd.n4837 vss 7.48fF $ **FLOATING
C652 vdd.n4838 vss 7.48fF $ **FLOATING
C653 vdd.n4839 vss 7.48fF $ **FLOATING
C654 vdd.n4840 vss 7.48fF $ **FLOATING
C655 vdd.n4841 vss 7.48fF $ **FLOATING
C656 vdd.n4842 vss 7.48fF $ **FLOATING
C657 vdd.n4843 vss 7.48fF $ **FLOATING
C658 vdd.n4844 vss 7.48fF $ **FLOATING
C659 vdd.n4845 vss 7.48fF $ **FLOATING
C660 vdd.n4846 vss 7.48fF $ **FLOATING
C661 vdd.n4847 vss 7.48fF $ **FLOATING
C662 vdd.n4848 vss 7.48fF $ **FLOATING
C663 vdd.n4856 vss 5.17fF $ **FLOATING
C664 vdd.n4857 vss 5.17fF $ **FLOATING
C665 vdd.n4859 vss 7.28fF $ **FLOATING
C666 vdd.n5005 vss 5.17fF $ **FLOATING
C667 vdd.n5006 vss 5.17fF $ **FLOATING
C668 vdd.n5010 vss 7.24fF $ **FLOATING
C669 vdd.n5011 vss 7.48fF $ **FLOATING
C670 vdd.n5012 vss 7.48fF $ **FLOATING
C671 vdd.n5013 vss 7.48fF $ **FLOATING
C672 vdd.n5014 vss 7.48fF $ **FLOATING
C673 vdd.n5015 vss 7.48fF $ **FLOATING
C674 vdd.n5016 vss 7.48fF $ **FLOATING
C675 vdd.n5017 vss 7.48fF $ **FLOATING
C676 vdd.n5018 vss 7.48fF $ **FLOATING
C677 vdd.n5019 vss 7.48fF $ **FLOATING
C678 vdd.n5020 vss 7.48fF $ **FLOATING
C679 vdd.n5021 vss 7.48fF $ **FLOATING
C680 vdd.n5022 vss 7.48fF $ **FLOATING
C681 vdd.n5023 vss 7.48fF $ **FLOATING
C682 vdd.n5024 vss 7.48fF $ **FLOATING
C683 vdd.n5025 vss 7.48fF $ **FLOATING
C684 vdd.n5026 vss 7.48fF $ **FLOATING
C685 vdd.n5027 vss 7.48fF $ **FLOATING
C686 vdd.n5028 vss 7.48fF $ **FLOATING
C687 vdd.n5036 vss 5.17fF $ **FLOATING
C688 vdd.n5037 vss 5.17fF $ **FLOATING
C689 vdd.n5039 vss 7.28fF $ **FLOATING
C690 vdd.n5185 vss 5.17fF $ **FLOATING
C691 vdd.n5186 vss 5.17fF $ **FLOATING
C692 vdd.n5190 vss 7.24fF $ **FLOATING
C693 vdd.n5191 vss 7.48fF $ **FLOATING
C694 vdd.n5192 vss 7.48fF $ **FLOATING
C695 vdd.n5193 vss 7.48fF $ **FLOATING
C696 vdd.n5194 vss 7.48fF $ **FLOATING
C697 vdd.n5195 vss 7.48fF $ **FLOATING
C698 vdd.n5196 vss 7.48fF $ **FLOATING
C699 vdd.n5197 vss 7.48fF $ **FLOATING
C700 vdd.n5198 vss 7.48fF $ **FLOATING
C701 vdd.n5199 vss 7.48fF $ **FLOATING
C702 vdd.n5200 vss 7.48fF $ **FLOATING
C703 vdd.n5201 vss 7.48fF $ **FLOATING
C704 vdd.n5202 vss 7.48fF $ **FLOATING
C705 vdd.n5203 vss 7.48fF $ **FLOATING
C706 vdd.n5204 vss 7.48fF $ **FLOATING
C707 vdd.n5205 vss 7.48fF $ **FLOATING
C708 vdd.n5206 vss 7.48fF $ **FLOATING
C709 vdd.n5207 vss 7.48fF $ **FLOATING
C710 vdd.n5208 vss 7.48fF $ **FLOATING
C711 vdd.n5216 vss 5.17fF $ **FLOATING
C712 vdd.n5217 vss 5.17fF $ **FLOATING
C713 vdd.n5219 vss 7.28fF $ **FLOATING
C714 vdd.n5365 vss 5.17fF $ **FLOATING
C715 vdd.n5366 vss 5.17fF $ **FLOATING
C716 vdd.n5370 vss 7.24fF $ **FLOATING
C717 vdd.n5371 vss 7.48fF $ **FLOATING
C718 vdd.n5372 vss 7.48fF $ **FLOATING
C719 vdd.n5373 vss 7.48fF $ **FLOATING
C720 vdd.n5374 vss 7.48fF $ **FLOATING
C721 vdd.n5375 vss 7.48fF $ **FLOATING
C722 vdd.n5376 vss 7.48fF $ **FLOATING
C723 vdd.n5377 vss 7.48fF $ **FLOATING
C724 vdd.n5378 vss 7.48fF $ **FLOATING
C725 vdd.n5379 vss 7.48fF $ **FLOATING
C726 vdd.n5380 vss 7.48fF $ **FLOATING
C727 vdd.n5381 vss 7.48fF $ **FLOATING
C728 vdd.n5382 vss 7.48fF $ **FLOATING
C729 vdd.n5383 vss 7.48fF $ **FLOATING
C730 vdd.n5384 vss 7.48fF $ **FLOATING
C731 vdd.n5385 vss 7.48fF $ **FLOATING
C732 vdd.n5386 vss 7.48fF $ **FLOATING
C733 vdd.n5387 vss 7.48fF $ **FLOATING
C734 vdd.n5388 vss 7.48fF $ **FLOATING
C735 vdd.n5396 vss 5.17fF $ **FLOATING
C736 vdd.n5397 vss 5.17fF $ **FLOATING
C737 vdd.n5399 vss 7.28fF $ **FLOATING
C738 vdd.n5545 vss 5.17fF $ **FLOATING
C739 vdd.n5546 vss 5.17fF $ **FLOATING
C740 vdd.n5550 vss 7.24fF $ **FLOATING
C741 vdd.n5551 vss 7.48fF $ **FLOATING
C742 vdd.n5552 vss 7.48fF $ **FLOATING
C743 vdd.n5553 vss 7.48fF $ **FLOATING
C744 vdd.n5554 vss 7.48fF $ **FLOATING
C745 vdd.n5555 vss 7.48fF $ **FLOATING
C746 vdd.n5556 vss 7.48fF $ **FLOATING
C747 vdd.n5557 vss 7.48fF $ **FLOATING
C748 vdd.n5558 vss 7.48fF $ **FLOATING
C749 vdd.n5559 vss 7.48fF $ **FLOATING
C750 vdd.n5560 vss 7.48fF $ **FLOATING
C751 vdd.n5561 vss 7.48fF $ **FLOATING
C752 vdd.n5562 vss 7.48fF $ **FLOATING
C753 vdd.n5563 vss 7.48fF $ **FLOATING
C754 vdd.n5564 vss 7.48fF $ **FLOATING
C755 vdd.n5565 vss 7.48fF $ **FLOATING
C756 vdd.n5566 vss 7.48fF $ **FLOATING
C757 vdd.n5567 vss 7.48fF $ **FLOATING
C758 vdd.n5568 vss 7.48fF $ **FLOATING
C759 vdd.n5576 vss 5.17fF $ **FLOATING
C760 vdd.n5577 vss 5.17fF $ **FLOATING
C761 vdd.n5579 vss 7.28fF $ **FLOATING
C762 vdd.n5725 vss 5.17fF $ **FLOATING
C763 vdd.n5726 vss 5.17fF $ **FLOATING
C764 vdd.n5730 vss 7.24fF $ **FLOATING
C765 vdd.n5731 vss 7.48fF $ **FLOATING
C766 vdd.n5732 vss 7.48fF $ **FLOATING
C767 vdd.n5733 vss 7.48fF $ **FLOATING
C768 vdd.n5734 vss 7.48fF $ **FLOATING
C769 vdd.n5735 vss 7.48fF $ **FLOATING
C770 vdd.n5736 vss 7.48fF $ **FLOATING
C771 vdd.n5737 vss 7.48fF $ **FLOATING
C772 vdd.n5738 vss 7.48fF $ **FLOATING
C773 vdd.n5739 vss 7.48fF $ **FLOATING
C774 vdd.n5740 vss 7.48fF $ **FLOATING
C775 vdd.n5741 vss 7.48fF $ **FLOATING
C776 vdd.n5742 vss 7.48fF $ **FLOATING
C777 vdd.n5743 vss 7.48fF $ **FLOATING
C778 vdd.n5744 vss 7.48fF $ **FLOATING
C779 vdd.n5745 vss 7.48fF $ **FLOATING
C780 vdd.n5746 vss 7.48fF $ **FLOATING
C781 vdd.n5747 vss 7.48fF $ **FLOATING
C782 vdd.n5748 vss 7.48fF $ **FLOATING
C783 vdd.n5756 vss 5.17fF $ **FLOATING
C784 vdd.n5757 vss 5.17fF $ **FLOATING
C785 vdd.n5759 vss 7.28fF $ **FLOATING
C786 vdd.n5905 vss 5.17fF $ **FLOATING
C787 vdd.n5906 vss 5.17fF $ **FLOATING
C788 vdd.n5910 vss 7.24fF $ **FLOATING
C789 vdd.n5911 vss 7.48fF $ **FLOATING
C790 vdd.n5912 vss 7.48fF $ **FLOATING
C791 vdd.n5913 vss 7.48fF $ **FLOATING
C792 vdd.n5914 vss 7.48fF $ **FLOATING
C793 vdd.n5915 vss 7.48fF $ **FLOATING
C794 vdd.n5916 vss 7.48fF $ **FLOATING
C795 vdd.n5917 vss 7.48fF $ **FLOATING
C796 vdd.n5918 vss 7.48fF $ **FLOATING
C797 vdd.n5919 vss 7.48fF $ **FLOATING
C798 vdd.n5920 vss 7.48fF $ **FLOATING
C799 vdd.n5921 vss 7.48fF $ **FLOATING
C800 vdd.n5922 vss 7.48fF $ **FLOATING
C801 vdd.n5923 vss 7.48fF $ **FLOATING
C802 vdd.n5924 vss 7.48fF $ **FLOATING
C803 vdd.n5925 vss 7.48fF $ **FLOATING
C804 vdd.n5926 vss 7.48fF $ **FLOATING
C805 vdd.n5927 vss 7.48fF $ **FLOATING
C806 vdd.n5928 vss 7.48fF $ **FLOATING
C807 vdd.n5936 vss 5.17fF $ **FLOATING
C808 vdd.n5937 vss 5.17fF $ **FLOATING
C809 vdd.n5939 vss 7.28fF $ **FLOATING
C810 vdd.n6085 vss 5.17fF $ **FLOATING
C811 vdd.n6086 vss 5.17fF $ **FLOATING
C812 vdd.n6090 vss 7.24fF $ **FLOATING
C813 vdd.n6091 vss 7.48fF $ **FLOATING
C814 vdd.n6092 vss 7.48fF $ **FLOATING
C815 vdd.n6093 vss 7.48fF $ **FLOATING
C816 vdd.n6094 vss 7.48fF $ **FLOATING
C817 vdd.n6095 vss 7.48fF $ **FLOATING
C818 vdd.n6096 vss 7.48fF $ **FLOATING
C819 vdd.n6097 vss 7.48fF $ **FLOATING
C820 vdd.n6098 vss 7.48fF $ **FLOATING
C821 vdd.n6099 vss 7.48fF $ **FLOATING
C822 vdd.n6100 vss 7.48fF $ **FLOATING
C823 vdd.n6101 vss 7.48fF $ **FLOATING
C824 vdd.n6102 vss 7.48fF $ **FLOATING
C825 vdd.n6103 vss 7.48fF $ **FLOATING
C826 vdd.n6104 vss 7.48fF $ **FLOATING
C827 vdd.n6105 vss 7.48fF $ **FLOATING
C828 vdd.n6106 vss 7.48fF $ **FLOATING
C829 vdd.n6107 vss 7.48fF $ **FLOATING
C830 vdd.n6108 vss 7.48fF $ **FLOATING
C831 vdd.n6116 vss 5.17fF $ **FLOATING
C832 vdd.n6117 vss 5.17fF $ **FLOATING
C833 vdd.n6119 vss 7.28fF $ **FLOATING
C834 vdd.n6265 vss 5.17fF $ **FLOATING
C835 vdd.n6266 vss 5.17fF $ **FLOATING
C836 vdd.n6270 vss 7.24fF $ **FLOATING
C837 vdd.n6271 vss 7.48fF $ **FLOATING
C838 vdd.n6272 vss 7.48fF $ **FLOATING
C839 vdd.n6273 vss 7.48fF $ **FLOATING
C840 vdd.n6274 vss 7.48fF $ **FLOATING
C841 vdd.n6275 vss 7.48fF $ **FLOATING
C842 vdd.n6276 vss 7.48fF $ **FLOATING
C843 vdd.n6277 vss 7.48fF $ **FLOATING
C844 vdd.n6278 vss 7.48fF $ **FLOATING
C845 vdd.n6279 vss 7.48fF $ **FLOATING
C846 vdd.n6280 vss 7.48fF $ **FLOATING
C847 vdd.n6281 vss 7.48fF $ **FLOATING
C848 vdd.n6282 vss 7.48fF $ **FLOATING
C849 vdd.n6283 vss 7.48fF $ **FLOATING
C850 vdd.n6284 vss 7.48fF $ **FLOATING
C851 vdd.n6285 vss 7.48fF $ **FLOATING
C852 vdd.n6286 vss 7.48fF $ **FLOATING
C853 vdd.n6287 vss 7.48fF $ **FLOATING
C854 vdd.n6288 vss 7.48fF $ **FLOATING
C855 vdd.n6296 vss 5.17fF $ **FLOATING
C856 vdd.n6297 vss 5.17fF $ **FLOATING
C857 vdd.n6299 vss 7.28fF $ **FLOATING
C858 vdd.n6445 vss 5.17fF $ **FLOATING
C859 vdd.n6446 vss 5.17fF $ **FLOATING
C860 vdd.n6450 vss 7.24fF $ **FLOATING
C861 vdd.n6451 vss 7.48fF $ **FLOATING
C862 vdd.n6452 vss 7.48fF $ **FLOATING
C863 vdd.n6453 vss 7.48fF $ **FLOATING
C864 vdd.n6454 vss 7.48fF $ **FLOATING
C865 vdd.n6455 vss 7.48fF $ **FLOATING
C866 vdd.n6456 vss 7.48fF $ **FLOATING
C867 vdd.n6457 vss 7.48fF $ **FLOATING
C868 vdd.n6458 vss 7.48fF $ **FLOATING
C869 vdd.n6459 vss 7.48fF $ **FLOATING
C870 vdd.n6460 vss 7.48fF $ **FLOATING
C871 vdd.n6461 vss 7.48fF $ **FLOATING
C872 vdd.n6462 vss 7.48fF $ **FLOATING
C873 vdd.n6463 vss 7.48fF $ **FLOATING
C874 vdd.n6464 vss 7.48fF $ **FLOATING
C875 vdd.n6465 vss 7.48fF $ **FLOATING
C876 vdd.n6466 vss 7.48fF $ **FLOATING
C877 vdd.n6467 vss 7.48fF $ **FLOATING
C878 vdd.n6468 vss 7.48fF $ **FLOATING
C879 vdd.n6476 vss 5.17fF $ **FLOATING
C880 vdd.n6477 vss 5.17fF $ **FLOATING
C881 vdd.n6479 vss 7.28fF $ **FLOATING
C882 vdd.n6625 vss 5.17fF $ **FLOATING
C883 vdd.n6626 vss 5.17fF $ **FLOATING
C884 vdd.n6630 vss 7.24fF $ **FLOATING
C885 vdd.n6631 vss 7.48fF $ **FLOATING
C886 vdd.n6632 vss 7.48fF $ **FLOATING
C887 vdd.n6633 vss 7.48fF $ **FLOATING
C888 vdd.n6634 vss 7.48fF $ **FLOATING
C889 vdd.n6635 vss 7.48fF $ **FLOATING
C890 vdd.n6636 vss 7.48fF $ **FLOATING
C891 vdd.n6637 vss 7.48fF $ **FLOATING
C892 vdd.n6638 vss 7.48fF $ **FLOATING
C893 vdd.n6639 vss 7.48fF $ **FLOATING
C894 vdd.n6640 vss 7.48fF $ **FLOATING
C895 vdd.n6641 vss 7.48fF $ **FLOATING
C896 vdd.n6642 vss 7.48fF $ **FLOATING
C897 vdd.n6643 vss 7.48fF $ **FLOATING
C898 vdd.n6644 vss 7.48fF $ **FLOATING
C899 vdd.n6645 vss 7.48fF $ **FLOATING
C900 vdd.n6646 vss 7.48fF $ **FLOATING
C901 vdd.n6647 vss 7.48fF $ **FLOATING
C902 vdd.n6648 vss 7.48fF $ **FLOATING
C903 vdd.n6656 vss 5.17fF $ **FLOATING
C904 vdd.n6657 vss 5.17fF $ **FLOATING
C905 vdd.n6659 vss 7.28fF $ **FLOATING
C906 vdd.n6805 vss 5.17fF $ **FLOATING
C907 vdd.n6806 vss 5.17fF $ **FLOATING
C908 vdd.n6810 vss 7.24fF $ **FLOATING
C909 vdd.n6811 vss 7.48fF $ **FLOATING
C910 vdd.n6812 vss 7.48fF $ **FLOATING
C911 vdd.n6813 vss 7.48fF $ **FLOATING
C912 vdd.n6814 vss 7.48fF $ **FLOATING
C913 vdd.n6815 vss 7.48fF $ **FLOATING
C914 vdd.n6816 vss 7.48fF $ **FLOATING
C915 vdd.n6817 vss 7.48fF $ **FLOATING
C916 vdd.n6818 vss 7.48fF $ **FLOATING
C917 vdd.n6819 vss 7.48fF $ **FLOATING
C918 vdd.n6820 vss 7.48fF $ **FLOATING
C919 vdd.n6821 vss 7.48fF $ **FLOATING
C920 vdd.n6822 vss 7.48fF $ **FLOATING
C921 vdd.n6823 vss 7.48fF $ **FLOATING
C922 vdd.n6824 vss 7.48fF $ **FLOATING
C923 vdd.n6825 vss 7.48fF $ **FLOATING
C924 vdd.n6826 vss 7.48fF $ **FLOATING
C925 vdd.n6827 vss 7.48fF $ **FLOATING
C926 vdd.n6828 vss 7.48fF $ **FLOATING
C927 vdd.n6836 vss 5.17fF $ **FLOATING
C928 vdd.n6837 vss 5.17fF $ **FLOATING
C929 vdd.n6839 vss 7.28fF $ **FLOATING
C930 vdd.n6985 vss 5.17fF $ **FLOATING
C931 vdd.n6986 vss 5.17fF $ **FLOATING
C932 vdd.n6990 vss 7.24fF $ **FLOATING
C933 vdd.n6991 vss 7.48fF $ **FLOATING
C934 vdd.n6992 vss 7.48fF $ **FLOATING
C935 vdd.n6993 vss 7.48fF $ **FLOATING
C936 vdd.n6994 vss 7.48fF $ **FLOATING
C937 vdd.n6995 vss 7.48fF $ **FLOATING
C938 vdd.n6996 vss 7.48fF $ **FLOATING
C939 vdd.n6997 vss 7.48fF $ **FLOATING
C940 vdd.n6998 vss 7.48fF $ **FLOATING
C941 vdd.n6999 vss 7.48fF $ **FLOATING
C942 vdd.n7000 vss 7.48fF $ **FLOATING
C943 vdd.n7001 vss 7.48fF $ **FLOATING
C944 vdd.n7002 vss 7.48fF $ **FLOATING
C945 vdd.n7003 vss 7.48fF $ **FLOATING
C946 vdd.n7004 vss 7.48fF $ **FLOATING
C947 vdd.n7005 vss 7.48fF $ **FLOATING
C948 vdd.n7006 vss 7.48fF $ **FLOATING
C949 vdd.n7007 vss 7.48fF $ **FLOATING
C950 vdd.n7008 vss 7.48fF $ **FLOATING
C951 vdd.n7016 vss 5.17fF $ **FLOATING
C952 vdd.n7017 vss 5.17fF $ **FLOATING
C953 vdd.n7019 vss 7.28fF $ **FLOATING
C954 vdd.n7165 vss 5.17fF $ **FLOATING
C955 vdd.n7166 vss 5.17fF $ **FLOATING
C956 vdd.n7170 vss 7.24fF $ **FLOATING
C957 vdd.n7171 vss 7.48fF $ **FLOATING
C958 vdd.n7172 vss 7.48fF $ **FLOATING
C959 vdd.n7173 vss 7.48fF $ **FLOATING
C960 vdd.n7174 vss 7.48fF $ **FLOATING
C961 vdd.n7175 vss 7.48fF $ **FLOATING
C962 vdd.n7176 vss 7.48fF $ **FLOATING
C963 vdd.n7177 vss 7.48fF $ **FLOATING
C964 vdd.n7178 vss 7.48fF $ **FLOATING
C965 vdd.n7179 vss 7.48fF $ **FLOATING
C966 vdd.n7180 vss 7.48fF $ **FLOATING
C967 vdd.n7181 vss 7.48fF $ **FLOATING
C968 vdd.n7182 vss 7.48fF $ **FLOATING
C969 vdd.n7183 vss 7.48fF $ **FLOATING
C970 vdd.n7184 vss 7.48fF $ **FLOATING
C971 vdd.n7185 vss 7.48fF $ **FLOATING
C972 vdd.n7186 vss 7.48fF $ **FLOATING
C973 vdd.n7187 vss 7.48fF $ **FLOATING
C974 vdd.n7188 vss 7.48fF $ **FLOATING
C975 vdd.n7196 vss 5.17fF $ **FLOATING
C976 vdd.n7197 vss 5.17fF $ **FLOATING
C977 vdd.n7199 vss 7.28fF $ **FLOATING
C978 vdd.n7345 vss 5.17fF $ **FLOATING
C979 vdd.n7346 vss 5.17fF $ **FLOATING
C980 vdd.n7350 vss 7.24fF $ **FLOATING
C981 vdd.n7351 vss 7.48fF $ **FLOATING
C982 vdd.n7352 vss 7.48fF $ **FLOATING
C983 vdd.n7353 vss 7.48fF $ **FLOATING
C984 vdd.n7354 vss 7.48fF $ **FLOATING
C985 vdd.n7355 vss 7.48fF $ **FLOATING
C986 vdd.n7356 vss 7.48fF $ **FLOATING
C987 vdd.n7357 vss 7.48fF $ **FLOATING
C988 vdd.n7358 vss 7.48fF $ **FLOATING
C989 vdd.n7359 vss 7.48fF $ **FLOATING
C990 vdd.n7360 vss 7.48fF $ **FLOATING
C991 vdd.n7361 vss 7.48fF $ **FLOATING
C992 vdd.n7362 vss 7.48fF $ **FLOATING
C993 vdd.n7363 vss 7.48fF $ **FLOATING
C994 vdd.n7364 vss 7.48fF $ **FLOATING
C995 vdd.n7365 vss 7.48fF $ **FLOATING
C996 vdd.n7366 vss 7.48fF $ **FLOATING
C997 vdd.n7367 vss 7.48fF $ **FLOATING
C998 vdd.n7368 vss 7.48fF $ **FLOATING
C999 vdd.n7376 vss 5.17fF $ **FLOATING
C1000 vdd.n7377 vss 5.17fF $ **FLOATING
C1001 vdd.n7379 vss 7.28fF $ **FLOATING
C1002 vdd.n7525 vss 5.17fF $ **FLOATING
C1003 vdd.n7526 vss 5.17fF $ **FLOATING
C1004 vdd.n7530 vss 7.24fF $ **FLOATING
C1005 vdd.n7531 vss 7.48fF $ **FLOATING
C1006 vdd.n7532 vss 7.48fF $ **FLOATING
C1007 vdd.n7533 vss 7.48fF $ **FLOATING
C1008 vdd.n7534 vss 7.48fF $ **FLOATING
C1009 vdd.n7535 vss 7.48fF $ **FLOATING
C1010 vdd.n7536 vss 7.48fF $ **FLOATING
C1011 vdd.n7537 vss 7.48fF $ **FLOATING
C1012 vdd.n7538 vss 7.48fF $ **FLOATING
C1013 vdd.n7539 vss 7.48fF $ **FLOATING
C1014 vdd.n7540 vss 7.48fF $ **FLOATING
C1015 vdd.n7541 vss 7.48fF $ **FLOATING
C1016 vdd.n7542 vss 7.48fF $ **FLOATING
C1017 vdd.n7543 vss 7.48fF $ **FLOATING
C1018 vdd.n7544 vss 7.48fF $ **FLOATING
C1019 vdd.n7545 vss 7.48fF $ **FLOATING
C1020 vdd.n7546 vss 7.48fF $ **FLOATING
C1021 vdd.n7547 vss 7.48fF $ **FLOATING
C1022 vdd.n7548 vss 7.48fF $ **FLOATING
C1023 vdd.n7556 vss 5.17fF $ **FLOATING
C1024 vdd.n7557 vss 5.17fF $ **FLOATING
C1025 vdd.n7559 vss 7.28fF $ **FLOATING
C1026 vdd.n7705 vss 5.17fF $ **FLOATING
C1027 vdd.n7706 vss 5.17fF $ **FLOATING
C1028 vdd.n7710 vss 7.24fF $ **FLOATING
C1029 vdd.n7711 vss 7.48fF $ **FLOATING
C1030 vdd.n7712 vss 7.48fF $ **FLOATING
C1031 vdd.n7713 vss 7.48fF $ **FLOATING
C1032 vdd.n7714 vss 7.48fF $ **FLOATING
C1033 vdd.n7715 vss 7.48fF $ **FLOATING
C1034 vdd.n7716 vss 7.48fF $ **FLOATING
C1035 vdd.n7717 vss 7.48fF $ **FLOATING
C1036 vdd.n7718 vss 7.48fF $ **FLOATING
C1037 vdd.n7719 vss 7.48fF $ **FLOATING
C1038 vdd.n7720 vss 7.48fF $ **FLOATING
C1039 vdd.n7721 vss 7.48fF $ **FLOATING
C1040 vdd.n7722 vss 7.48fF $ **FLOATING
C1041 vdd.n7723 vss 7.48fF $ **FLOATING
C1042 vdd.n7724 vss 7.48fF $ **FLOATING
C1043 vdd.n7725 vss 7.48fF $ **FLOATING
C1044 vdd.n7726 vss 7.48fF $ **FLOATING
C1045 vdd.n7727 vss 7.48fF $ **FLOATING
C1046 vdd.n7728 vss 7.48fF $ **FLOATING
C1047 vdd.n7736 vss 5.17fF $ **FLOATING
C1048 vdd.n7737 vss 5.17fF $ **FLOATING
C1049 vdd.n7739 vss 7.28fF $ **FLOATING
C1050 vdd.n7885 vss 5.17fF $ **FLOATING
C1051 vdd.n7886 vss 5.17fF $ **FLOATING
C1052 vdd.n7890 vss 7.24fF $ **FLOATING
C1053 vdd.n7891 vss 7.48fF $ **FLOATING
C1054 vdd.n7892 vss 7.48fF $ **FLOATING
C1055 vdd.n7893 vss 7.48fF $ **FLOATING
C1056 vdd.n7894 vss 7.48fF $ **FLOATING
C1057 vdd.n7895 vss 7.48fF $ **FLOATING
C1058 vdd.n7896 vss 7.48fF $ **FLOATING
C1059 vdd.n7897 vss 7.48fF $ **FLOATING
C1060 vdd.n7898 vss 7.48fF $ **FLOATING
C1061 vdd.n7899 vss 7.48fF $ **FLOATING
C1062 vdd.n7900 vss 7.48fF $ **FLOATING
C1063 vdd.n7901 vss 7.48fF $ **FLOATING
C1064 vdd.n7902 vss 7.48fF $ **FLOATING
C1065 vdd.n7903 vss 7.48fF $ **FLOATING
C1066 vdd.n7904 vss 7.48fF $ **FLOATING
C1067 vdd.n7905 vss 7.48fF $ **FLOATING
C1068 vdd.n7906 vss 7.48fF $ **FLOATING
C1069 vdd.n7907 vss 7.48fF $ **FLOATING
C1070 vdd.n7908 vss 7.48fF $ **FLOATING
C1071 vdd.n7916 vss 5.17fF $ **FLOATING
C1072 vdd.n7917 vss 5.17fF $ **FLOATING
C1073 vdd.n7919 vss 7.28fF $ **FLOATING
C1074 vdd.n8065 vss 5.17fF $ **FLOATING
C1075 vdd.n8066 vss 5.17fF $ **FLOATING
C1076 vdd.n8070 vss 7.24fF $ **FLOATING
C1077 vdd.n8071 vss 7.48fF $ **FLOATING
C1078 vdd.n8072 vss 7.48fF $ **FLOATING
C1079 vdd.n8073 vss 7.48fF $ **FLOATING
C1080 vdd.n8074 vss 7.48fF $ **FLOATING
C1081 vdd.n8075 vss 7.48fF $ **FLOATING
C1082 vdd.n8076 vss 7.48fF $ **FLOATING
C1083 vdd.n8077 vss 7.48fF $ **FLOATING
C1084 vdd.n8078 vss 7.48fF $ **FLOATING
C1085 vdd.n8079 vss 7.48fF $ **FLOATING
C1086 vdd.n8080 vss 7.48fF $ **FLOATING
C1087 vdd.n8081 vss 7.48fF $ **FLOATING
C1088 vdd.n8082 vss 7.48fF $ **FLOATING
C1089 vdd.n8083 vss 7.48fF $ **FLOATING
C1090 vdd.n8084 vss 7.48fF $ **FLOATING
C1091 vdd.n8085 vss 7.48fF $ **FLOATING
C1092 vdd.n8086 vss 7.48fF $ **FLOATING
C1093 vdd.n8087 vss 7.48fF $ **FLOATING
C1094 vdd.n8088 vss 7.48fF $ **FLOATING
C1095 vdd.n8096 vss 5.17fF $ **FLOATING
C1096 vdd.n8097 vss 5.17fF $ **FLOATING
C1097 vdd.n8099 vss 7.28fF $ **FLOATING
C1098 vdd.n8245 vss 5.17fF $ **FLOATING
C1099 vdd.n8246 vss 5.17fF $ **FLOATING
C1100 vdd.n8250 vss 7.24fF $ **FLOATING
C1101 vdd.n8251 vss 7.48fF $ **FLOATING
C1102 vdd.n8252 vss 7.48fF $ **FLOATING
C1103 vdd.n8253 vss 7.48fF $ **FLOATING
C1104 vdd.n8254 vss 7.48fF $ **FLOATING
C1105 vdd.n8255 vss 7.48fF $ **FLOATING
C1106 vdd.n8256 vss 7.48fF $ **FLOATING
C1107 vdd.n8257 vss 7.48fF $ **FLOATING
C1108 vdd.n8258 vss 7.48fF $ **FLOATING
C1109 vdd.n8259 vss 7.48fF $ **FLOATING
C1110 vdd.n8260 vss 7.48fF $ **FLOATING
C1111 vdd.n8261 vss 7.48fF $ **FLOATING
C1112 vdd.n8262 vss 7.48fF $ **FLOATING
C1113 vdd.n8263 vss 7.48fF $ **FLOATING
C1114 vdd.n8264 vss 7.48fF $ **FLOATING
C1115 vdd.n8265 vss 7.48fF $ **FLOATING
C1116 vdd.n8266 vss 7.48fF $ **FLOATING
C1117 vdd.n8267 vss 7.48fF $ **FLOATING
C1118 vdd.n8268 vss 7.48fF $ **FLOATING
C1119 vdd.n8276 vss 5.17fF $ **FLOATING
C1120 vdd.n8277 vss 5.17fF $ **FLOATING
C1121 vdd.n8279 vss 7.28fF $ **FLOATING
C1122 vdd.n8425 vss 5.17fF $ **FLOATING
C1123 vdd.n8426 vss 5.17fF $ **FLOATING
C1124 vdd.n8430 vss 7.24fF $ **FLOATING
C1125 vdd.n8431 vss 7.48fF $ **FLOATING
C1126 vdd.n8432 vss 7.48fF $ **FLOATING
C1127 vdd.n8433 vss 7.48fF $ **FLOATING
C1128 vdd.n8434 vss 7.48fF $ **FLOATING
C1129 vdd.n8435 vss 7.48fF $ **FLOATING
C1130 vdd.n8436 vss 7.48fF $ **FLOATING
C1131 vdd.n8437 vss 7.48fF $ **FLOATING
C1132 vdd.n8438 vss 7.48fF $ **FLOATING
C1133 vdd.n8439 vss 7.48fF $ **FLOATING
C1134 vdd.n8440 vss 7.48fF $ **FLOATING
C1135 vdd.n8441 vss 7.48fF $ **FLOATING
C1136 vdd.n8442 vss 7.48fF $ **FLOATING
C1137 vdd.n8443 vss 7.48fF $ **FLOATING
C1138 vdd.n8444 vss 7.48fF $ **FLOATING
C1139 vdd.n8445 vss 7.48fF $ **FLOATING
C1140 vdd.n8446 vss 7.48fF $ **FLOATING
C1141 vdd.n8447 vss 7.48fF $ **FLOATING
C1142 vdd.n8448 vss 7.48fF $ **FLOATING
C1143 vdd.n8456 vss 5.17fF $ **FLOATING
C1144 vdd.n8457 vss 5.17fF $ **FLOATING
C1145 vdd.n8459 vss 7.28fF $ **FLOATING
C1146 vdd.n8605 vss 5.17fF $ **FLOATING
C1147 vdd.n8606 vss 5.17fF $ **FLOATING
C1148 vdd.n8610 vss 7.24fF $ **FLOATING
C1149 vdd.n8611 vss 7.48fF $ **FLOATING
C1150 vdd.n8612 vss 7.48fF $ **FLOATING
C1151 vdd.n8613 vss 7.48fF $ **FLOATING
C1152 vdd.n8614 vss 7.48fF $ **FLOATING
C1153 vdd.n8615 vss 7.48fF $ **FLOATING
C1154 vdd.n8616 vss 7.48fF $ **FLOATING
C1155 vdd.n8617 vss 7.48fF $ **FLOATING
C1156 vdd.n8618 vss 7.48fF $ **FLOATING
C1157 vdd.n8619 vss 7.48fF $ **FLOATING
C1158 vdd.n8620 vss 7.48fF $ **FLOATING
C1159 vdd.n8621 vss 7.48fF $ **FLOATING
C1160 vdd.n8622 vss 7.48fF $ **FLOATING
C1161 vdd.n8623 vss 7.48fF $ **FLOATING
C1162 vdd.n8624 vss 7.48fF $ **FLOATING
C1163 vdd.n8625 vss 7.48fF $ **FLOATING
C1164 vdd.n8626 vss 7.48fF $ **FLOATING
C1165 vdd.n8627 vss 7.48fF $ **FLOATING
C1166 vdd.n8628 vss 7.48fF $ **FLOATING
C1167 vdd.n8636 vss 5.17fF $ **FLOATING
C1168 vdd.n8637 vss 5.17fF $ **FLOATING
C1169 vdd.n8639 vss 7.28fF $ **FLOATING
C1170 vdd.n8785 vss 5.17fF $ **FLOATING
C1171 vdd.n8786 vss 5.17fF $ **FLOATING
C1172 vdd.n8790 vss 7.24fF $ **FLOATING
C1173 vdd.n8791 vss 7.48fF $ **FLOATING
C1174 vdd.n8792 vss 7.48fF $ **FLOATING
C1175 vdd.n8793 vss 7.48fF $ **FLOATING
C1176 vdd.n8794 vss 7.48fF $ **FLOATING
C1177 vdd.n8795 vss 7.48fF $ **FLOATING
C1178 vdd.n8796 vss 7.48fF $ **FLOATING
C1179 vdd.n8797 vss 7.48fF $ **FLOATING
C1180 vdd.n8798 vss 7.48fF $ **FLOATING
C1181 vdd.n8799 vss 7.48fF $ **FLOATING
C1182 vdd.n8800 vss 7.48fF $ **FLOATING
C1183 vdd.n8801 vss 7.48fF $ **FLOATING
C1184 vdd.n8802 vss 7.48fF $ **FLOATING
C1185 vdd.n8803 vss 7.48fF $ **FLOATING
C1186 vdd.n8804 vss 7.48fF $ **FLOATING
C1187 vdd.n8805 vss 7.48fF $ **FLOATING
C1188 vdd.n8806 vss 7.48fF $ **FLOATING
C1189 vdd.n8807 vss 7.48fF $ **FLOATING
C1190 vdd.n8808 vss 7.48fF $ **FLOATING
C1191 vdd.n8816 vss 5.17fF $ **FLOATING
C1192 vdd.n8817 vss 5.17fF $ **FLOATING
C1193 vdd.n8819 vss 7.28fF $ **FLOATING
C1194 vdd.n8965 vss 5.17fF $ **FLOATING
C1195 vdd.n8966 vss 5.17fF $ **FLOATING
C1196 vdd.n8970 vss 7.24fF $ **FLOATING
C1197 vdd.n8971 vss 7.48fF $ **FLOATING
C1198 vdd.n8972 vss 7.48fF $ **FLOATING
C1199 vdd.n8973 vss 7.48fF $ **FLOATING
C1200 vdd.n8974 vss 7.48fF $ **FLOATING
C1201 vdd.n8975 vss 7.48fF $ **FLOATING
C1202 vdd.n8976 vss 7.48fF $ **FLOATING
C1203 vdd.n8977 vss 7.48fF $ **FLOATING
C1204 vdd.n8978 vss 7.48fF $ **FLOATING
C1205 vdd.n8979 vss 7.48fF $ **FLOATING
C1206 vdd.n8980 vss 7.48fF $ **FLOATING
C1207 vdd.n8981 vss 7.48fF $ **FLOATING
C1208 vdd.n8982 vss 7.48fF $ **FLOATING
C1209 vdd.n8983 vss 7.48fF $ **FLOATING
C1210 vdd.n8984 vss 7.48fF $ **FLOATING
C1211 vdd.n8985 vss 7.48fF $ **FLOATING
C1212 vdd.n8986 vss 7.48fF $ **FLOATING
C1213 vdd.n8987 vss 7.48fF $ **FLOATING
C1214 vdd.n8988 vss 7.48fF $ **FLOATING
C1215 vdd.n8996 vss 5.17fF $ **FLOATING
C1216 vdd.n8997 vss 5.17fF $ **FLOATING
C1217 vdd.n8999 vss 7.28fF $ **FLOATING
C1218 vdd.n9145 vss 5.17fF $ **FLOATING
C1219 vdd.n9146 vss 5.17fF $ **FLOATING
C1220 vdd.n9150 vss 7.24fF $ **FLOATING
C1221 vdd.n9151 vss 7.48fF $ **FLOATING
C1222 vdd.n9152 vss 7.48fF $ **FLOATING
C1223 vdd.n9153 vss 7.48fF $ **FLOATING
C1224 vdd.n9154 vss 7.48fF $ **FLOATING
C1225 vdd.n9155 vss 7.48fF $ **FLOATING
C1226 vdd.n9156 vss 7.48fF $ **FLOATING
C1227 vdd.n9157 vss 7.48fF $ **FLOATING
C1228 vdd.n9158 vss 7.48fF $ **FLOATING
C1229 vdd.n9159 vss 7.48fF $ **FLOATING
C1230 vdd.n9160 vss 7.48fF $ **FLOATING
C1231 vdd.n9161 vss 7.48fF $ **FLOATING
C1232 vdd.n9162 vss 7.48fF $ **FLOATING
C1233 vdd.n9163 vss 7.48fF $ **FLOATING
C1234 vdd.n9164 vss 7.48fF $ **FLOATING
C1235 vdd.n9165 vss 7.48fF $ **FLOATING
C1236 vdd.n9166 vss 7.48fF $ **FLOATING
C1237 vdd.n9167 vss 7.48fF $ **FLOATING
C1238 vdd.n9168 vss 7.48fF $ **FLOATING
C1239 vdd.n9176 vss 5.17fF $ **FLOATING
C1240 vdd.n9177 vss 5.17fF $ **FLOATING
C1241 vdd.n9179 vss 7.28fF $ **FLOATING
C1242 vdd.n9325 vss 5.17fF $ **FLOATING
C1243 vdd.n9326 vss 5.17fF $ **FLOATING
C1244 vdd.n9330 vss 7.24fF $ **FLOATING
C1245 vdd.n9331 vss 7.48fF $ **FLOATING
C1246 vdd.n9332 vss 7.48fF $ **FLOATING
C1247 vdd.n9333 vss 7.48fF $ **FLOATING
C1248 vdd.n9334 vss 7.48fF $ **FLOATING
C1249 vdd.n9335 vss 7.48fF $ **FLOATING
C1250 vdd.n9336 vss 7.48fF $ **FLOATING
C1251 vdd.n9337 vss 7.48fF $ **FLOATING
C1252 vdd.n9338 vss 7.48fF $ **FLOATING
C1253 vdd.n9339 vss 7.48fF $ **FLOATING
C1254 vdd.n9340 vss 7.48fF $ **FLOATING
C1255 vdd.n9341 vss 7.48fF $ **FLOATING
C1256 vdd.n9342 vss 7.48fF $ **FLOATING
C1257 vdd.n9343 vss 7.48fF $ **FLOATING
C1258 vdd.n9344 vss 7.48fF $ **FLOATING
C1259 vdd.n9345 vss 7.48fF $ **FLOATING
C1260 vdd.n9346 vss 7.48fF $ **FLOATING
C1261 vdd.n9347 vss 7.48fF $ **FLOATING
C1262 vdd.n9348 vss 7.48fF $ **FLOATING
C1263 vdd.n9356 vss 5.17fF $ **FLOATING
C1264 vdd.n9357 vss 5.17fF $ **FLOATING
C1265 vdd.n9359 vss 7.28fF $ **FLOATING
C1266 vdd.n9505 vss 5.17fF $ **FLOATING
C1267 vdd.n9506 vss 5.17fF $ **FLOATING
C1268 vdd.n9510 vss 7.24fF $ **FLOATING
C1269 vdd.n9511 vss 7.48fF $ **FLOATING
C1270 vdd.n9512 vss 7.48fF $ **FLOATING
C1271 vdd.n9513 vss 7.48fF $ **FLOATING
C1272 vdd.n9514 vss 7.48fF $ **FLOATING
C1273 vdd.n9515 vss 7.48fF $ **FLOATING
C1274 vdd.n9516 vss 7.48fF $ **FLOATING
C1275 vdd.n9517 vss 7.48fF $ **FLOATING
C1276 vdd.n9518 vss 7.48fF $ **FLOATING
C1277 vdd.n9519 vss 7.48fF $ **FLOATING
C1278 vdd.n9520 vss 7.48fF $ **FLOATING
C1279 vdd.n9521 vss 7.48fF $ **FLOATING
C1280 vdd.n9522 vss 7.48fF $ **FLOATING
C1281 vdd.n9523 vss 7.48fF $ **FLOATING
C1282 vdd.n9524 vss 7.48fF $ **FLOATING
C1283 vdd.n9525 vss 7.48fF $ **FLOATING
C1284 vdd.n9526 vss 7.48fF $ **FLOATING
C1285 vdd.n9527 vss 7.48fF $ **FLOATING
C1286 vdd.n9528 vss 7.48fF $ **FLOATING
C1287 vdd.n9536 vss 5.17fF $ **FLOATING
C1288 vdd.n9537 vss 5.17fF $ **FLOATING
C1289 vdd.n9539 vss 7.28fF $ **FLOATING
C1290 vdd.n9685 vss 5.17fF $ **FLOATING
C1291 vdd.n9686 vss 5.17fF $ **FLOATING
C1292 vdd.n9690 vss 7.24fF $ **FLOATING
C1293 vdd.n9691 vss 7.48fF $ **FLOATING
C1294 vdd.n9692 vss 7.48fF $ **FLOATING
C1295 vdd.n9693 vss 7.48fF $ **FLOATING
C1296 vdd.n9694 vss 7.48fF $ **FLOATING
C1297 vdd.n9695 vss 7.48fF $ **FLOATING
C1298 vdd.n9696 vss 7.48fF $ **FLOATING
C1299 vdd.n9697 vss 7.48fF $ **FLOATING
C1300 vdd.n9698 vss 7.48fF $ **FLOATING
C1301 vdd.n9699 vss 7.48fF $ **FLOATING
C1302 vdd.n9700 vss 7.48fF $ **FLOATING
C1303 vdd.n9701 vss 7.48fF $ **FLOATING
C1304 vdd.n9702 vss 7.48fF $ **FLOATING
C1305 vdd.n9703 vss 7.48fF $ **FLOATING
C1306 vdd.n9704 vss 7.48fF $ **FLOATING
C1307 vdd.n9705 vss 7.48fF $ **FLOATING
C1308 vdd.n9706 vss 7.48fF $ **FLOATING
C1309 vdd.n9707 vss 7.48fF $ **FLOATING
C1310 vdd.n9708 vss 7.48fF $ **FLOATING
C1311 vdd.n9716 vss 5.17fF $ **FLOATING
C1312 vdd.n9717 vss 5.17fF $ **FLOATING
C1313 vdd.n9719 vss 7.28fF $ **FLOATING
C1314 vdd.n9865 vss 5.17fF $ **FLOATING
C1315 vdd.n9866 vss 5.17fF $ **FLOATING
C1316 vdd.n9870 vss 7.24fF $ **FLOATING
C1317 vdd.n9871 vss 7.48fF $ **FLOATING
C1318 vdd.n9872 vss 7.48fF $ **FLOATING
C1319 vdd.n9873 vss 7.48fF $ **FLOATING
C1320 vdd.n9874 vss 7.48fF $ **FLOATING
C1321 vdd.n9875 vss 7.48fF $ **FLOATING
C1322 vdd.n9876 vss 7.48fF $ **FLOATING
C1323 vdd.n9877 vss 7.48fF $ **FLOATING
C1324 vdd.n9878 vss 7.48fF $ **FLOATING
C1325 vdd.n9879 vss 7.48fF $ **FLOATING
C1326 vdd.n9880 vss 7.48fF $ **FLOATING
C1327 vdd.n9881 vss 7.48fF $ **FLOATING
C1328 vdd.n9882 vss 7.48fF $ **FLOATING
C1329 vdd.n9883 vss 7.48fF $ **FLOATING
C1330 vdd.n9884 vss 7.48fF $ **FLOATING
C1331 vdd.n9885 vss 7.48fF $ **FLOATING
C1332 vdd.n9886 vss 7.48fF $ **FLOATING
C1333 vdd.n9887 vss 7.48fF $ **FLOATING
C1334 vdd.n9888 vss 7.48fF $ **FLOATING
C1335 vdd.n9896 vss 5.17fF $ **FLOATING
C1336 vdd.n9897 vss 5.17fF $ **FLOATING
C1337 vdd.n9899 vss 7.28fF $ **FLOATING
C1338 vdd.n10045 vss 5.17fF $ **FLOATING
C1339 vdd.n10046 vss 5.17fF $ **FLOATING
C1340 vdd.n10050 vss 7.24fF $ **FLOATING
C1341 vdd.n10051 vss 7.48fF $ **FLOATING
C1342 vdd.n10052 vss 7.48fF $ **FLOATING
C1343 vdd.n10053 vss 7.48fF $ **FLOATING
C1344 vdd.n10054 vss 7.48fF $ **FLOATING
C1345 vdd.n10055 vss 7.48fF $ **FLOATING
C1346 vdd.n10056 vss 7.48fF $ **FLOATING
C1347 vdd.n10057 vss 7.48fF $ **FLOATING
C1348 vdd.n10058 vss 7.48fF $ **FLOATING
C1349 vdd.n10059 vss 7.48fF $ **FLOATING
C1350 vdd.n10060 vss 7.48fF $ **FLOATING
C1351 vdd.n10061 vss 7.48fF $ **FLOATING
C1352 vdd.n10062 vss 7.48fF $ **FLOATING
C1353 vdd.n10063 vss 7.48fF $ **FLOATING
C1354 vdd.n10064 vss 7.48fF $ **FLOATING
C1355 vdd.n10065 vss 7.48fF $ **FLOATING
C1356 vdd.n10066 vss 7.48fF $ **FLOATING
C1357 vdd.n10067 vss 7.48fF $ **FLOATING
C1358 vdd.n10068 vss 7.48fF $ **FLOATING
C1359 vdd.n10076 vss 5.17fF $ **FLOATING
C1360 vdd.n10077 vss 5.17fF $ **FLOATING
C1361 vdd.n10079 vss 7.28fF $ **FLOATING
C1362 vdd.n10225 vss 5.17fF $ **FLOATING
C1363 vdd.n10226 vss 5.17fF $ **FLOATING
C1364 vdd.n10230 vss 7.24fF $ **FLOATING
C1365 vdd.n10231 vss 7.48fF $ **FLOATING
C1366 vdd.n10232 vss 7.48fF $ **FLOATING
C1367 vdd.n10233 vss 7.48fF $ **FLOATING
C1368 vdd.n10234 vss 7.48fF $ **FLOATING
C1369 vdd.n10235 vss 7.48fF $ **FLOATING
C1370 vdd.n10236 vss 7.48fF $ **FLOATING
C1371 vdd.n10237 vss 7.48fF $ **FLOATING
C1372 vdd.n10238 vss 7.48fF $ **FLOATING
C1373 vdd.n10239 vss 7.48fF $ **FLOATING
C1374 vdd.n10240 vss 7.48fF $ **FLOATING
C1375 vdd.n10241 vss 7.48fF $ **FLOATING
C1376 vdd.n10242 vss 7.48fF $ **FLOATING
C1377 vdd.n10243 vss 7.48fF $ **FLOATING
C1378 vdd.n10244 vss 7.48fF $ **FLOATING
C1379 vdd.n10245 vss 7.48fF $ **FLOATING
C1380 vdd.n10246 vss 7.48fF $ **FLOATING
C1381 vdd.n10247 vss 7.48fF $ **FLOATING
C1382 vdd.n10248 vss 7.48fF $ **FLOATING
C1383 vdd.n10256 vss 5.17fF $ **FLOATING
C1384 vdd.n10257 vss 5.17fF $ **FLOATING
C1385 vdd.n10259 vss 7.28fF $ **FLOATING
C1386 vdd.n10405 vss 5.17fF $ **FLOATING
C1387 vdd.n10406 vss 5.17fF $ **FLOATING
C1388 vdd.n10410 vss 7.24fF $ **FLOATING
C1389 vdd.n10411 vss 7.48fF $ **FLOATING
C1390 vdd.n10412 vss 7.48fF $ **FLOATING
C1391 vdd.n10413 vss 7.48fF $ **FLOATING
C1392 vdd.n10414 vss 7.48fF $ **FLOATING
C1393 vdd.n10415 vss 7.48fF $ **FLOATING
C1394 vdd.n10416 vss 7.48fF $ **FLOATING
C1395 vdd.n10417 vss 7.48fF $ **FLOATING
C1396 vdd.n10418 vss 7.48fF $ **FLOATING
C1397 vdd.n10419 vss 7.48fF $ **FLOATING
C1398 vdd.n10420 vss 7.48fF $ **FLOATING
C1399 vdd.n10421 vss 7.48fF $ **FLOATING
C1400 vdd.n10422 vss 7.48fF $ **FLOATING
C1401 vdd.n10423 vss 7.48fF $ **FLOATING
C1402 vdd.n10424 vss 7.48fF $ **FLOATING
C1403 vdd.n10425 vss 7.48fF $ **FLOATING
C1404 vdd.n10426 vss 7.48fF $ **FLOATING
C1405 vdd.n10427 vss 7.48fF $ **FLOATING
C1406 vdd.n10428 vss 7.48fF $ **FLOATING
C1407 vdd.n10436 vss 5.17fF $ **FLOATING
C1408 vdd.n10437 vss 5.17fF $ **FLOATING
C1409 vdd.n10439 vss 7.28fF $ **FLOATING
C1410 vdd.n10585 vss 5.17fF $ **FLOATING
C1411 vdd.n10586 vss 5.17fF $ **FLOATING
C1412 vdd.n10590 vss 7.24fF $ **FLOATING
C1413 vdd.n10591 vss 7.48fF $ **FLOATING
C1414 vdd.n10592 vss 7.48fF $ **FLOATING
C1415 vdd.n10593 vss 7.48fF $ **FLOATING
C1416 vdd.n10594 vss 7.48fF $ **FLOATING
C1417 vdd.n10595 vss 7.48fF $ **FLOATING
C1418 vdd.n10596 vss 7.48fF $ **FLOATING
C1419 vdd.n10597 vss 7.48fF $ **FLOATING
C1420 vdd.n10598 vss 7.48fF $ **FLOATING
C1421 vdd.n10599 vss 7.48fF $ **FLOATING
C1422 vdd.n10600 vss 7.48fF $ **FLOATING
C1423 vdd.n10601 vss 7.48fF $ **FLOATING
C1424 vdd.n10602 vss 7.48fF $ **FLOATING
C1425 vdd.n10603 vss 7.48fF $ **FLOATING
C1426 vdd.n10604 vss 7.48fF $ **FLOATING
C1427 vdd.n10605 vss 7.48fF $ **FLOATING
C1428 vdd.n10606 vss 7.48fF $ **FLOATING
C1429 vdd.n10607 vss 7.48fF $ **FLOATING
C1430 vdd.n10608 vss 7.48fF $ **FLOATING
C1431 vdd.n10616 vss 5.17fF $ **FLOATING
C1432 vdd.n10617 vss 5.17fF $ **FLOATING
C1433 vdd.n10619 vss 7.28fF $ **FLOATING
C1434 vdd.n10765 vss 5.17fF $ **FLOATING
C1435 vdd.n10766 vss 5.17fF $ **FLOATING
C1436 vdd.n10770 vss 7.24fF $ **FLOATING
C1437 vdd.n10771 vss 7.48fF $ **FLOATING
C1438 vdd.n10772 vss 7.48fF $ **FLOATING
C1439 vdd.n10773 vss 7.48fF $ **FLOATING
C1440 vdd.n10774 vss 7.48fF $ **FLOATING
C1441 vdd.n10775 vss 7.48fF $ **FLOATING
C1442 vdd.n10776 vss 7.48fF $ **FLOATING
C1443 vdd.n10777 vss 7.48fF $ **FLOATING
C1444 vdd.n10778 vss 7.48fF $ **FLOATING
C1445 vdd.n10779 vss 7.48fF $ **FLOATING
C1446 vdd.n10780 vss 7.48fF $ **FLOATING
C1447 vdd.n10781 vss 7.48fF $ **FLOATING
C1448 vdd.n10782 vss 7.48fF $ **FLOATING
C1449 vdd.n10783 vss 7.48fF $ **FLOATING
C1450 vdd.n10784 vss 7.48fF $ **FLOATING
C1451 vdd.n10785 vss 7.48fF $ **FLOATING
C1452 vdd.n10786 vss 7.48fF $ **FLOATING
C1453 vdd.n10787 vss 7.48fF $ **FLOATING
C1454 vdd.n10788 vss 7.48fF $ **FLOATING
C1455 vdd.n10796 vss 5.17fF $ **FLOATING
C1456 vdd.n10797 vss 5.17fF $ **FLOATING
C1457 vdd.n10799 vss 7.28fF $ **FLOATING
C1458 vdd.n10945 vss 5.17fF $ **FLOATING
C1459 vdd.n10946 vss 5.17fF $ **FLOATING
C1460 vdd.n10950 vss 7.24fF $ **FLOATING
C1461 vdd.n10951 vss 7.48fF $ **FLOATING
C1462 vdd.n10952 vss 7.48fF $ **FLOATING
C1463 vdd.n10953 vss 7.48fF $ **FLOATING
C1464 vdd.n10954 vss 7.48fF $ **FLOATING
C1465 vdd.n10955 vss 7.48fF $ **FLOATING
C1466 vdd.n10956 vss 7.48fF $ **FLOATING
C1467 vdd.n10957 vss 7.48fF $ **FLOATING
C1468 vdd.n10958 vss 7.48fF $ **FLOATING
C1469 vdd.n10959 vss 7.48fF $ **FLOATING
C1470 vdd.n10960 vss 7.48fF $ **FLOATING
C1471 vdd.n10961 vss 7.48fF $ **FLOATING
C1472 vdd.n10962 vss 7.48fF $ **FLOATING
C1473 vdd.n10963 vss 7.48fF $ **FLOATING
C1474 vdd.n10964 vss 7.48fF $ **FLOATING
C1475 vdd.n10965 vss 7.48fF $ **FLOATING
C1476 vdd.n10966 vss 7.48fF $ **FLOATING
C1477 vdd.n10967 vss 7.48fF $ **FLOATING
C1478 vdd.n10968 vss 7.48fF $ **FLOATING
C1479 vdd.n10976 vss 5.17fF $ **FLOATING
C1480 vdd.n10977 vss 5.17fF $ **FLOATING
C1481 vdd.n10979 vss 7.28fF $ **FLOATING
C1482 vdd.n11125 vss 5.17fF $ **FLOATING
C1483 vdd.n11126 vss 5.17fF $ **FLOATING
C1484 vdd.n11130 vss 7.24fF $ **FLOATING
C1485 vdd.n11131 vss 7.48fF $ **FLOATING
C1486 vdd.n11132 vss 7.48fF $ **FLOATING
C1487 vdd.n11133 vss 7.48fF $ **FLOATING
C1488 vdd.n11134 vss 7.48fF $ **FLOATING
C1489 vdd.n11135 vss 7.48fF $ **FLOATING
C1490 vdd.n11136 vss 7.48fF $ **FLOATING
C1491 vdd.n11137 vss 7.48fF $ **FLOATING
C1492 vdd.n11138 vss 7.48fF $ **FLOATING
C1493 vdd.n11139 vss 7.48fF $ **FLOATING
C1494 vdd.n11140 vss 7.48fF $ **FLOATING
C1495 vdd.n11141 vss 7.48fF $ **FLOATING
C1496 vdd.n11142 vss 7.48fF $ **FLOATING
C1497 vdd.n11143 vss 7.48fF $ **FLOATING
C1498 vdd.n11144 vss 7.48fF $ **FLOATING
C1499 vdd.n11145 vss 7.48fF $ **FLOATING
C1500 vdd.n11146 vss 7.48fF $ **FLOATING
C1501 vdd.n11147 vss 7.48fF $ **FLOATING
C1502 vdd.n11148 vss 7.48fF $ **FLOATING
C1503 vdd.n11156 vss 5.17fF $ **FLOATING
C1504 vdd.n11157 vss 5.17fF $ **FLOATING
C1505 vdd.n11159 vss 7.28fF $ **FLOATING
C1506 vdd.n11305 vss 5.17fF $ **FLOATING
C1507 vdd.n11306 vss 5.17fF $ **FLOATING
C1508 vdd.n11310 vss 7.24fF $ **FLOATING
C1509 vdd.n11311 vss 7.48fF $ **FLOATING
C1510 vdd.n11312 vss 7.48fF $ **FLOATING
C1511 vdd.n11313 vss 7.48fF $ **FLOATING
C1512 vdd.n11314 vss 7.48fF $ **FLOATING
C1513 vdd.n11315 vss 7.48fF $ **FLOATING
C1514 vdd.n11316 vss 7.48fF $ **FLOATING
C1515 vdd.n11317 vss 7.48fF $ **FLOATING
C1516 vdd.n11318 vss 7.48fF $ **FLOATING
C1517 vdd.n11319 vss 7.48fF $ **FLOATING
C1518 vdd.n11320 vss 7.48fF $ **FLOATING
C1519 vdd.n11321 vss 7.48fF $ **FLOATING
C1520 vdd.n11322 vss 7.48fF $ **FLOATING
C1521 vdd.n11323 vss 7.48fF $ **FLOATING
C1522 vdd.n11324 vss 7.48fF $ **FLOATING
C1523 vdd.n11325 vss 7.48fF $ **FLOATING
C1524 vdd.n11326 vss 7.48fF $ **FLOATING
C1525 vdd.n11327 vss 7.48fF $ **FLOATING
C1526 vdd.n11328 vss 7.48fF $ **FLOATING
C1527 vdd.n11336 vss 5.17fF $ **FLOATING
C1528 vdd.n11337 vss 5.17fF $ **FLOATING
C1529 vdd.n11339 vss 7.28fF $ **FLOATING
C1530 vdd.n11358 vss 5.36fF $ **FLOATING
C1531 vdd.n11359 vss 4.13fF $ **FLOATING
C1532 vdd.n11362 vss 4.31fF $ **FLOATING
C1533 vdd.n11365 vss 4.31fF $ **FLOATING
C1534 vdd.n11368 vss 4.31fF $ **FLOATING
C1535 vdd.n11371 vss 4.31fF $ **FLOATING
C1536 vdd.n11374 vss 4.31fF $ **FLOATING
C1537 vdd.n11377 vss 4.31fF $ **FLOATING
C1538 vdd.n11380 vss 4.31fF $ **FLOATING
C1539 vdd.n11383 vss 4.31fF $ **FLOATING
C1540 vdd.n11386 vss 4.31fF $ **FLOATING
C1541 vdd.n11387 vss 4.31fF $ **FLOATING
C1542 vdd.n11390 vss 4.31fF $ **FLOATING
C1543 vdd.n11393 vss 4.31fF $ **FLOATING
C1544 vdd.n11396 vss 4.31fF $ **FLOATING
C1545 vdd.n11399 vss 4.31fF $ **FLOATING
C1546 vdd.n11402 vss 4.31fF $ **FLOATING
C1547 vdd.n11405 vss 4.31fF $ **FLOATING
C1548 vdd.n11408 vss 4.31fF $ **FLOATING
C1549 vdd.n11411 vss 4.31fF $ **FLOATING
C1550 vdd.n11414 vss 5.36fF $ **FLOATING
C1551 vdd.n11415 vss 4.78fF $ **FLOATING
C1552 vdd.n11416 vss 136.24fF $ **FLOATING
C1553 vdd.n11417 vss 76.29fF $ **FLOATING
C1554 vdd.n11418 vss 76.29fF $ **FLOATING
C1555 vdd.n11419 vss 76.29fF $ **FLOATING
C1556 vdd.n11420 vss 76.29fF $ **FLOATING
C1557 vdd.n11421 vss 76.29fF $ **FLOATING
C1558 vdd.n11422 vss 76.29fF $ **FLOATING
C1559 vdd.n11423 vss 76.29fF $ **FLOATING
C1560 vdd.n11424 vss 76.29fF $ **FLOATING
C1561 vdd.n11425 vss 76.29fF $ **FLOATING
C1562 vdd.n11426 vss 76.29fF $ **FLOATING
C1563 vdd.n11427 vss 76.29fF $ **FLOATING
C1564 vdd.n11428 vss 76.29fF $ **FLOATING
C1565 vdd.n11429 vss 76.29fF $ **FLOATING
C1566 vdd.n11430 vss 76.29fF $ **FLOATING
C1567 vdd.n11431 vss 76.29fF $ **FLOATING
C1568 vdd.n11432 vss 76.29fF $ **FLOATING
C1569 vdd.n11433 vss 76.29fF $ **FLOATING
C1570 vdd.n11434 vss 76.29fF $ **FLOATING
C1571 vdd.n11435 vss 76.29fF $ **FLOATING
C1572 vdd.n11436 vss 76.29fF $ **FLOATING
C1573 vdd.n11437 vss 76.29fF $ **FLOATING
C1574 vdd.n11438 vss 76.29fF $ **FLOATING
C1575 vdd.n11439 vss 76.29fF $ **FLOATING
C1576 vdd.n11440 vss 76.29fF $ **FLOATING
C1577 vdd.n11441 vss 76.29fF $ **FLOATING
C1578 vdd.n11442 vss 76.29fF $ **FLOATING
C1579 vdd.n11443 vss 76.29fF $ **FLOATING
C1580 vdd.n11444 vss 76.29fF $ **FLOATING
C1581 vdd.n11445 vss 76.29fF $ **FLOATING
C1582 vdd.n11446 vss 76.29fF $ **FLOATING
C1583 vdd.n11447 vss 76.29fF $ **FLOATING
C1584 vdd.n11448 vss 76.29fF $ **FLOATING
C1585 vdd.n11449 vss 76.29fF $ **FLOATING
C1586 vdd.n11450 vss 76.29fF $ **FLOATING
C1587 vdd.n11451 vss 76.29fF $ **FLOATING
C1588 vdd.n11452 vss 76.29fF $ **FLOATING
C1589 vdd.n11453 vss 76.29fF $ **FLOATING
C1590 vdd.n11454 vss 76.29fF $ **FLOATING
C1591 vdd.n11455 vss 76.29fF $ **FLOATING
C1592 vdd.n11456 vss 76.29fF $ **FLOATING
C1593 vdd.n11457 vss 76.29fF $ **FLOATING
C1594 vdd.n11458 vss 76.29fF $ **FLOATING
C1595 vdd.n11459 vss 76.29fF $ **FLOATING
C1596 vdd.n11460 vss 76.29fF $ **FLOATING
C1597 vdd.n11461 vss 76.29fF $ **FLOATING
C1598 vdd.n11462 vss 76.29fF $ **FLOATING
C1599 vdd.n11463 vss 76.29fF $ **FLOATING
C1600 vdd.n11464 vss 76.29fF $ **FLOATING
C1601 vdd.n11465 vss 76.29fF $ **FLOATING
C1602 vdd.n11466 vss 76.29fF $ **FLOATING
C1603 vdd.n11467 vss 76.29fF $ **FLOATING
C1604 vdd.n11468 vss 76.29fF $ **FLOATING
C1605 vdd.n11469 vss 76.29fF $ **FLOATING
C1606 vdd.n11470 vss 76.29fF $ **FLOATING
C1607 vdd.n11471 vss 76.29fF $ **FLOATING
C1608 vdd.n11472 vss 76.29fF $ **FLOATING
C1609 vdd.n11473 vss 76.29fF $ **FLOATING
C1610 vdd.n11474 vss 76.29fF $ **FLOATING
C1611 vdd.n11475 vss 76.29fF $ **FLOATING
C1612 vdd.n11476 vss 76.29fF $ **FLOATING
C1613 vdd.n11477 vss 76.29fF $ **FLOATING
C1614 vdd.n11478 vss 52.84fF $ **FLOATING
C1615 vdd.n11624 vss 5.17fF $ **FLOATING
C1616 vdd.n11625 vss 5.17fF $ **FLOATING
C1617 vdd.n11629 vss 7.24fF $ **FLOATING
C1618 vdd.n11630 vss 7.48fF $ **FLOATING
C1619 vdd.n11631 vss 7.48fF $ **FLOATING
C1620 vdd.n11632 vss 7.48fF $ **FLOATING
C1621 vdd.n11633 vss 7.48fF $ **FLOATING
C1622 vdd.n11634 vss 7.48fF $ **FLOATING
C1623 vdd.n11635 vss 7.48fF $ **FLOATING
C1624 vdd.n11636 vss 7.48fF $ **FLOATING
C1625 vdd.n11637 vss 7.48fF $ **FLOATING
C1626 vdd.n11638 vss 7.48fF $ **FLOATING
C1627 vdd.n11639 vss 7.48fF $ **FLOATING
C1628 vdd.n11640 vss 7.48fF $ **FLOATING
C1629 vdd.n11641 vss 7.48fF $ **FLOATING
C1630 vdd.n11642 vss 7.48fF $ **FLOATING
C1631 vdd.n11643 vss 7.48fF $ **FLOATING
C1632 vdd.n11644 vss 7.48fF $ **FLOATING
C1633 vdd.n11645 vss 7.48fF $ **FLOATING
C1634 vdd.n11646 vss 7.48fF $ **FLOATING
C1635 vdd.n11647 vss 7.48fF $ **FLOATING
C1636 vdd.n11655 vss 5.17fF $ **FLOATING
C1637 vdd.n11656 vss 5.17fF $ **FLOATING
C1638 vdd.n11658 vss 7.28fF $ **FLOATING
C1639 vdd.n11804 vss 5.17fF $ **FLOATING
C1640 vdd.n11805 vss 5.17fF $ **FLOATING
C1641 vdd.n11809 vss 7.24fF $ **FLOATING
C1642 vdd.n11810 vss 7.48fF $ **FLOATING
C1643 vdd.n11811 vss 7.48fF $ **FLOATING
C1644 vdd.n11812 vss 7.48fF $ **FLOATING
C1645 vdd.n11813 vss 7.48fF $ **FLOATING
C1646 vdd.n11814 vss 7.48fF $ **FLOATING
C1647 vdd.n11815 vss 7.48fF $ **FLOATING
C1648 vdd.n11816 vss 7.48fF $ **FLOATING
C1649 vdd.n11817 vss 7.48fF $ **FLOATING
C1650 vdd.n11818 vss 7.48fF $ **FLOATING
C1651 vdd.n11819 vss 7.48fF $ **FLOATING
C1652 vdd.n11820 vss 7.48fF $ **FLOATING
C1653 vdd.n11821 vss 7.48fF $ **FLOATING
C1654 vdd.n11822 vss 7.48fF $ **FLOATING
C1655 vdd.n11823 vss 7.48fF $ **FLOATING
C1656 vdd.n11824 vss 7.48fF $ **FLOATING
C1657 vdd.n11825 vss 7.48fF $ **FLOATING
C1658 vdd.n11826 vss 7.48fF $ **FLOATING
C1659 vdd.n11827 vss 7.48fF $ **FLOATING
C1660 vdd.n11835 vss 5.17fF $ **FLOATING
C1661 vdd.n11836 vss 5.17fF $ **FLOATING
C1662 vdd.n11838 vss 7.28fF $ **FLOATING
C1663 vdd.n11984 vss 5.17fF $ **FLOATING
C1664 vdd.n11985 vss 5.17fF $ **FLOATING
C1665 vdd.n11989 vss 7.24fF $ **FLOATING
C1666 vdd.n11990 vss 7.48fF $ **FLOATING
C1667 vdd.n11991 vss 7.48fF $ **FLOATING
C1668 vdd.n11992 vss 7.48fF $ **FLOATING
C1669 vdd.n11993 vss 7.48fF $ **FLOATING
C1670 vdd.n11994 vss 7.48fF $ **FLOATING
C1671 vdd.n11995 vss 7.48fF $ **FLOATING
C1672 vdd.n11996 vss 7.48fF $ **FLOATING
C1673 vdd.n11997 vss 7.48fF $ **FLOATING
C1674 vdd.n11998 vss 7.48fF $ **FLOATING
C1675 vdd.n11999 vss 7.48fF $ **FLOATING
C1676 vdd.n12000 vss 7.48fF $ **FLOATING
C1677 vdd.n12001 vss 7.48fF $ **FLOATING
C1678 vdd.n12002 vss 7.48fF $ **FLOATING
C1679 vdd.n12003 vss 7.48fF $ **FLOATING
C1680 vdd.n12004 vss 7.48fF $ **FLOATING
C1681 vdd.n12005 vss 7.48fF $ **FLOATING
C1682 vdd.n12006 vss 7.48fF $ **FLOATING
C1683 vdd.n12007 vss 7.48fF $ **FLOATING
C1684 vdd.n12015 vss 5.17fF $ **FLOATING
C1685 vdd.n12016 vss 5.17fF $ **FLOATING
C1686 vdd.n12018 vss 7.28fF $ **FLOATING
C1687 vdd.n12164 vss 5.17fF $ **FLOATING
C1688 vdd.n12165 vss 5.17fF $ **FLOATING
C1689 vdd.n12169 vss 7.24fF $ **FLOATING
C1690 vdd.n12170 vss 7.48fF $ **FLOATING
C1691 vdd.n12171 vss 7.48fF $ **FLOATING
C1692 vdd.n12172 vss 7.48fF $ **FLOATING
C1693 vdd.n12173 vss 7.48fF $ **FLOATING
C1694 vdd.n12174 vss 7.48fF $ **FLOATING
C1695 vdd.n12175 vss 7.48fF $ **FLOATING
C1696 vdd.n12176 vss 7.48fF $ **FLOATING
C1697 vdd.n12177 vss 7.48fF $ **FLOATING
C1698 vdd.n12178 vss 7.48fF $ **FLOATING
C1699 vdd.n12179 vss 7.48fF $ **FLOATING
C1700 vdd.n12180 vss 7.48fF $ **FLOATING
C1701 vdd.n12181 vss 7.48fF $ **FLOATING
C1702 vdd.n12182 vss 7.48fF $ **FLOATING
C1703 vdd.n12183 vss 7.48fF $ **FLOATING
C1704 vdd.n12184 vss 7.48fF $ **FLOATING
C1705 vdd.n12185 vss 7.48fF $ **FLOATING
C1706 vdd.n12186 vss 7.48fF $ **FLOATING
C1707 vdd.n12187 vss 7.48fF $ **FLOATING
C1708 vdd.n12195 vss 5.17fF $ **FLOATING
C1709 vdd.n12196 vss 5.17fF $ **FLOATING
C1710 vdd.n12198 vss 7.28fF $ **FLOATING
C1711 vdd.n12344 vss 5.17fF $ **FLOATING
C1712 vdd.n12345 vss 5.17fF $ **FLOATING
C1713 vdd.n12349 vss 7.24fF $ **FLOATING
C1714 vdd.n12350 vss 7.48fF $ **FLOATING
C1715 vdd.n12351 vss 7.48fF $ **FLOATING
C1716 vdd.n12352 vss 7.48fF $ **FLOATING
C1717 vdd.n12353 vss 7.48fF $ **FLOATING
C1718 vdd.n12354 vss 7.48fF $ **FLOATING
C1719 vdd.n12355 vss 7.48fF $ **FLOATING
C1720 vdd.n12356 vss 7.48fF $ **FLOATING
C1721 vdd.n12357 vss 7.48fF $ **FLOATING
C1722 vdd.n12358 vss 7.48fF $ **FLOATING
C1723 vdd.n12359 vss 7.48fF $ **FLOATING
C1724 vdd.n12360 vss 7.48fF $ **FLOATING
C1725 vdd.n12361 vss 7.48fF $ **FLOATING
C1726 vdd.n12362 vss 7.48fF $ **FLOATING
C1727 vdd.n12363 vss 7.48fF $ **FLOATING
C1728 vdd.n12364 vss 7.48fF $ **FLOATING
C1729 vdd.n12365 vss 7.48fF $ **FLOATING
C1730 vdd.n12366 vss 7.48fF $ **FLOATING
C1731 vdd.n12367 vss 7.48fF $ **FLOATING
C1732 vdd.n12375 vss 5.17fF $ **FLOATING
C1733 vdd.n12376 vss 5.17fF $ **FLOATING
C1734 vdd.n12378 vss 7.28fF $ **FLOATING
C1735 vdd.n12524 vss 5.17fF $ **FLOATING
C1736 vdd.n12525 vss 5.17fF $ **FLOATING
C1737 vdd.n12529 vss 7.24fF $ **FLOATING
C1738 vdd.n12530 vss 7.48fF $ **FLOATING
C1739 vdd.n12531 vss 7.48fF $ **FLOATING
C1740 vdd.n12532 vss 7.48fF $ **FLOATING
C1741 vdd.n12533 vss 7.48fF $ **FLOATING
C1742 vdd.n12534 vss 7.48fF $ **FLOATING
C1743 vdd.n12535 vss 7.48fF $ **FLOATING
C1744 vdd.n12536 vss 7.48fF $ **FLOATING
C1745 vdd.n12537 vss 7.48fF $ **FLOATING
C1746 vdd.n12538 vss 7.48fF $ **FLOATING
C1747 vdd.n12539 vss 7.48fF $ **FLOATING
C1748 vdd.n12540 vss 7.48fF $ **FLOATING
C1749 vdd.n12541 vss 7.48fF $ **FLOATING
C1750 vdd.n12542 vss 7.48fF $ **FLOATING
C1751 vdd.n12543 vss 7.48fF $ **FLOATING
C1752 vdd.n12544 vss 7.48fF $ **FLOATING
C1753 vdd.n12545 vss 7.48fF $ **FLOATING
C1754 vdd.n12546 vss 7.48fF $ **FLOATING
C1755 vdd.n12547 vss 7.48fF $ **FLOATING
C1756 vdd.n12555 vss 5.17fF $ **FLOATING
C1757 vdd.n12556 vss 5.17fF $ **FLOATING
C1758 vdd.n12558 vss 7.28fF $ **FLOATING
C1759 vdd.n12704 vss 5.17fF $ **FLOATING
C1760 vdd.n12705 vss 5.17fF $ **FLOATING
C1761 vdd.n12709 vss 7.24fF $ **FLOATING
C1762 vdd.n12710 vss 7.48fF $ **FLOATING
C1763 vdd.n12711 vss 7.48fF $ **FLOATING
C1764 vdd.n12712 vss 7.48fF $ **FLOATING
C1765 vdd.n12713 vss 7.48fF $ **FLOATING
C1766 vdd.n12714 vss 7.48fF $ **FLOATING
C1767 vdd.n12715 vss 7.48fF $ **FLOATING
C1768 vdd.n12716 vss 7.48fF $ **FLOATING
C1769 vdd.n12717 vss 7.48fF $ **FLOATING
C1770 vdd.n12718 vss 7.48fF $ **FLOATING
C1771 vdd.n12719 vss 7.48fF $ **FLOATING
C1772 vdd.n12720 vss 7.48fF $ **FLOATING
C1773 vdd.n12721 vss 7.48fF $ **FLOATING
C1774 vdd.n12722 vss 7.48fF $ **FLOATING
C1775 vdd.n12723 vss 7.48fF $ **FLOATING
C1776 vdd.n12724 vss 7.48fF $ **FLOATING
C1777 vdd.n12725 vss 7.48fF $ **FLOATING
C1778 vdd.n12726 vss 7.48fF $ **FLOATING
C1779 vdd.n12727 vss 7.48fF $ **FLOATING
C1780 vdd.n12735 vss 5.17fF $ **FLOATING
C1781 vdd.n12736 vss 5.17fF $ **FLOATING
C1782 vdd.n12738 vss 7.28fF $ **FLOATING
C1783 vdd.n12884 vss 5.17fF $ **FLOATING
C1784 vdd.n12885 vss 5.17fF $ **FLOATING
C1785 vdd.n12889 vss 7.24fF $ **FLOATING
C1786 vdd.n12890 vss 7.48fF $ **FLOATING
C1787 vdd.n12891 vss 7.48fF $ **FLOATING
C1788 vdd.n12892 vss 7.48fF $ **FLOATING
C1789 vdd.n12893 vss 7.48fF $ **FLOATING
C1790 vdd.n12894 vss 7.48fF $ **FLOATING
C1791 vdd.n12895 vss 7.48fF $ **FLOATING
C1792 vdd.n12896 vss 7.48fF $ **FLOATING
C1793 vdd.n12897 vss 7.48fF $ **FLOATING
C1794 vdd.n12898 vss 7.48fF $ **FLOATING
C1795 vdd.n12899 vss 7.48fF $ **FLOATING
C1796 vdd.n12900 vss 7.48fF $ **FLOATING
C1797 vdd.n12901 vss 7.48fF $ **FLOATING
C1798 vdd.n12902 vss 7.48fF $ **FLOATING
C1799 vdd.n12903 vss 7.48fF $ **FLOATING
C1800 vdd.n12904 vss 7.48fF $ **FLOATING
C1801 vdd.n12905 vss 7.48fF $ **FLOATING
C1802 vdd.n12906 vss 7.48fF $ **FLOATING
C1803 vdd.n12907 vss 7.48fF $ **FLOATING
C1804 vdd.n12915 vss 5.17fF $ **FLOATING
C1805 vdd.n12916 vss 5.17fF $ **FLOATING
C1806 vdd.n12918 vss 7.28fF $ **FLOATING
C1807 vdd.n13064 vss 5.17fF $ **FLOATING
C1808 vdd.n13065 vss 5.17fF $ **FLOATING
C1809 vdd.n13069 vss 7.24fF $ **FLOATING
C1810 vdd.n13070 vss 7.48fF $ **FLOATING
C1811 vdd.n13071 vss 7.48fF $ **FLOATING
C1812 vdd.n13072 vss 7.48fF $ **FLOATING
C1813 vdd.n13073 vss 7.48fF $ **FLOATING
C1814 vdd.n13074 vss 7.48fF $ **FLOATING
C1815 vdd.n13075 vss 7.48fF $ **FLOATING
C1816 vdd.n13076 vss 7.48fF $ **FLOATING
C1817 vdd.n13077 vss 7.48fF $ **FLOATING
C1818 vdd.n13078 vss 7.48fF $ **FLOATING
C1819 vdd.n13079 vss 7.48fF $ **FLOATING
C1820 vdd.n13080 vss 7.48fF $ **FLOATING
C1821 vdd.n13081 vss 7.48fF $ **FLOATING
C1822 vdd.n13082 vss 7.48fF $ **FLOATING
C1823 vdd.n13083 vss 7.48fF $ **FLOATING
C1824 vdd.n13084 vss 7.48fF $ **FLOATING
C1825 vdd.n13085 vss 7.48fF $ **FLOATING
C1826 vdd.n13086 vss 7.48fF $ **FLOATING
C1827 vdd.n13087 vss 7.48fF $ **FLOATING
C1828 vdd.n13095 vss 5.17fF $ **FLOATING
C1829 vdd.n13096 vss 5.17fF $ **FLOATING
C1830 vdd.n13098 vss 7.28fF $ **FLOATING
C1831 vdd.n13244 vss 5.17fF $ **FLOATING
C1832 vdd.n13245 vss 5.17fF $ **FLOATING
C1833 vdd.n13249 vss 7.24fF $ **FLOATING
C1834 vdd.n13250 vss 7.48fF $ **FLOATING
C1835 vdd.n13251 vss 7.48fF $ **FLOATING
C1836 vdd.n13252 vss 7.48fF $ **FLOATING
C1837 vdd.n13253 vss 7.48fF $ **FLOATING
C1838 vdd.n13254 vss 7.48fF $ **FLOATING
C1839 vdd.n13255 vss 7.48fF $ **FLOATING
C1840 vdd.n13256 vss 7.48fF $ **FLOATING
C1841 vdd.n13257 vss 7.48fF $ **FLOATING
C1842 vdd.n13258 vss 7.48fF $ **FLOATING
C1843 vdd.n13259 vss 7.48fF $ **FLOATING
C1844 vdd.n13260 vss 7.48fF $ **FLOATING
C1845 vdd.n13261 vss 7.48fF $ **FLOATING
C1846 vdd.n13262 vss 7.48fF $ **FLOATING
C1847 vdd.n13263 vss 7.48fF $ **FLOATING
C1848 vdd.n13264 vss 7.48fF $ **FLOATING
C1849 vdd.n13265 vss 7.48fF $ **FLOATING
C1850 vdd.n13266 vss 7.48fF $ **FLOATING
C1851 vdd.n13267 vss 7.48fF $ **FLOATING
C1852 vdd.n13275 vss 5.17fF $ **FLOATING
C1853 vdd.n13276 vss 5.17fF $ **FLOATING
C1854 vdd.n13278 vss 7.28fF $ **FLOATING
C1855 vdd.n13424 vss 5.17fF $ **FLOATING
C1856 vdd.n13425 vss 5.17fF $ **FLOATING
C1857 vdd.n13429 vss 7.24fF $ **FLOATING
C1858 vdd.n13430 vss 7.48fF $ **FLOATING
C1859 vdd.n13431 vss 7.48fF $ **FLOATING
C1860 vdd.n13432 vss 7.48fF $ **FLOATING
C1861 vdd.n13433 vss 7.48fF $ **FLOATING
C1862 vdd.n13434 vss 7.48fF $ **FLOATING
C1863 vdd.n13435 vss 7.48fF $ **FLOATING
C1864 vdd.n13436 vss 7.48fF $ **FLOATING
C1865 vdd.n13437 vss 7.48fF $ **FLOATING
C1866 vdd.n13438 vss 7.48fF $ **FLOATING
C1867 vdd.n13439 vss 7.48fF $ **FLOATING
C1868 vdd.n13440 vss 7.48fF $ **FLOATING
C1869 vdd.n13441 vss 7.48fF $ **FLOATING
C1870 vdd.n13442 vss 7.48fF $ **FLOATING
C1871 vdd.n13443 vss 7.48fF $ **FLOATING
C1872 vdd.n13444 vss 7.48fF $ **FLOATING
C1873 vdd.n13445 vss 7.48fF $ **FLOATING
C1874 vdd.n13446 vss 7.48fF $ **FLOATING
C1875 vdd.n13447 vss 7.48fF $ **FLOATING
C1876 vdd.n13455 vss 5.17fF $ **FLOATING
C1877 vdd.n13456 vss 5.17fF $ **FLOATING
C1878 vdd.n13458 vss 7.28fF $ **FLOATING
C1879 vdd.n13477 vss 5.36fF $ **FLOATING
C1880 vdd.n13478 vss 4.17fF $ **FLOATING
C1881 vdd.n13481 vss 4.34fF $ **FLOATING
C1882 vdd.n13484 vss 4.34fF $ **FLOATING
C1883 vdd.n13487 vss 4.34fF $ **FLOATING
C1884 vdd.n13490 vss 4.34fF $ **FLOATING
C1885 vdd.n13493 vss 4.34fF $ **FLOATING
C1886 vdd.n13496 vss 4.34fF $ **FLOATING
C1887 vdd.n13499 vss 4.34fF $ **FLOATING
C1888 vdd.n13502 vss 4.34fF $ **FLOATING
C1889 vdd.n13505 vss 4.34fF $ **FLOATING
C1890 vdd.n13506 vss 4.34fF $ **FLOATING
C1891 vdd.n13509 vss 4.34fF $ **FLOATING
C1892 vdd.n13512 vss 4.34fF $ **FLOATING
C1893 vdd.n13515 vss 4.34fF $ **FLOATING
C1894 vdd.n13518 vss 4.34fF $ **FLOATING
C1895 vdd.n13521 vss 4.34fF $ **FLOATING
C1896 vdd.n13524 vss 4.34fF $ **FLOATING
C1897 vdd.n13527 vss 4.34fF $ **FLOATING
C1898 vdd.n13530 vss 4.34fF $ **FLOATING
C1899 vdd.n13533 vss 5.36fF $ **FLOATING
C1900 vdd.n13534 vss 5.68fF $ **FLOATING
C1901 vdd.n13535 vss 172.67fF $ **FLOATING
C1902 vdd.n13536 vss 76.29fF $ **FLOATING
C1903 vdd.n13537 vss 76.29fF $ **FLOATING
C1904 vdd.n13538 vss 76.29fF $ **FLOATING
C1905 vdd.n13539 vss 76.29fF $ **FLOATING
C1906 vdd.n13540 vss 76.29fF $ **FLOATING
C1907 vdd.n13541 vss 76.29fF $ **FLOATING
C1908 vdd.n13542 vss 76.29fF $ **FLOATING
C1909 vdd.n13543 vss 76.29fF $ **FLOATING
C1910 vdd.n13544 vss 76.29fF $ **FLOATING
C1911 vdd.n13545 vss 62.46fF $ **FLOATING
C1912 out_p.n0 vss 4.40fF $ **FLOATING
C1913 out_p.n1 vss 4.56fF $ **FLOATING
C1914 out_p.n2 vss 4.56fF $ **FLOATING
C1915 out_p.n3 vss 4.56fF $ **FLOATING
C1916 out_p.n4 vss 4.56fF $ **FLOATING
C1917 out_p.n5 vss 4.56fF $ **FLOATING
C1918 out_p.n6 vss 4.56fF $ **FLOATING
C1919 out_p.n7 vss 4.56fF $ **FLOATING
C1920 out_p.n8 vss 4.56fF $ **FLOATING
C1921 out_p.n9 vss 4.56fF $ **FLOATING
C1922 out_p.n10 vss 4.56fF $ **FLOATING
C1923 out_p.n11 vss 4.56fF $ **FLOATING
C1924 out_p.n12 vss 4.56fF $ **FLOATING
C1925 out_p.n13 vss 4.56fF $ **FLOATING
C1926 out_p.n14 vss 4.56fF $ **FLOATING
C1927 out_p.n15 vss 4.56fF $ **FLOATING
C1928 out_p.n16 vss 4.56fF $ **FLOATING
C1929 out_p.n17 vss 4.56fF $ **FLOATING
C1930 out_p.n18 vss 4.56fF $ **FLOATING
C1931 out_p.n19 vss 4.27fF $ **FLOATING
C1932 out_p.n20 vss 4.37fF $ **FLOATING
C1933 out_p.n21 vss 4.53fF $ **FLOATING
C1934 out_p.n22 vss 4.53fF $ **FLOATING
C1935 out_p.n23 vss 4.26fF $ **FLOATING
C1936 out_p.n24 vss 4.40fF $ **FLOATING
C1937 out_p.n25 vss 4.56fF $ **FLOATING
C1938 out_p.n26 vss 4.56fF $ **FLOATING
C1939 out_p.n27 vss 4.56fF $ **FLOATING
C1940 out_p.n28 vss 4.56fF $ **FLOATING
C1941 out_p.n29 vss 4.56fF $ **FLOATING
C1942 out_p.n30 vss 4.56fF $ **FLOATING
C1943 out_p.n31 vss 4.56fF $ **FLOATING
C1944 out_p.n32 vss 4.56fF $ **FLOATING
C1945 out_p.n33 vss 4.56fF $ **FLOATING
C1946 out_p.n34 vss 4.56fF $ **FLOATING
C1947 out_p.n35 vss 4.56fF $ **FLOATING
C1948 out_p.n36 vss 4.56fF $ **FLOATING
C1949 out_p.n37 vss 4.56fF $ **FLOATING
C1950 out_p.n38 vss 4.56fF $ **FLOATING
C1951 out_p.n39 vss 4.56fF $ **FLOATING
C1952 out_p.n40 vss 4.56fF $ **FLOATING
C1953 out_p.n41 vss 4.56fF $ **FLOATING
C1954 out_p.n42 vss 4.56fF $ **FLOATING
C1955 out_p.n43 vss 4.27fF $ **FLOATING
C1956 out_p.n44 vss 4.37fF $ **FLOATING
C1957 out_p.n45 vss 4.53fF $ **FLOATING
C1958 out_p.n46 vss 4.53fF $ **FLOATING
C1959 out_p.n47 vss 4.26fF $ **FLOATING
C1960 out_p.n48 vss 4.40fF $ **FLOATING
C1961 out_p.n49 vss 4.56fF $ **FLOATING
C1962 out_p.n50 vss 4.56fF $ **FLOATING
C1963 out_p.n51 vss 4.56fF $ **FLOATING
C1964 out_p.n52 vss 4.56fF $ **FLOATING
C1965 out_p.n53 vss 4.56fF $ **FLOATING
C1966 out_p.n54 vss 4.56fF $ **FLOATING
C1967 out_p.n55 vss 4.56fF $ **FLOATING
C1968 out_p.n56 vss 4.56fF $ **FLOATING
C1969 out_p.n57 vss 4.56fF $ **FLOATING
C1970 out_p.n58 vss 4.56fF $ **FLOATING
C1971 out_p.n59 vss 4.56fF $ **FLOATING
C1972 out_p.n60 vss 4.56fF $ **FLOATING
C1973 out_p.n61 vss 4.56fF $ **FLOATING
C1974 out_p.n62 vss 4.56fF $ **FLOATING
C1975 out_p.n63 vss 4.56fF $ **FLOATING
C1976 out_p.n64 vss 4.56fF $ **FLOATING
C1977 out_p.n65 vss 4.56fF $ **FLOATING
C1978 out_p.n66 vss 4.56fF $ **FLOATING
C1979 out_p.n67 vss 4.27fF $ **FLOATING
C1980 out_p.n68 vss 4.37fF $ **FLOATING
C1981 out_p.n69 vss 4.53fF $ **FLOATING
C1982 out_p.n70 vss 4.53fF $ **FLOATING
C1983 out_p.n71 vss 4.26fF $ **FLOATING
C1984 out_p.n72 vss 4.40fF $ **FLOATING
C1985 out_p.n73 vss 4.56fF $ **FLOATING
C1986 out_p.n74 vss 4.56fF $ **FLOATING
C1987 out_p.n75 vss 4.56fF $ **FLOATING
C1988 out_p.n76 vss 4.56fF $ **FLOATING
C1989 out_p.n77 vss 4.56fF $ **FLOATING
C1990 out_p.n78 vss 4.56fF $ **FLOATING
C1991 out_p.n79 vss 4.56fF $ **FLOATING
C1992 out_p.n80 vss 4.56fF $ **FLOATING
C1993 out_p.n81 vss 4.56fF $ **FLOATING
C1994 out_p.n82 vss 4.56fF $ **FLOATING
C1995 out_p.n83 vss 4.56fF $ **FLOATING
C1996 out_p.n84 vss 4.56fF $ **FLOATING
C1997 out_p.n85 vss 4.56fF $ **FLOATING
C1998 out_p.n86 vss 4.56fF $ **FLOATING
C1999 out_p.n87 vss 4.56fF $ **FLOATING
C2000 out_p.n88 vss 4.56fF $ **FLOATING
C2001 out_p.n89 vss 4.56fF $ **FLOATING
C2002 out_p.n90 vss 4.56fF $ **FLOATING
C2003 out_p.n91 vss 4.27fF $ **FLOATING
C2004 out_p.n92 vss 4.37fF $ **FLOATING
C2005 out_p.n93 vss 4.53fF $ **FLOATING
C2006 out_p.n94 vss 4.53fF $ **FLOATING
C2007 out_p.n95 vss 4.26fF $ **FLOATING
C2008 out_p.n96 vss 4.40fF $ **FLOATING
C2009 out_p.n97 vss 4.56fF $ **FLOATING
C2010 out_p.n98 vss 4.56fF $ **FLOATING
C2011 out_p.n99 vss 4.56fF $ **FLOATING
C2012 out_p.n100 vss 4.56fF $ **FLOATING
C2013 out_p.n101 vss 4.56fF $ **FLOATING
C2014 out_p.n102 vss 4.56fF $ **FLOATING
C2015 out_p.n103 vss 4.56fF $ **FLOATING
C2016 out_p.n104 vss 4.56fF $ **FLOATING
C2017 out_p.n105 vss 4.56fF $ **FLOATING
C2018 out_p.n106 vss 4.56fF $ **FLOATING
C2019 out_p.n107 vss 4.56fF $ **FLOATING
C2020 out_p.n108 vss 4.56fF $ **FLOATING
C2021 out_p.n109 vss 4.56fF $ **FLOATING
C2022 out_p.n110 vss 4.56fF $ **FLOATING
C2023 out_p.n111 vss 4.56fF $ **FLOATING
C2024 out_p.n112 vss 4.56fF $ **FLOATING
C2025 out_p.n113 vss 4.56fF $ **FLOATING
C2026 out_p.n114 vss 4.56fF $ **FLOATING
C2027 out_p.n115 vss 4.27fF $ **FLOATING
C2028 out_p.n116 vss 4.37fF $ **FLOATING
C2029 out_p.n117 vss 4.53fF $ **FLOATING
C2030 out_p.n118 vss 4.53fF $ **FLOATING
C2031 out_p.n119 vss 4.26fF $ **FLOATING
C2032 out_p.n120 vss 4.40fF $ **FLOATING
C2033 out_p.n121 vss 4.56fF $ **FLOATING
C2034 out_p.n122 vss 4.56fF $ **FLOATING
C2035 out_p.n123 vss 4.56fF $ **FLOATING
C2036 out_p.n124 vss 4.56fF $ **FLOATING
C2037 out_p.n125 vss 4.56fF $ **FLOATING
C2038 out_p.n126 vss 4.56fF $ **FLOATING
C2039 out_p.n127 vss 4.56fF $ **FLOATING
C2040 out_p.n128 vss 4.56fF $ **FLOATING
C2041 out_p.n129 vss 4.56fF $ **FLOATING
C2042 out_p.n130 vss 4.56fF $ **FLOATING
C2043 out_p.n131 vss 4.56fF $ **FLOATING
C2044 out_p.n132 vss 4.56fF $ **FLOATING
C2045 out_p.n133 vss 4.56fF $ **FLOATING
C2046 out_p.n134 vss 4.56fF $ **FLOATING
C2047 out_p.n135 vss 4.56fF $ **FLOATING
C2048 out_p.n136 vss 4.56fF $ **FLOATING
C2049 out_p.n137 vss 4.56fF $ **FLOATING
C2050 out_p.n138 vss 4.56fF $ **FLOATING
C2051 out_p.n139 vss 4.27fF $ **FLOATING
C2052 out_p.n140 vss 4.37fF $ **FLOATING
C2053 out_p.n141 vss 4.53fF $ **FLOATING
C2054 out_p.n142 vss 4.53fF $ **FLOATING
C2055 out_p.n143 vss 4.26fF $ **FLOATING
C2056 out_p.n144 vss 4.40fF $ **FLOATING
C2057 out_p.n145 vss 4.56fF $ **FLOATING
C2058 out_p.n146 vss 4.56fF $ **FLOATING
C2059 out_p.n147 vss 4.56fF $ **FLOATING
C2060 out_p.n148 vss 4.56fF $ **FLOATING
C2061 out_p.n149 vss 4.56fF $ **FLOATING
C2062 out_p.n150 vss 4.56fF $ **FLOATING
C2063 out_p.n151 vss 4.56fF $ **FLOATING
C2064 out_p.n152 vss 4.56fF $ **FLOATING
C2065 out_p.n153 vss 4.56fF $ **FLOATING
C2066 out_p.n154 vss 4.56fF $ **FLOATING
C2067 out_p.n155 vss 4.56fF $ **FLOATING
C2068 out_p.n156 vss 4.56fF $ **FLOATING
C2069 out_p.n157 vss 4.56fF $ **FLOATING
C2070 out_p.n158 vss 4.56fF $ **FLOATING
C2071 out_p.n159 vss 4.56fF $ **FLOATING
C2072 out_p.n160 vss 4.56fF $ **FLOATING
C2073 out_p.n161 vss 4.56fF $ **FLOATING
C2074 out_p.n162 vss 4.56fF $ **FLOATING
C2075 out_p.n163 vss 4.27fF $ **FLOATING
C2076 out_p.n164 vss 4.37fF $ **FLOATING
C2077 out_p.n165 vss 4.53fF $ **FLOATING
C2078 out_p.n166 vss 4.53fF $ **FLOATING
C2079 out_p.n167 vss 4.26fF $ **FLOATING
C2080 out_p.n168 vss 4.40fF $ **FLOATING
C2081 out_p.n169 vss 4.56fF $ **FLOATING
C2082 out_p.n170 vss 4.56fF $ **FLOATING
C2083 out_p.n171 vss 4.56fF $ **FLOATING
C2084 out_p.n172 vss 4.56fF $ **FLOATING
C2085 out_p.n173 vss 4.56fF $ **FLOATING
C2086 out_p.n174 vss 4.56fF $ **FLOATING
C2087 out_p.n175 vss 4.56fF $ **FLOATING
C2088 out_p.n176 vss 4.56fF $ **FLOATING
C2089 out_p.n177 vss 4.56fF $ **FLOATING
C2090 out_p.n178 vss 4.56fF $ **FLOATING
C2091 out_p.n179 vss 4.56fF $ **FLOATING
C2092 out_p.n180 vss 4.56fF $ **FLOATING
C2093 out_p.n181 vss 4.56fF $ **FLOATING
C2094 out_p.n182 vss 4.56fF $ **FLOATING
C2095 out_p.n183 vss 4.56fF $ **FLOATING
C2096 out_p.n184 vss 4.56fF $ **FLOATING
C2097 out_p.n185 vss 4.56fF $ **FLOATING
C2098 out_p.n186 vss 4.56fF $ **FLOATING
C2099 out_p.n187 vss 4.27fF $ **FLOATING
C2100 out_p.n188 vss 4.37fF $ **FLOATING
C2101 out_p.n189 vss 4.53fF $ **FLOATING
C2102 out_p.n190 vss 4.53fF $ **FLOATING
C2103 out_p.n191 vss 4.26fF $ **FLOATING
C2104 out_p.n192 vss 4.40fF $ **FLOATING
C2105 out_p.n193 vss 4.56fF $ **FLOATING
C2106 out_p.n194 vss 4.56fF $ **FLOATING
C2107 out_p.n195 vss 4.56fF $ **FLOATING
C2108 out_p.n196 vss 4.56fF $ **FLOATING
C2109 out_p.n197 vss 4.56fF $ **FLOATING
C2110 out_p.n198 vss 4.56fF $ **FLOATING
C2111 out_p.n199 vss 4.56fF $ **FLOATING
C2112 out_p.n200 vss 4.56fF $ **FLOATING
C2113 out_p.n201 vss 4.56fF $ **FLOATING
C2114 out_p.n202 vss 4.56fF $ **FLOATING
C2115 out_p.n203 vss 4.56fF $ **FLOATING
C2116 out_p.n204 vss 4.56fF $ **FLOATING
C2117 out_p.n205 vss 4.56fF $ **FLOATING
C2118 out_p.n206 vss 4.56fF $ **FLOATING
C2119 out_p.n207 vss 4.56fF $ **FLOATING
C2120 out_p.n208 vss 4.56fF $ **FLOATING
C2121 out_p.n209 vss 4.56fF $ **FLOATING
C2122 out_p.n210 vss 4.56fF $ **FLOATING
C2123 out_p.n211 vss 4.27fF $ **FLOATING
C2124 out_p.n212 vss 4.37fF $ **FLOATING
C2125 out_p.n213 vss 4.53fF $ **FLOATING
C2126 out_p.n214 vss 4.53fF $ **FLOATING
C2127 out_p.n215 vss 4.26fF $ **FLOATING
C2128 out_p.n216 vss 4.40fF $ **FLOATING
C2129 out_p.n217 vss 4.56fF $ **FLOATING
C2130 out_p.n218 vss 4.56fF $ **FLOATING
C2131 out_p.n219 vss 4.56fF $ **FLOATING
C2132 out_p.n220 vss 4.56fF $ **FLOATING
C2133 out_p.n221 vss 4.56fF $ **FLOATING
C2134 out_p.n222 vss 4.56fF $ **FLOATING
C2135 out_p.n223 vss 4.56fF $ **FLOATING
C2136 out_p.n224 vss 4.56fF $ **FLOATING
C2137 out_p.n225 vss 4.56fF $ **FLOATING
C2138 out_p.n226 vss 4.56fF $ **FLOATING
C2139 out_p.n227 vss 4.56fF $ **FLOATING
C2140 out_p.n228 vss 4.56fF $ **FLOATING
C2141 out_p.n229 vss 4.56fF $ **FLOATING
C2142 out_p.n230 vss 4.56fF $ **FLOATING
C2143 out_p.n231 vss 4.56fF $ **FLOATING
C2144 out_p.n232 vss 4.56fF $ **FLOATING
C2145 out_p.n233 vss 4.56fF $ **FLOATING
C2146 out_p.n234 vss 4.56fF $ **FLOATING
C2147 out_p.n235 vss 4.27fF $ **FLOATING
C2148 out_p.n236 vss 4.37fF $ **FLOATING
C2149 out_p.n237 vss 4.53fF $ **FLOATING
C2150 out_p.n238 vss 4.53fF $ **FLOATING
C2151 out_p.n239 vss 4.26fF $ **FLOATING
C2152 out_p.n240 vss 4.40fF $ **FLOATING
C2153 out_p.n241 vss 4.56fF $ **FLOATING
C2154 out_p.n242 vss 4.56fF $ **FLOATING
C2155 out_p.n243 vss 4.56fF $ **FLOATING
C2156 out_p.n244 vss 4.56fF $ **FLOATING
C2157 out_p.n245 vss 4.56fF $ **FLOATING
C2158 out_p.n246 vss 4.56fF $ **FLOATING
C2159 out_p.n247 vss 4.56fF $ **FLOATING
C2160 out_p.n248 vss 4.56fF $ **FLOATING
C2161 out_p.n249 vss 4.56fF $ **FLOATING
C2162 out_p.n250 vss 4.56fF $ **FLOATING
C2163 out_p.n251 vss 4.56fF $ **FLOATING
C2164 out_p.n252 vss 4.56fF $ **FLOATING
C2165 out_p.n253 vss 4.56fF $ **FLOATING
C2166 out_p.n254 vss 4.56fF $ **FLOATING
C2167 out_p.n255 vss 4.56fF $ **FLOATING
C2168 out_p.n256 vss 4.56fF $ **FLOATING
C2169 out_p.n257 vss 4.56fF $ **FLOATING
C2170 out_p.n258 vss 4.56fF $ **FLOATING
C2171 out_p.n259 vss 4.27fF $ **FLOATING
C2172 out_p.n260 vss 4.37fF $ **FLOATING
C2173 out_p.n261 vss 4.53fF $ **FLOATING
C2174 out_p.n262 vss 4.53fF $ **FLOATING
C2175 out_p.n263 vss 4.26fF $ **FLOATING
C2176 out_p.n264 vss 4.40fF $ **FLOATING
C2177 out_p.n265 vss 4.56fF $ **FLOATING
C2178 out_p.n266 vss 4.56fF $ **FLOATING
C2179 out_p.n267 vss 4.56fF $ **FLOATING
C2180 out_p.n268 vss 4.56fF $ **FLOATING
C2181 out_p.n269 vss 4.56fF $ **FLOATING
C2182 out_p.n270 vss 4.56fF $ **FLOATING
C2183 out_p.n271 vss 4.56fF $ **FLOATING
C2184 out_p.n272 vss 4.56fF $ **FLOATING
C2185 out_p.n273 vss 4.56fF $ **FLOATING
C2186 out_p.n274 vss 4.56fF $ **FLOATING
C2187 out_p.n275 vss 4.56fF $ **FLOATING
C2188 out_p.n276 vss 4.56fF $ **FLOATING
C2189 out_p.n277 vss 4.56fF $ **FLOATING
C2190 out_p.n278 vss 4.56fF $ **FLOATING
C2191 out_p.n279 vss 4.56fF $ **FLOATING
C2192 out_p.n280 vss 4.56fF $ **FLOATING
C2193 out_p.n281 vss 4.56fF $ **FLOATING
C2194 out_p.n282 vss 4.56fF $ **FLOATING
C2195 out_p.n283 vss 4.27fF $ **FLOATING
C2196 out_p.n284 vss 4.37fF $ **FLOATING
C2197 out_p.n285 vss 4.53fF $ **FLOATING
C2198 out_p.n286 vss 4.53fF $ **FLOATING
C2199 out_p.n287 vss 4.26fF $ **FLOATING
C2200 out_p.n288 vss 4.40fF $ **FLOATING
C2201 out_p.n289 vss 4.56fF $ **FLOATING
C2202 out_p.n290 vss 4.56fF $ **FLOATING
C2203 out_p.n291 vss 4.56fF $ **FLOATING
C2204 out_p.n292 vss 4.56fF $ **FLOATING
C2205 out_p.n293 vss 4.56fF $ **FLOATING
C2206 out_p.n294 vss 4.56fF $ **FLOATING
C2207 out_p.n295 vss 4.56fF $ **FLOATING
C2208 out_p.n296 vss 4.56fF $ **FLOATING
C2209 out_p.n297 vss 4.56fF $ **FLOATING
C2210 out_p.n298 vss 4.56fF $ **FLOATING
C2211 out_p.n299 vss 4.56fF $ **FLOATING
C2212 out_p.n300 vss 4.56fF $ **FLOATING
C2213 out_p.n301 vss 4.56fF $ **FLOATING
C2214 out_p.n302 vss 4.56fF $ **FLOATING
C2215 out_p.n303 vss 4.56fF $ **FLOATING
C2216 out_p.n304 vss 4.56fF $ **FLOATING
C2217 out_p.n305 vss 4.56fF $ **FLOATING
C2218 out_p.n306 vss 4.56fF $ **FLOATING
C2219 out_p.n307 vss 4.27fF $ **FLOATING
C2220 out_p.n308 vss 4.37fF $ **FLOATING
C2221 out_p.n309 vss 4.53fF $ **FLOATING
C2222 out_p.n310 vss 4.53fF $ **FLOATING
C2223 out_p.n311 vss 4.26fF $ **FLOATING
C2224 out_p.n312 vss 4.40fF $ **FLOATING
C2225 out_p.n313 vss 4.56fF $ **FLOATING
C2226 out_p.n314 vss 4.56fF $ **FLOATING
C2227 out_p.n315 vss 4.56fF $ **FLOATING
C2228 out_p.n316 vss 4.56fF $ **FLOATING
C2229 out_p.n317 vss 4.56fF $ **FLOATING
C2230 out_p.n318 vss 4.56fF $ **FLOATING
C2231 out_p.n319 vss 4.56fF $ **FLOATING
C2232 out_p.n320 vss 4.56fF $ **FLOATING
C2233 out_p.n321 vss 4.56fF $ **FLOATING
C2234 out_p.n322 vss 4.56fF $ **FLOATING
C2235 out_p.n323 vss 4.56fF $ **FLOATING
C2236 out_p.n324 vss 4.56fF $ **FLOATING
C2237 out_p.n325 vss 4.56fF $ **FLOATING
C2238 out_p.n326 vss 4.56fF $ **FLOATING
C2239 out_p.n327 vss 4.56fF $ **FLOATING
C2240 out_p.n328 vss 4.56fF $ **FLOATING
C2241 out_p.n329 vss 4.56fF $ **FLOATING
C2242 out_p.n330 vss 4.56fF $ **FLOATING
C2243 out_p.n331 vss 4.27fF $ **FLOATING
C2244 out_p.n332 vss 4.37fF $ **FLOATING
C2245 out_p.n333 vss 4.53fF $ **FLOATING
C2246 out_p.n334 vss 4.53fF $ **FLOATING
C2247 out_p.n335 vss 4.26fF $ **FLOATING
C2248 out_p.n336 vss 4.40fF $ **FLOATING
C2249 out_p.n337 vss 4.56fF $ **FLOATING
C2250 out_p.n338 vss 4.56fF $ **FLOATING
C2251 out_p.n339 vss 4.56fF $ **FLOATING
C2252 out_p.n340 vss 4.56fF $ **FLOATING
C2253 out_p.n341 vss 4.56fF $ **FLOATING
C2254 out_p.n342 vss 4.56fF $ **FLOATING
C2255 out_p.n343 vss 4.56fF $ **FLOATING
C2256 out_p.n344 vss 4.56fF $ **FLOATING
C2257 out_p.n345 vss 4.56fF $ **FLOATING
C2258 out_p.n346 vss 4.56fF $ **FLOATING
C2259 out_p.n347 vss 4.56fF $ **FLOATING
C2260 out_p.n348 vss 4.56fF $ **FLOATING
C2261 out_p.n349 vss 4.56fF $ **FLOATING
C2262 out_p.n350 vss 4.56fF $ **FLOATING
C2263 out_p.n351 vss 4.56fF $ **FLOATING
C2264 out_p.n352 vss 4.56fF $ **FLOATING
C2265 out_p.n353 vss 4.56fF $ **FLOATING
C2266 out_p.n354 vss 4.56fF $ **FLOATING
C2267 out_p.n355 vss 4.27fF $ **FLOATING
C2268 out_p.n356 vss 4.37fF $ **FLOATING
C2269 out_p.n357 vss 4.53fF $ **FLOATING
C2270 out_p.n358 vss 4.53fF $ **FLOATING
C2271 out_p.n359 vss 4.26fF $ **FLOATING
C2272 out_p.n360 vss 4.40fF $ **FLOATING
C2273 out_p.n361 vss 4.56fF $ **FLOATING
C2274 out_p.n362 vss 4.56fF $ **FLOATING
C2275 out_p.n363 vss 4.56fF $ **FLOATING
C2276 out_p.n364 vss 4.56fF $ **FLOATING
C2277 out_p.n365 vss 4.56fF $ **FLOATING
C2278 out_p.n366 vss 4.56fF $ **FLOATING
C2279 out_p.n367 vss 4.56fF $ **FLOATING
C2280 out_p.n368 vss 4.56fF $ **FLOATING
C2281 out_p.n369 vss 4.56fF $ **FLOATING
C2282 out_p.n370 vss 4.56fF $ **FLOATING
C2283 out_p.n371 vss 4.56fF $ **FLOATING
C2284 out_p.n372 vss 4.56fF $ **FLOATING
C2285 out_p.n373 vss 4.56fF $ **FLOATING
C2286 out_p.n374 vss 4.56fF $ **FLOATING
C2287 out_p.n375 vss 4.56fF $ **FLOATING
C2288 out_p.n376 vss 4.56fF $ **FLOATING
C2289 out_p.n377 vss 4.56fF $ **FLOATING
C2290 out_p.n378 vss 4.56fF $ **FLOATING
C2291 out_p.n379 vss 4.27fF $ **FLOATING
C2292 out_p.n380 vss 4.37fF $ **FLOATING
C2293 out_p.n381 vss 4.53fF $ **FLOATING
C2294 out_p.n382 vss 4.53fF $ **FLOATING
C2295 out_p.n383 vss 4.26fF $ **FLOATING
C2296 out_p.n384 vss 4.40fF $ **FLOATING
C2297 out_p.n385 vss 4.56fF $ **FLOATING
C2298 out_p.n386 vss 4.56fF $ **FLOATING
C2299 out_p.n387 vss 4.56fF $ **FLOATING
C2300 out_p.n388 vss 4.56fF $ **FLOATING
C2301 out_p.n389 vss 4.56fF $ **FLOATING
C2302 out_p.n390 vss 4.56fF $ **FLOATING
C2303 out_p.n391 vss 4.56fF $ **FLOATING
C2304 out_p.n392 vss 4.56fF $ **FLOATING
C2305 out_p.n393 vss 4.56fF $ **FLOATING
C2306 out_p.n394 vss 4.56fF $ **FLOATING
C2307 out_p.n395 vss 4.56fF $ **FLOATING
C2308 out_p.n396 vss 4.56fF $ **FLOATING
C2309 out_p.n397 vss 4.56fF $ **FLOATING
C2310 out_p.n398 vss 4.56fF $ **FLOATING
C2311 out_p.n399 vss 4.56fF $ **FLOATING
C2312 out_p.n400 vss 4.56fF $ **FLOATING
C2313 out_p.n401 vss 4.56fF $ **FLOATING
C2314 out_p.n402 vss 4.56fF $ **FLOATING
C2315 out_p.n403 vss 4.27fF $ **FLOATING
C2316 out_p.n404 vss 4.37fF $ **FLOATING
C2317 out_p.n405 vss 4.53fF $ **FLOATING
C2318 out_p.n406 vss 4.53fF $ **FLOATING
C2319 out_p.n407 vss 4.26fF $ **FLOATING
C2320 out_p.n408 vss 4.40fF $ **FLOATING
C2321 out_p.n409 vss 4.56fF $ **FLOATING
C2322 out_p.n410 vss 4.56fF $ **FLOATING
C2323 out_p.n411 vss 4.56fF $ **FLOATING
C2324 out_p.n412 vss 4.56fF $ **FLOATING
C2325 out_p.n413 vss 4.56fF $ **FLOATING
C2326 out_p.n414 vss 4.56fF $ **FLOATING
C2327 out_p.n415 vss 4.56fF $ **FLOATING
C2328 out_p.n416 vss 4.56fF $ **FLOATING
C2329 out_p.n417 vss 4.56fF $ **FLOATING
C2330 out_p.n418 vss 4.56fF $ **FLOATING
C2331 out_p.n419 vss 4.56fF $ **FLOATING
C2332 out_p.n420 vss 4.56fF $ **FLOATING
C2333 out_p.n421 vss 4.56fF $ **FLOATING
C2334 out_p.n422 vss 4.56fF $ **FLOATING
C2335 out_p.n423 vss 4.56fF $ **FLOATING
C2336 out_p.n424 vss 4.56fF $ **FLOATING
C2337 out_p.n425 vss 4.56fF $ **FLOATING
C2338 out_p.n426 vss 4.56fF $ **FLOATING
C2339 out_p.n427 vss 4.27fF $ **FLOATING
C2340 out_p.n428 vss 4.37fF $ **FLOATING
C2341 out_p.n429 vss 4.53fF $ **FLOATING
C2342 out_p.n430 vss 4.53fF $ **FLOATING
C2343 out_p.n431 vss 4.26fF $ **FLOATING
C2344 out_p.n432 vss 4.40fF $ **FLOATING
C2345 out_p.n433 vss 4.56fF $ **FLOATING
C2346 out_p.n434 vss 4.56fF $ **FLOATING
C2347 out_p.n435 vss 4.56fF $ **FLOATING
C2348 out_p.n436 vss 4.56fF $ **FLOATING
C2349 out_p.n437 vss 4.56fF $ **FLOATING
C2350 out_p.n438 vss 4.56fF $ **FLOATING
C2351 out_p.n439 vss 4.56fF $ **FLOATING
C2352 out_p.n440 vss 4.56fF $ **FLOATING
C2353 out_p.n441 vss 4.56fF $ **FLOATING
C2354 out_p.n442 vss 4.56fF $ **FLOATING
C2355 out_p.n443 vss 4.56fF $ **FLOATING
C2356 out_p.n444 vss 4.56fF $ **FLOATING
C2357 out_p.n445 vss 4.56fF $ **FLOATING
C2358 out_p.n446 vss 4.56fF $ **FLOATING
C2359 out_p.n447 vss 4.56fF $ **FLOATING
C2360 out_p.n448 vss 4.56fF $ **FLOATING
C2361 out_p.n449 vss 4.56fF $ **FLOATING
C2362 out_p.n450 vss 4.56fF $ **FLOATING
C2363 out_p.n451 vss 4.27fF $ **FLOATING
C2364 out_p.n452 vss 4.37fF $ **FLOATING
C2365 out_p.n453 vss 4.53fF $ **FLOATING
C2366 out_p.n454 vss 4.53fF $ **FLOATING
C2367 out_p.n455 vss 4.26fF $ **FLOATING
C2368 out_p.n456 vss 4.40fF $ **FLOATING
C2369 out_p.n457 vss 4.56fF $ **FLOATING
C2370 out_p.n458 vss 4.56fF $ **FLOATING
C2371 out_p.n459 vss 4.56fF $ **FLOATING
C2372 out_p.n460 vss 4.56fF $ **FLOATING
C2373 out_p.n461 vss 4.56fF $ **FLOATING
C2374 out_p.n462 vss 4.56fF $ **FLOATING
C2375 out_p.n463 vss 4.56fF $ **FLOATING
C2376 out_p.n464 vss 4.56fF $ **FLOATING
C2377 out_p.n465 vss 4.56fF $ **FLOATING
C2378 out_p.n466 vss 4.56fF $ **FLOATING
C2379 out_p.n467 vss 4.56fF $ **FLOATING
C2380 out_p.n468 vss 4.56fF $ **FLOATING
C2381 out_p.n469 vss 4.56fF $ **FLOATING
C2382 out_p.n470 vss 4.56fF $ **FLOATING
C2383 out_p.n471 vss 4.56fF $ **FLOATING
C2384 out_p.n472 vss 4.56fF $ **FLOATING
C2385 out_p.n473 vss 4.56fF $ **FLOATING
C2386 out_p.n474 vss 4.56fF $ **FLOATING
C2387 out_p.n475 vss 4.27fF $ **FLOATING
C2388 out_p.n476 vss 4.37fF $ **FLOATING
C2389 out_p.n477 vss 4.53fF $ **FLOATING
C2390 out_p.n478 vss 4.53fF $ **FLOATING
C2391 out_p.n479 vss 4.26fF $ **FLOATING
C2392 out_p.n480 vss 4.40fF $ **FLOATING
C2393 out_p.n481 vss 4.56fF $ **FLOATING
C2394 out_p.n482 vss 4.56fF $ **FLOATING
C2395 out_p.n483 vss 4.56fF $ **FLOATING
C2396 out_p.n484 vss 4.56fF $ **FLOATING
C2397 out_p.n485 vss 4.56fF $ **FLOATING
C2398 out_p.n486 vss 4.56fF $ **FLOATING
C2399 out_p.n487 vss 4.56fF $ **FLOATING
C2400 out_p.n488 vss 4.56fF $ **FLOATING
C2401 out_p.n489 vss 4.56fF $ **FLOATING
C2402 out_p.n490 vss 4.56fF $ **FLOATING
C2403 out_p.n491 vss 4.56fF $ **FLOATING
C2404 out_p.n492 vss 4.56fF $ **FLOATING
C2405 out_p.n493 vss 4.56fF $ **FLOATING
C2406 out_p.n494 vss 4.56fF $ **FLOATING
C2407 out_p.n495 vss 4.56fF $ **FLOATING
C2408 out_p.n496 vss 4.56fF $ **FLOATING
C2409 out_p.n497 vss 4.56fF $ **FLOATING
C2410 out_p.n498 vss 4.56fF $ **FLOATING
C2411 out_p.n499 vss 4.27fF $ **FLOATING
C2412 out_p.n500 vss 4.37fF $ **FLOATING
C2413 out_p.n501 vss 4.53fF $ **FLOATING
C2414 out_p.n502 vss 4.53fF $ **FLOATING
C2415 out_p.n503 vss 4.26fF $ **FLOATING
C2416 out_p.n504 vss 4.40fF $ **FLOATING
C2417 out_p.n505 vss 4.56fF $ **FLOATING
C2418 out_p.n506 vss 4.56fF $ **FLOATING
C2419 out_p.n507 vss 4.56fF $ **FLOATING
C2420 out_p.n508 vss 4.56fF $ **FLOATING
C2421 out_p.n509 vss 4.56fF $ **FLOATING
C2422 out_p.n510 vss 4.56fF $ **FLOATING
C2423 out_p.n511 vss 4.56fF $ **FLOATING
C2424 out_p.n512 vss 4.56fF $ **FLOATING
C2425 out_p.n513 vss 4.56fF $ **FLOATING
C2426 out_p.n514 vss 4.56fF $ **FLOATING
C2427 out_p.n515 vss 4.56fF $ **FLOATING
C2428 out_p.n516 vss 4.56fF $ **FLOATING
C2429 out_p.n517 vss 4.56fF $ **FLOATING
C2430 out_p.n518 vss 4.56fF $ **FLOATING
C2431 out_p.n519 vss 4.56fF $ **FLOATING
C2432 out_p.n520 vss 4.56fF $ **FLOATING
C2433 out_p.n521 vss 4.56fF $ **FLOATING
C2434 out_p.n522 vss 4.56fF $ **FLOATING
C2435 out_p.n523 vss 4.27fF $ **FLOATING
C2436 out_p.n524 vss 4.37fF $ **FLOATING
C2437 out_p.n525 vss 4.53fF $ **FLOATING
C2438 out_p.n526 vss 4.53fF $ **FLOATING
C2439 out_p.n527 vss 4.26fF $ **FLOATING
C2440 out_p.n528 vss 4.40fF $ **FLOATING
C2441 out_p.n529 vss 4.56fF $ **FLOATING
C2442 out_p.n530 vss 4.56fF $ **FLOATING
C2443 out_p.n531 vss 4.56fF $ **FLOATING
C2444 out_p.n532 vss 4.56fF $ **FLOATING
C2445 out_p.n533 vss 4.56fF $ **FLOATING
C2446 out_p.n534 vss 4.56fF $ **FLOATING
C2447 out_p.n535 vss 4.56fF $ **FLOATING
C2448 out_p.n536 vss 4.56fF $ **FLOATING
C2449 out_p.n537 vss 4.56fF $ **FLOATING
C2450 out_p.n538 vss 4.56fF $ **FLOATING
C2451 out_p.n539 vss 4.56fF $ **FLOATING
C2452 out_p.n540 vss 4.56fF $ **FLOATING
C2453 out_p.n541 vss 4.56fF $ **FLOATING
C2454 out_p.n542 vss 4.56fF $ **FLOATING
C2455 out_p.n543 vss 4.56fF $ **FLOATING
C2456 out_p.n544 vss 4.56fF $ **FLOATING
C2457 out_p.n545 vss 4.56fF $ **FLOATING
C2458 out_p.n546 vss 4.56fF $ **FLOATING
C2459 out_p.n547 vss 4.27fF $ **FLOATING
C2460 out_p.n548 vss 4.37fF $ **FLOATING
C2461 out_p.n549 vss 4.53fF $ **FLOATING
C2462 out_p.n550 vss 4.53fF $ **FLOATING
C2463 out_p.n551 vss 4.26fF $ **FLOATING
C2464 out_p.n552 vss 4.40fF $ **FLOATING
C2465 out_p.n553 vss 4.56fF $ **FLOATING
C2466 out_p.n554 vss 4.56fF $ **FLOATING
C2467 out_p.n555 vss 4.56fF $ **FLOATING
C2468 out_p.n556 vss 4.56fF $ **FLOATING
C2469 out_p.n557 vss 4.56fF $ **FLOATING
C2470 out_p.n558 vss 4.56fF $ **FLOATING
C2471 out_p.n559 vss 4.56fF $ **FLOATING
C2472 out_p.n560 vss 4.56fF $ **FLOATING
C2473 out_p.n561 vss 4.56fF $ **FLOATING
C2474 out_p.n562 vss 4.56fF $ **FLOATING
C2475 out_p.n563 vss 4.56fF $ **FLOATING
C2476 out_p.n564 vss 4.56fF $ **FLOATING
C2477 out_p.n565 vss 4.56fF $ **FLOATING
C2478 out_p.n566 vss 4.56fF $ **FLOATING
C2479 out_p.n567 vss 4.56fF $ **FLOATING
C2480 out_p.n568 vss 4.56fF $ **FLOATING
C2481 out_p.n569 vss 4.56fF $ **FLOATING
C2482 out_p.n570 vss 4.56fF $ **FLOATING
C2483 out_p.n571 vss 4.27fF $ **FLOATING
C2484 out_p.n572 vss 4.37fF $ **FLOATING
C2485 out_p.n573 vss 4.53fF $ **FLOATING
C2486 out_p.n574 vss 4.53fF $ **FLOATING
C2487 out_p.n575 vss 4.26fF $ **FLOATING
C2488 out_p.n576 vss 4.40fF $ **FLOATING
C2489 out_p.n577 vss 4.56fF $ **FLOATING
C2490 out_p.n578 vss 4.56fF $ **FLOATING
C2491 out_p.n579 vss 4.56fF $ **FLOATING
C2492 out_p.n580 vss 4.56fF $ **FLOATING
C2493 out_p.n581 vss 4.56fF $ **FLOATING
C2494 out_p.n582 vss 4.56fF $ **FLOATING
C2495 out_p.n583 vss 4.56fF $ **FLOATING
C2496 out_p.n584 vss 4.56fF $ **FLOATING
C2497 out_p.n585 vss 4.56fF $ **FLOATING
C2498 out_p.n586 vss 4.56fF $ **FLOATING
C2499 out_p.n587 vss 4.56fF $ **FLOATING
C2500 out_p.n588 vss 4.56fF $ **FLOATING
C2501 out_p.n589 vss 4.56fF $ **FLOATING
C2502 out_p.n590 vss 4.56fF $ **FLOATING
C2503 out_p.n591 vss 4.56fF $ **FLOATING
C2504 out_p.n592 vss 4.56fF $ **FLOATING
C2505 out_p.n593 vss 4.56fF $ **FLOATING
C2506 out_p.n594 vss 4.56fF $ **FLOATING
C2507 out_p.n595 vss 4.27fF $ **FLOATING
C2508 out_p.n596 vss 4.37fF $ **FLOATING
C2509 out_p.n597 vss 4.53fF $ **FLOATING
C2510 out_p.n598 vss 4.53fF $ **FLOATING
C2511 out_p.n599 vss 4.26fF $ **FLOATING
C2512 out_p.n600 vss 4.40fF $ **FLOATING
C2513 out_p.n601 vss 4.56fF $ **FLOATING
C2514 out_p.n602 vss 4.56fF $ **FLOATING
C2515 out_p.n603 vss 4.56fF $ **FLOATING
C2516 out_p.n604 vss 4.56fF $ **FLOATING
C2517 out_p.n605 vss 4.56fF $ **FLOATING
C2518 out_p.n606 vss 4.56fF $ **FLOATING
C2519 out_p.n607 vss 4.56fF $ **FLOATING
C2520 out_p.n608 vss 4.56fF $ **FLOATING
C2521 out_p.n609 vss 4.56fF $ **FLOATING
C2522 out_p.n610 vss 4.56fF $ **FLOATING
C2523 out_p.n611 vss 4.56fF $ **FLOATING
C2524 out_p.n612 vss 4.56fF $ **FLOATING
C2525 out_p.n613 vss 4.56fF $ **FLOATING
C2526 out_p.n614 vss 4.56fF $ **FLOATING
C2527 out_p.n615 vss 4.56fF $ **FLOATING
C2528 out_p.n616 vss 4.56fF $ **FLOATING
C2529 out_p.n617 vss 4.56fF $ **FLOATING
C2530 out_p.n618 vss 4.56fF $ **FLOATING
C2531 out_p.n619 vss 4.27fF $ **FLOATING
C2532 out_p.n620 vss 4.37fF $ **FLOATING
C2533 out_p.n621 vss 4.53fF $ **FLOATING
C2534 out_p.n622 vss 4.53fF $ **FLOATING
C2535 out_p.n623 vss 4.26fF $ **FLOATING
C2536 out_p.n624 vss 4.40fF $ **FLOATING
C2537 out_p.n625 vss 4.56fF $ **FLOATING
C2538 out_p.n626 vss 4.56fF $ **FLOATING
C2539 out_p.n627 vss 4.56fF $ **FLOATING
C2540 out_p.n628 vss 4.56fF $ **FLOATING
C2541 out_p.n629 vss 4.56fF $ **FLOATING
C2542 out_p.n630 vss 4.56fF $ **FLOATING
C2543 out_p.n631 vss 4.56fF $ **FLOATING
C2544 out_p.n632 vss 4.56fF $ **FLOATING
C2545 out_p.n633 vss 4.56fF $ **FLOATING
C2546 out_p.n634 vss 4.56fF $ **FLOATING
C2547 out_p.n635 vss 4.56fF $ **FLOATING
C2548 out_p.n636 vss 4.56fF $ **FLOATING
C2549 out_p.n637 vss 4.56fF $ **FLOATING
C2550 out_p.n638 vss 4.56fF $ **FLOATING
C2551 out_p.n639 vss 4.56fF $ **FLOATING
C2552 out_p.n640 vss 4.56fF $ **FLOATING
C2553 out_p.n641 vss 4.56fF $ **FLOATING
C2554 out_p.n642 vss 4.56fF $ **FLOATING
C2555 out_p.n643 vss 4.27fF $ **FLOATING
C2556 out_p.n644 vss 4.37fF $ **FLOATING
C2557 out_p.n645 vss 4.53fF $ **FLOATING
C2558 out_p.n646 vss 4.53fF $ **FLOATING
C2559 out_p.n647 vss 4.26fF $ **FLOATING
C2560 out_p.n648 vss 4.40fF $ **FLOATING
C2561 out_p.n649 vss 4.56fF $ **FLOATING
C2562 out_p.n650 vss 4.56fF $ **FLOATING
C2563 out_p.n651 vss 4.56fF $ **FLOATING
C2564 out_p.n652 vss 4.56fF $ **FLOATING
C2565 out_p.n653 vss 4.56fF $ **FLOATING
C2566 out_p.n654 vss 4.56fF $ **FLOATING
C2567 out_p.n655 vss 4.56fF $ **FLOATING
C2568 out_p.n656 vss 4.56fF $ **FLOATING
C2569 out_p.n657 vss 4.56fF $ **FLOATING
C2570 out_p.n658 vss 4.56fF $ **FLOATING
C2571 out_p.n659 vss 4.56fF $ **FLOATING
C2572 out_p.n660 vss 4.56fF $ **FLOATING
C2573 out_p.n661 vss 4.56fF $ **FLOATING
C2574 out_p.n662 vss 4.56fF $ **FLOATING
C2575 out_p.n663 vss 4.56fF $ **FLOATING
C2576 out_p.n664 vss 4.56fF $ **FLOATING
C2577 out_p.n665 vss 4.56fF $ **FLOATING
C2578 out_p.n666 vss 4.56fF $ **FLOATING
C2579 out_p.n667 vss 4.27fF $ **FLOATING
C2580 out_p.n668 vss 4.37fF $ **FLOATING
C2581 out_p.n669 vss 4.53fF $ **FLOATING
C2582 out_p.n670 vss 4.53fF $ **FLOATING
C2583 out_p.n671 vss 4.26fF $ **FLOATING
C2584 out_p.n672 vss 4.40fF $ **FLOATING
C2585 out_p.n673 vss 4.56fF $ **FLOATING
C2586 out_p.n674 vss 4.56fF $ **FLOATING
C2587 out_p.n675 vss 4.56fF $ **FLOATING
C2588 out_p.n676 vss 4.56fF $ **FLOATING
C2589 out_p.n677 vss 4.56fF $ **FLOATING
C2590 out_p.n678 vss 4.56fF $ **FLOATING
C2591 out_p.n679 vss 4.56fF $ **FLOATING
C2592 out_p.n680 vss 4.56fF $ **FLOATING
C2593 out_p.n681 vss 4.56fF $ **FLOATING
C2594 out_p.n682 vss 4.56fF $ **FLOATING
C2595 out_p.n683 vss 4.56fF $ **FLOATING
C2596 out_p.n684 vss 4.56fF $ **FLOATING
C2597 out_p.n685 vss 4.56fF $ **FLOATING
C2598 out_p.n686 vss 4.56fF $ **FLOATING
C2599 out_p.n687 vss 4.56fF $ **FLOATING
C2600 out_p.n688 vss 4.56fF $ **FLOATING
C2601 out_p.n689 vss 4.56fF $ **FLOATING
C2602 out_p.n690 vss 4.56fF $ **FLOATING
C2603 out_p.n691 vss 4.27fF $ **FLOATING
C2604 out_p.n692 vss 4.37fF $ **FLOATING
C2605 out_p.n693 vss 4.53fF $ **FLOATING
C2606 out_p.n694 vss 4.53fF $ **FLOATING
C2607 out_p.n695 vss 4.26fF $ **FLOATING
C2608 out_p.n696 vss 4.40fF $ **FLOATING
C2609 out_p.n697 vss 4.56fF $ **FLOATING
C2610 out_p.n698 vss 4.56fF $ **FLOATING
C2611 out_p.n699 vss 4.56fF $ **FLOATING
C2612 out_p.n700 vss 4.56fF $ **FLOATING
C2613 out_p.n701 vss 4.56fF $ **FLOATING
C2614 out_p.n702 vss 4.56fF $ **FLOATING
C2615 out_p.n703 vss 4.56fF $ **FLOATING
C2616 out_p.n704 vss 4.56fF $ **FLOATING
C2617 out_p.n705 vss 4.56fF $ **FLOATING
C2618 out_p.n706 vss 4.56fF $ **FLOATING
C2619 out_p.n707 vss 4.56fF $ **FLOATING
C2620 out_p.n708 vss 4.56fF $ **FLOATING
C2621 out_p.n709 vss 4.56fF $ **FLOATING
C2622 out_p.n710 vss 4.56fF $ **FLOATING
C2623 out_p.n711 vss 4.56fF $ **FLOATING
C2624 out_p.n712 vss 4.56fF $ **FLOATING
C2625 out_p.n713 vss 4.56fF $ **FLOATING
C2626 out_p.n714 vss 4.56fF $ **FLOATING
C2627 out_p.n715 vss 4.27fF $ **FLOATING
C2628 out_p.n716 vss 4.37fF $ **FLOATING
C2629 out_p.n717 vss 4.53fF $ **FLOATING
C2630 out_p.n718 vss 4.53fF $ **FLOATING
C2631 out_p.n719 vss 4.26fF $ **FLOATING
C2632 out_p.n720 vss 4.40fF $ **FLOATING
C2633 out_p.n721 vss 4.56fF $ **FLOATING
C2634 out_p.n722 vss 4.56fF $ **FLOATING
C2635 out_p.n723 vss 4.56fF $ **FLOATING
C2636 out_p.n724 vss 4.56fF $ **FLOATING
C2637 out_p.n725 vss 4.56fF $ **FLOATING
C2638 out_p.n726 vss 4.56fF $ **FLOATING
C2639 out_p.n727 vss 4.56fF $ **FLOATING
C2640 out_p.n728 vss 4.56fF $ **FLOATING
C2641 out_p.n729 vss 4.56fF $ **FLOATING
C2642 out_p.n730 vss 4.56fF $ **FLOATING
C2643 out_p.n731 vss 4.56fF $ **FLOATING
C2644 out_p.n732 vss 4.56fF $ **FLOATING
C2645 out_p.n733 vss 4.56fF $ **FLOATING
C2646 out_p.n734 vss 4.56fF $ **FLOATING
C2647 out_p.n735 vss 4.56fF $ **FLOATING
C2648 out_p.n736 vss 4.56fF $ **FLOATING
C2649 out_p.n737 vss 4.56fF $ **FLOATING
C2650 out_p.n738 vss 4.56fF $ **FLOATING
C2651 out_p.n739 vss 4.27fF $ **FLOATING
C2652 out_p.n740 vss 4.37fF $ **FLOATING
C2653 out_p.n741 vss 4.53fF $ **FLOATING
C2654 out_p.n742 vss 4.53fF $ **FLOATING
C2655 out_p.n743 vss 4.26fF $ **FLOATING
C2656 out_p.n744 vss 4.34fF $ **FLOATING
C2657 out_p.n745 vss 4.22fF $ **FLOATING
C2658 out_p.n747 vss 4.04fF $ **FLOATING
C2659 out_p.n748 vss 4.23fF $ **FLOATING
C2660 out_p.n749 vss 4.40fF $ **FLOATING
C2661 out_p.n750 vss 4.56fF $ **FLOATING
C2662 out_p.n751 vss 4.56fF $ **FLOATING
C2663 out_p.n752 vss 4.56fF $ **FLOATING
C2664 out_p.n753 vss 4.56fF $ **FLOATING
C2665 out_p.n754 vss 4.56fF $ **FLOATING
C2666 out_p.n755 vss 4.56fF $ **FLOATING
C2667 out_p.n756 vss 4.56fF $ **FLOATING
C2668 out_p.n757 vss 4.56fF $ **FLOATING
C2669 out_p.n758 vss 4.56fF $ **FLOATING
C2670 out_p.n759 vss 4.56fF $ **FLOATING
C2671 out_p.n760 vss 4.56fF $ **FLOATING
C2672 out_p.n761 vss 4.56fF $ **FLOATING
C2673 out_p.n762 vss 4.56fF $ **FLOATING
C2674 out_p.n763 vss 4.56fF $ **FLOATING
C2675 out_p.n764 vss 4.56fF $ **FLOATING
C2676 out_p.n765 vss 4.56fF $ **FLOATING
C2677 out_p.n766 vss 4.56fF $ **FLOATING
C2678 out_p.n767 vss 4.56fF $ **FLOATING
C2679 out_p.n768 vss 4.27fF $ **FLOATING
C2680 out_p.n769 vss 59.03fF $ **FLOATING
C2681 out_p.n770 vss 85.73fF $ **FLOATING
C2682 out_p.n771 vss 85.93fF $ **FLOATING
C2683 out_p.n772 vss 85.93fF $ **FLOATING
C2684 out_p.n773 vss 85.93fF $ **FLOATING
C2685 out_p.n774 vss 85.93fF $ **FLOATING
C2686 out_p.n775 vss 85.93fF $ **FLOATING
C2687 out_p.n776 vss 85.93fF $ **FLOATING
C2688 out_p.n777 vss 85.93fF $ **FLOATING
C2689 out_p.n778 vss 85.93fF $ **FLOATING
C2690 out_p.n779 vss 85.93fF $ **FLOATING
C2691 out_p.n780 vss 85.93fF $ **FLOATING
C2692 out_p.n781 vss 85.93fF $ **FLOATING
C2693 out_p.n782 vss 85.93fF $ **FLOATING
C2694 out_p.n783 vss 85.93fF $ **FLOATING
C2695 out_p.n784 vss 85.93fF $ **FLOATING
C2696 out_p.n785 vss 85.93fF $ **FLOATING
C2697 out_p.n786 vss 85.93fF $ **FLOATING
C2698 out_p.n787 vss 85.93fF $ **FLOATING
C2699 out_p.n788 vss 85.93fF $ **FLOATING
C2700 out_p.n789 vss 85.93fF $ **FLOATING
C2701 out_p.n790 vss 85.93fF $ **FLOATING
C2702 out_p.n791 vss 85.93fF $ **FLOATING
C2703 out_p.n792 vss 85.93fF $ **FLOATING
C2704 out_p.n793 vss 85.93fF $ **FLOATING
C2705 out_p.n794 vss 85.93fF $ **FLOATING
C2706 out_p.n795 vss 85.93fF $ **FLOATING
C2707 out_p.n796 vss 85.93fF $ **FLOATING
C2708 out_p.n797 vss 85.93fF $ **FLOATING
C2709 out_p.n798 vss 85.93fF $ **FLOATING
C2710 out_p.n799 vss 85.93fF $ **FLOATING
C2711 out_p.n800 vss 85.93fF $ **FLOATING
C2712 out_p.n801 vss 4.37fF $ **FLOATING
C2713 out_p.n802 vss 4.53fF $ **FLOATING
C2714 out_p.n803 vss 4.53fF $ **FLOATING
C2715 out_p.n804 vss 4.26fF $ **FLOATING
C2716 out_p.n805 vss 4.40fF $ **FLOATING
C2717 out_p.n806 vss 4.56fF $ **FLOATING
C2718 out_p.n807 vss 4.56fF $ **FLOATING
C2719 out_p.n808 vss 4.56fF $ **FLOATING
C2720 out_p.n809 vss 4.56fF $ **FLOATING
C2721 out_p.n810 vss 4.56fF $ **FLOATING
C2722 out_p.n811 vss 4.56fF $ **FLOATING
C2723 out_p.n812 vss 4.56fF $ **FLOATING
C2724 out_p.n813 vss 4.56fF $ **FLOATING
C2725 out_p.n814 vss 4.56fF $ **FLOATING
C2726 out_p.n815 vss 4.56fF $ **FLOATING
C2727 out_p.n816 vss 4.56fF $ **FLOATING
C2728 out_p.n817 vss 4.56fF $ **FLOATING
C2729 out_p.n818 vss 4.56fF $ **FLOATING
C2730 out_p.n819 vss 4.56fF $ **FLOATING
C2731 out_p.n820 vss 4.56fF $ **FLOATING
C2732 out_p.n821 vss 4.56fF $ **FLOATING
C2733 out_p.n822 vss 4.56fF $ **FLOATING
C2734 out_p.n823 vss 4.56fF $ **FLOATING
C2735 out_p.n824 vss 4.27fF $ **FLOATING
C2736 out_p.n825 vss 4.40fF $ **FLOATING
C2737 out_p.n826 vss 4.56fF $ **FLOATING
C2738 out_p.n827 vss 4.56fF $ **FLOATING
C2739 out_p.n828 vss 4.56fF $ **FLOATING
C2740 out_p.n829 vss 4.56fF $ **FLOATING
C2741 out_p.n830 vss 4.56fF $ **FLOATING
C2742 out_p.n831 vss 4.56fF $ **FLOATING
C2743 out_p.n832 vss 4.56fF $ **FLOATING
C2744 out_p.n833 vss 4.56fF $ **FLOATING
C2745 out_p.n834 vss 4.56fF $ **FLOATING
C2746 out_p.n835 vss 4.56fF $ **FLOATING
C2747 out_p.n836 vss 4.56fF $ **FLOATING
C2748 out_p.n837 vss 4.56fF $ **FLOATING
C2749 out_p.n838 vss 4.56fF $ **FLOATING
C2750 out_p.n839 vss 4.56fF $ **FLOATING
C2751 out_p.n840 vss 4.56fF $ **FLOATING
C2752 out_p.n841 vss 4.56fF $ **FLOATING
C2753 out_p.n842 vss 4.56fF $ **FLOATING
C2754 out_p.n843 vss 4.56fF $ **FLOATING
C2755 out_p.n844 vss 4.27fF $ **FLOATING
C2756 out_p.n845 vss 4.37fF $ **FLOATING
C2757 out_p.n846 vss 4.53fF $ **FLOATING
C2758 out_p.n847 vss 4.53fF $ **FLOATING
C2759 out_p.n848 vss 4.26fF $ **FLOATING
C2760 out_p.n849 vss 4.40fF $ **FLOATING
C2761 out_p.n850 vss 4.56fF $ **FLOATING
C2762 out_p.n851 vss 4.56fF $ **FLOATING
C2763 out_p.n852 vss 4.56fF $ **FLOATING
C2764 out_p.n853 vss 4.56fF $ **FLOATING
C2765 out_p.n854 vss 4.56fF $ **FLOATING
C2766 out_p.n855 vss 4.56fF $ **FLOATING
C2767 out_p.n856 vss 4.56fF $ **FLOATING
C2768 out_p.n857 vss 4.56fF $ **FLOATING
C2769 out_p.n858 vss 4.56fF $ **FLOATING
C2770 out_p.n859 vss 4.56fF $ **FLOATING
C2771 out_p.n860 vss 4.56fF $ **FLOATING
C2772 out_p.n861 vss 4.56fF $ **FLOATING
C2773 out_p.n862 vss 4.56fF $ **FLOATING
C2774 out_p.n863 vss 4.56fF $ **FLOATING
C2775 out_p.n864 vss 4.56fF $ **FLOATING
C2776 out_p.n865 vss 4.56fF $ **FLOATING
C2777 out_p.n866 vss 4.56fF $ **FLOATING
C2778 out_p.n867 vss 4.56fF $ **FLOATING
C2779 out_p.n868 vss 4.27fF $ **FLOATING
C2780 out_p.n869 vss 4.37fF $ **FLOATING
C2781 out_p.n870 vss 4.53fF $ **FLOATING
C2782 out_p.n871 vss 4.53fF $ **FLOATING
C2783 out_p.n872 vss 4.26fF $ **FLOATING
C2784 out_p.n873 vss 4.40fF $ **FLOATING
C2785 out_p.n874 vss 4.56fF $ **FLOATING
C2786 out_p.n875 vss 4.56fF $ **FLOATING
C2787 out_p.n876 vss 4.56fF $ **FLOATING
C2788 out_p.n877 vss 4.56fF $ **FLOATING
C2789 out_p.n878 vss 4.56fF $ **FLOATING
C2790 out_p.n879 vss 4.56fF $ **FLOATING
C2791 out_p.n880 vss 4.56fF $ **FLOATING
C2792 out_p.n881 vss 4.56fF $ **FLOATING
C2793 out_p.n882 vss 4.56fF $ **FLOATING
C2794 out_p.n883 vss 4.56fF $ **FLOATING
C2795 out_p.n884 vss 4.56fF $ **FLOATING
C2796 out_p.n885 vss 4.56fF $ **FLOATING
C2797 out_p.n886 vss 4.56fF $ **FLOATING
C2798 out_p.n887 vss 4.56fF $ **FLOATING
C2799 out_p.n888 vss 4.56fF $ **FLOATING
C2800 out_p.n889 vss 4.56fF $ **FLOATING
C2801 out_p.n890 vss 4.56fF $ **FLOATING
C2802 out_p.n891 vss 4.56fF $ **FLOATING
C2803 out_p.n892 vss 4.27fF $ **FLOATING
C2804 out_p.n893 vss 4.37fF $ **FLOATING
C2805 out_p.n894 vss 4.53fF $ **FLOATING
C2806 out_p.n895 vss 4.53fF $ **FLOATING
C2807 out_p.n896 vss 4.26fF $ **FLOATING
C2808 out_p.n897 vss 4.40fF $ **FLOATING
C2809 out_p.n898 vss 4.56fF $ **FLOATING
C2810 out_p.n899 vss 4.56fF $ **FLOATING
C2811 out_p.n900 vss 4.56fF $ **FLOATING
C2812 out_p.n901 vss 4.56fF $ **FLOATING
C2813 out_p.n902 vss 4.56fF $ **FLOATING
C2814 out_p.n903 vss 4.56fF $ **FLOATING
C2815 out_p.n904 vss 4.56fF $ **FLOATING
C2816 out_p.n905 vss 4.56fF $ **FLOATING
C2817 out_p.n906 vss 4.56fF $ **FLOATING
C2818 out_p.n907 vss 4.56fF $ **FLOATING
C2819 out_p.n908 vss 4.56fF $ **FLOATING
C2820 out_p.n909 vss 4.56fF $ **FLOATING
C2821 out_p.n910 vss 4.56fF $ **FLOATING
C2822 out_p.n911 vss 4.56fF $ **FLOATING
C2823 out_p.n912 vss 4.56fF $ **FLOATING
C2824 out_p.n913 vss 4.56fF $ **FLOATING
C2825 out_p.n914 vss 4.56fF $ **FLOATING
C2826 out_p.n915 vss 4.56fF $ **FLOATING
C2827 out_p.n916 vss 4.27fF $ **FLOATING
C2828 out_p.n917 vss 4.37fF $ **FLOATING
C2829 out_p.n918 vss 4.53fF $ **FLOATING
C2830 out_p.n919 vss 4.53fF $ **FLOATING
C2831 out_p.n920 vss 4.26fF $ **FLOATING
C2832 out_p.n921 vss 4.40fF $ **FLOATING
C2833 out_p.n922 vss 4.56fF $ **FLOATING
C2834 out_p.n923 vss 4.56fF $ **FLOATING
C2835 out_p.n924 vss 4.56fF $ **FLOATING
C2836 out_p.n925 vss 4.56fF $ **FLOATING
C2837 out_p.n926 vss 4.56fF $ **FLOATING
C2838 out_p.n927 vss 4.56fF $ **FLOATING
C2839 out_p.n928 vss 4.56fF $ **FLOATING
C2840 out_p.n929 vss 4.56fF $ **FLOATING
C2841 out_p.n930 vss 4.56fF $ **FLOATING
C2842 out_p.n931 vss 4.56fF $ **FLOATING
C2843 out_p.n932 vss 4.56fF $ **FLOATING
C2844 out_p.n933 vss 4.56fF $ **FLOATING
C2845 out_p.n934 vss 4.56fF $ **FLOATING
C2846 out_p.n935 vss 4.56fF $ **FLOATING
C2847 out_p.n936 vss 4.56fF $ **FLOATING
C2848 out_p.n937 vss 4.56fF $ **FLOATING
C2849 out_p.n938 vss 4.56fF $ **FLOATING
C2850 out_p.n939 vss 4.56fF $ **FLOATING
C2851 out_p.n940 vss 4.27fF $ **FLOATING
C2852 out_p.n941 vss 4.37fF $ **FLOATING
C2853 out_p.n942 vss 4.53fF $ **FLOATING
C2854 out_p.n943 vss 4.53fF $ **FLOATING
C2855 out_p.n944 vss 4.26fF $ **FLOATING
C2856 out_p.n945 vss 4.40fF $ **FLOATING
C2857 out_p.n946 vss 4.56fF $ **FLOATING
C2858 out_p.n947 vss 4.56fF $ **FLOATING
C2859 out_p.n948 vss 4.56fF $ **FLOATING
C2860 out_p.n949 vss 4.56fF $ **FLOATING
C2861 out_p.n950 vss 4.56fF $ **FLOATING
C2862 out_p.n951 vss 4.56fF $ **FLOATING
C2863 out_p.n952 vss 4.56fF $ **FLOATING
C2864 out_p.n953 vss 4.56fF $ **FLOATING
C2865 out_p.n954 vss 4.56fF $ **FLOATING
C2866 out_p.n955 vss 4.56fF $ **FLOATING
C2867 out_p.n956 vss 4.56fF $ **FLOATING
C2868 out_p.n957 vss 4.56fF $ **FLOATING
C2869 out_p.n958 vss 4.56fF $ **FLOATING
C2870 out_p.n959 vss 4.56fF $ **FLOATING
C2871 out_p.n960 vss 4.56fF $ **FLOATING
C2872 out_p.n961 vss 4.56fF $ **FLOATING
C2873 out_p.n962 vss 4.56fF $ **FLOATING
C2874 out_p.n963 vss 4.56fF $ **FLOATING
C2875 out_p.n964 vss 4.27fF $ **FLOATING
C2876 out_p.n965 vss 4.37fF $ **FLOATING
C2877 out_p.n966 vss 4.53fF $ **FLOATING
C2878 out_p.n967 vss 4.53fF $ **FLOATING
C2879 out_p.n968 vss 4.26fF $ **FLOATING
C2880 out_p.n969 vss 4.40fF $ **FLOATING
C2881 out_p.n970 vss 4.56fF $ **FLOATING
C2882 out_p.n971 vss 4.56fF $ **FLOATING
C2883 out_p.n972 vss 4.56fF $ **FLOATING
C2884 out_p.n973 vss 4.56fF $ **FLOATING
C2885 out_p.n974 vss 4.56fF $ **FLOATING
C2886 out_p.n975 vss 4.56fF $ **FLOATING
C2887 out_p.n976 vss 4.56fF $ **FLOATING
C2888 out_p.n977 vss 4.56fF $ **FLOATING
C2889 out_p.n978 vss 4.56fF $ **FLOATING
C2890 out_p.n979 vss 4.56fF $ **FLOATING
C2891 out_p.n980 vss 4.56fF $ **FLOATING
C2892 out_p.n981 vss 4.56fF $ **FLOATING
C2893 out_p.n982 vss 4.56fF $ **FLOATING
C2894 out_p.n983 vss 4.56fF $ **FLOATING
C2895 out_p.n984 vss 4.56fF $ **FLOATING
C2896 out_p.n985 vss 4.56fF $ **FLOATING
C2897 out_p.n986 vss 4.56fF $ **FLOATING
C2898 out_p.n987 vss 4.56fF $ **FLOATING
C2899 out_p.n988 vss 4.27fF $ **FLOATING
C2900 out_p.n989 vss 4.37fF $ **FLOATING
C2901 out_p.n990 vss 4.53fF $ **FLOATING
C2902 out_p.n991 vss 4.53fF $ **FLOATING
C2903 out_p.n992 vss 4.26fF $ **FLOATING
C2904 out_p.n993 vss 4.40fF $ **FLOATING
C2905 out_p.n994 vss 4.56fF $ **FLOATING
C2906 out_p.n995 vss 4.56fF $ **FLOATING
C2907 out_p.n996 vss 4.56fF $ **FLOATING
C2908 out_p.n997 vss 4.56fF $ **FLOATING
C2909 out_p.n998 vss 4.56fF $ **FLOATING
C2910 out_p.n999 vss 4.56fF $ **FLOATING
C2911 out_p.n1000 vss 4.56fF $ **FLOATING
C2912 out_p.n1001 vss 4.56fF $ **FLOATING
C2913 out_p.n1002 vss 4.56fF $ **FLOATING
C2914 out_p.n1003 vss 4.56fF $ **FLOATING
C2915 out_p.n1004 vss 4.56fF $ **FLOATING
C2916 out_p.n1005 vss 4.56fF $ **FLOATING
C2917 out_p.n1006 vss 4.56fF $ **FLOATING
C2918 out_p.n1007 vss 4.56fF $ **FLOATING
C2919 out_p.n1008 vss 4.56fF $ **FLOATING
C2920 out_p.n1009 vss 4.56fF $ **FLOATING
C2921 out_p.n1010 vss 4.56fF $ **FLOATING
C2922 out_p.n1011 vss 4.56fF $ **FLOATING
C2923 out_p.n1012 vss 4.27fF $ **FLOATING
C2924 out_p.n1013 vss 4.37fF $ **FLOATING
C2925 out_p.n1014 vss 4.53fF $ **FLOATING
C2926 out_p.n1015 vss 4.53fF $ **FLOATING
C2927 out_p.n1016 vss 4.26fF $ **FLOATING
C2928 out_p.n1017 vss 4.40fF $ **FLOATING
C2929 out_p.n1018 vss 4.56fF $ **FLOATING
C2930 out_p.n1019 vss 4.56fF $ **FLOATING
C2931 out_p.n1020 vss 4.56fF $ **FLOATING
C2932 out_p.n1021 vss 4.56fF $ **FLOATING
C2933 out_p.n1022 vss 4.56fF $ **FLOATING
C2934 out_p.n1023 vss 4.56fF $ **FLOATING
C2935 out_p.n1024 vss 4.56fF $ **FLOATING
C2936 out_p.n1025 vss 4.56fF $ **FLOATING
C2937 out_p.n1026 vss 4.56fF $ **FLOATING
C2938 out_p.n1027 vss 4.56fF $ **FLOATING
C2939 out_p.n1028 vss 4.56fF $ **FLOATING
C2940 out_p.n1029 vss 4.56fF $ **FLOATING
C2941 out_p.n1030 vss 4.56fF $ **FLOATING
C2942 out_p.n1031 vss 4.56fF $ **FLOATING
C2943 out_p.n1032 vss 4.56fF $ **FLOATING
C2944 out_p.n1033 vss 4.56fF $ **FLOATING
C2945 out_p.n1034 vss 4.56fF $ **FLOATING
C2946 out_p.n1035 vss 4.56fF $ **FLOATING
C2947 out_p.n1036 vss 4.27fF $ **FLOATING
C2948 out_p.n1037 vss 4.37fF $ **FLOATING
C2949 out_p.n1038 vss 4.53fF $ **FLOATING
C2950 out_p.n1039 vss 4.53fF $ **FLOATING
C2951 out_p.n1040 vss 4.26fF $ **FLOATING
C2952 out_p.n1041 vss 4.40fF $ **FLOATING
C2953 out_p.n1042 vss 4.56fF $ **FLOATING
C2954 out_p.n1043 vss 4.56fF $ **FLOATING
C2955 out_p.n1044 vss 4.56fF $ **FLOATING
C2956 out_p.n1045 vss 4.56fF $ **FLOATING
C2957 out_p.n1046 vss 4.56fF $ **FLOATING
C2958 out_p.n1047 vss 4.56fF $ **FLOATING
C2959 out_p.n1048 vss 4.56fF $ **FLOATING
C2960 out_p.n1049 vss 4.56fF $ **FLOATING
C2961 out_p.n1050 vss 4.56fF $ **FLOATING
C2962 out_p.n1051 vss 4.56fF $ **FLOATING
C2963 out_p.n1052 vss 4.56fF $ **FLOATING
C2964 out_p.n1053 vss 4.56fF $ **FLOATING
C2965 out_p.n1054 vss 4.56fF $ **FLOATING
C2966 out_p.n1055 vss 4.56fF $ **FLOATING
C2967 out_p.n1056 vss 4.56fF $ **FLOATING
C2968 out_p.n1057 vss 4.56fF $ **FLOATING
C2969 out_p.n1058 vss 4.56fF $ **FLOATING
C2970 out_p.n1059 vss 4.56fF $ **FLOATING
C2971 out_p.n1060 vss 4.27fF $ **FLOATING
C2972 out_p.n1061 vss 4.37fF $ **FLOATING
C2973 out_p.n1062 vss 4.53fF $ **FLOATING
C2974 out_p.n1063 vss 4.53fF $ **FLOATING
C2975 out_p.n1064 vss 4.26fF $ **FLOATING
C2976 out_p.n1065 vss 4.40fF $ **FLOATING
C2977 out_p.n1066 vss 4.56fF $ **FLOATING
C2978 out_p.n1067 vss 4.56fF $ **FLOATING
C2979 out_p.n1068 vss 4.56fF $ **FLOATING
C2980 out_p.n1069 vss 4.56fF $ **FLOATING
C2981 out_p.n1070 vss 4.56fF $ **FLOATING
C2982 out_p.n1071 vss 4.56fF $ **FLOATING
C2983 out_p.n1072 vss 4.56fF $ **FLOATING
C2984 out_p.n1073 vss 4.56fF $ **FLOATING
C2985 out_p.n1074 vss 4.56fF $ **FLOATING
C2986 out_p.n1075 vss 4.56fF $ **FLOATING
C2987 out_p.n1076 vss 4.56fF $ **FLOATING
C2988 out_p.n1077 vss 4.56fF $ **FLOATING
C2989 out_p.n1078 vss 4.56fF $ **FLOATING
C2990 out_p.n1079 vss 4.56fF $ **FLOATING
C2991 out_p.n1080 vss 4.56fF $ **FLOATING
C2992 out_p.n1081 vss 4.56fF $ **FLOATING
C2993 out_p.n1082 vss 4.56fF $ **FLOATING
C2994 out_p.n1083 vss 4.56fF $ **FLOATING
C2995 out_p.n1084 vss 4.27fF $ **FLOATING
C2996 out_p.n1085 vss 4.37fF $ **FLOATING
C2997 out_p.n1086 vss 4.53fF $ **FLOATING
C2998 out_p.n1087 vss 4.53fF $ **FLOATING
C2999 out_p.n1088 vss 4.26fF $ **FLOATING
C3000 out_p.n1089 vss 4.40fF $ **FLOATING
C3001 out_p.n1090 vss 4.56fF $ **FLOATING
C3002 out_p.n1091 vss 4.56fF $ **FLOATING
C3003 out_p.n1092 vss 4.56fF $ **FLOATING
C3004 out_p.n1093 vss 4.56fF $ **FLOATING
C3005 out_p.n1094 vss 4.56fF $ **FLOATING
C3006 out_p.n1095 vss 4.56fF $ **FLOATING
C3007 out_p.n1096 vss 4.56fF $ **FLOATING
C3008 out_p.n1097 vss 4.56fF $ **FLOATING
C3009 out_p.n1098 vss 4.56fF $ **FLOATING
C3010 out_p.n1099 vss 4.56fF $ **FLOATING
C3011 out_p.n1100 vss 4.56fF $ **FLOATING
C3012 out_p.n1101 vss 4.56fF $ **FLOATING
C3013 out_p.n1102 vss 4.56fF $ **FLOATING
C3014 out_p.n1103 vss 4.56fF $ **FLOATING
C3015 out_p.n1104 vss 4.56fF $ **FLOATING
C3016 out_p.n1105 vss 4.56fF $ **FLOATING
C3017 out_p.n1106 vss 4.56fF $ **FLOATING
C3018 out_p.n1107 vss 4.56fF $ **FLOATING
C3019 out_p.n1108 vss 4.27fF $ **FLOATING
C3020 out_p.n1109 vss 4.37fF $ **FLOATING
C3021 out_p.n1110 vss 4.53fF $ **FLOATING
C3022 out_p.n1111 vss 4.53fF $ **FLOATING
C3023 out_p.n1112 vss 4.26fF $ **FLOATING
C3024 out_p.n1113 vss 4.40fF $ **FLOATING
C3025 out_p.n1114 vss 4.56fF $ **FLOATING
C3026 out_p.n1115 vss 4.56fF $ **FLOATING
C3027 out_p.n1116 vss 4.56fF $ **FLOATING
C3028 out_p.n1117 vss 4.56fF $ **FLOATING
C3029 out_p.n1118 vss 4.56fF $ **FLOATING
C3030 out_p.n1119 vss 4.56fF $ **FLOATING
C3031 out_p.n1120 vss 4.56fF $ **FLOATING
C3032 out_p.n1121 vss 4.56fF $ **FLOATING
C3033 out_p.n1122 vss 4.56fF $ **FLOATING
C3034 out_p.n1123 vss 4.56fF $ **FLOATING
C3035 out_p.n1124 vss 4.56fF $ **FLOATING
C3036 out_p.n1125 vss 4.56fF $ **FLOATING
C3037 out_p.n1126 vss 4.56fF $ **FLOATING
C3038 out_p.n1127 vss 4.56fF $ **FLOATING
C3039 out_p.n1128 vss 4.56fF $ **FLOATING
C3040 out_p.n1129 vss 4.56fF $ **FLOATING
C3041 out_p.n1130 vss 4.56fF $ **FLOATING
C3042 out_p.n1131 vss 4.56fF $ **FLOATING
C3043 out_p.n1132 vss 4.27fF $ **FLOATING
C3044 out_p.n1133 vss 4.37fF $ **FLOATING
C3045 out_p.n1134 vss 4.53fF $ **FLOATING
C3046 out_p.n1135 vss 4.53fF $ **FLOATING
C3047 out_p.n1136 vss 4.26fF $ **FLOATING
C3048 out_p.n1137 vss 4.40fF $ **FLOATING
C3049 out_p.n1138 vss 4.56fF $ **FLOATING
C3050 out_p.n1139 vss 4.56fF $ **FLOATING
C3051 out_p.n1140 vss 4.56fF $ **FLOATING
C3052 out_p.n1141 vss 4.56fF $ **FLOATING
C3053 out_p.n1142 vss 4.56fF $ **FLOATING
C3054 out_p.n1143 vss 4.56fF $ **FLOATING
C3055 out_p.n1144 vss 4.56fF $ **FLOATING
C3056 out_p.n1145 vss 4.56fF $ **FLOATING
C3057 out_p.n1146 vss 4.56fF $ **FLOATING
C3058 out_p.n1147 vss 4.56fF $ **FLOATING
C3059 out_p.n1148 vss 4.56fF $ **FLOATING
C3060 out_p.n1149 vss 4.56fF $ **FLOATING
C3061 out_p.n1150 vss 4.56fF $ **FLOATING
C3062 out_p.n1151 vss 4.56fF $ **FLOATING
C3063 out_p.n1152 vss 4.56fF $ **FLOATING
C3064 out_p.n1153 vss 4.56fF $ **FLOATING
C3065 out_p.n1154 vss 4.56fF $ **FLOATING
C3066 out_p.n1155 vss 4.56fF $ **FLOATING
C3067 out_p.n1156 vss 4.27fF $ **FLOATING
C3068 out_p.n1157 vss 4.37fF $ **FLOATING
C3069 out_p.n1158 vss 4.53fF $ **FLOATING
C3070 out_p.n1159 vss 4.53fF $ **FLOATING
C3071 out_p.n1160 vss 4.26fF $ **FLOATING
C3072 out_p.n1161 vss 4.40fF $ **FLOATING
C3073 out_p.n1162 vss 4.56fF $ **FLOATING
C3074 out_p.n1163 vss 4.56fF $ **FLOATING
C3075 out_p.n1164 vss 4.56fF $ **FLOATING
C3076 out_p.n1165 vss 4.56fF $ **FLOATING
C3077 out_p.n1166 vss 4.56fF $ **FLOATING
C3078 out_p.n1167 vss 4.56fF $ **FLOATING
C3079 out_p.n1168 vss 4.56fF $ **FLOATING
C3080 out_p.n1169 vss 4.56fF $ **FLOATING
C3081 out_p.n1170 vss 4.56fF $ **FLOATING
C3082 out_p.n1171 vss 4.56fF $ **FLOATING
C3083 out_p.n1172 vss 4.56fF $ **FLOATING
C3084 out_p.n1173 vss 4.56fF $ **FLOATING
C3085 out_p.n1174 vss 4.56fF $ **FLOATING
C3086 out_p.n1175 vss 4.56fF $ **FLOATING
C3087 out_p.n1176 vss 4.56fF $ **FLOATING
C3088 out_p.n1177 vss 4.56fF $ **FLOATING
C3089 out_p.n1178 vss 4.56fF $ **FLOATING
C3090 out_p.n1179 vss 4.56fF $ **FLOATING
C3091 out_p.n1180 vss 4.27fF $ **FLOATING
C3092 out_p.n1181 vss 4.37fF $ **FLOATING
C3093 out_p.n1182 vss 4.53fF $ **FLOATING
C3094 out_p.n1183 vss 4.53fF $ **FLOATING
C3095 out_p.n1184 vss 4.26fF $ **FLOATING
C3096 out_p.n1185 vss 4.40fF $ **FLOATING
C3097 out_p.n1186 vss 4.56fF $ **FLOATING
C3098 out_p.n1187 vss 4.56fF $ **FLOATING
C3099 out_p.n1188 vss 4.56fF $ **FLOATING
C3100 out_p.n1189 vss 4.56fF $ **FLOATING
C3101 out_p.n1190 vss 4.56fF $ **FLOATING
C3102 out_p.n1191 vss 4.56fF $ **FLOATING
C3103 out_p.n1192 vss 4.56fF $ **FLOATING
C3104 out_p.n1193 vss 4.56fF $ **FLOATING
C3105 out_p.n1194 vss 4.56fF $ **FLOATING
C3106 out_p.n1195 vss 4.56fF $ **FLOATING
C3107 out_p.n1196 vss 4.56fF $ **FLOATING
C3108 out_p.n1197 vss 4.56fF $ **FLOATING
C3109 out_p.n1198 vss 4.56fF $ **FLOATING
C3110 out_p.n1199 vss 4.56fF $ **FLOATING
C3111 out_p.n1200 vss 4.56fF $ **FLOATING
C3112 out_p.n1201 vss 4.56fF $ **FLOATING
C3113 out_p.n1202 vss 4.56fF $ **FLOATING
C3114 out_p.n1203 vss 4.56fF $ **FLOATING
C3115 out_p.n1204 vss 4.27fF $ **FLOATING
C3116 out_p.n1205 vss 4.37fF $ **FLOATING
C3117 out_p.n1206 vss 4.53fF $ **FLOATING
C3118 out_p.n1207 vss 4.53fF $ **FLOATING
C3119 out_p.n1208 vss 4.26fF $ **FLOATING
C3120 out_p.n1209 vss 4.40fF $ **FLOATING
C3121 out_p.n1210 vss 4.56fF $ **FLOATING
C3122 out_p.n1211 vss 4.56fF $ **FLOATING
C3123 out_p.n1212 vss 4.56fF $ **FLOATING
C3124 out_p.n1213 vss 4.56fF $ **FLOATING
C3125 out_p.n1214 vss 4.56fF $ **FLOATING
C3126 out_p.n1215 vss 4.56fF $ **FLOATING
C3127 out_p.n1216 vss 4.56fF $ **FLOATING
C3128 out_p.n1217 vss 4.56fF $ **FLOATING
C3129 out_p.n1218 vss 4.56fF $ **FLOATING
C3130 out_p.n1219 vss 4.56fF $ **FLOATING
C3131 out_p.n1220 vss 4.56fF $ **FLOATING
C3132 out_p.n1221 vss 4.56fF $ **FLOATING
C3133 out_p.n1222 vss 4.56fF $ **FLOATING
C3134 out_p.n1223 vss 4.56fF $ **FLOATING
C3135 out_p.n1224 vss 4.56fF $ **FLOATING
C3136 out_p.n1225 vss 4.56fF $ **FLOATING
C3137 out_p.n1226 vss 4.56fF $ **FLOATING
C3138 out_p.n1227 vss 4.56fF $ **FLOATING
C3139 out_p.n1228 vss 4.27fF $ **FLOATING
C3140 out_p.n1229 vss 4.37fF $ **FLOATING
C3141 out_p.n1230 vss 4.53fF $ **FLOATING
C3142 out_p.n1231 vss 4.53fF $ **FLOATING
C3143 out_p.n1232 vss 4.26fF $ **FLOATING
C3144 out_p.n1233 vss 4.40fF $ **FLOATING
C3145 out_p.n1234 vss 4.56fF $ **FLOATING
C3146 out_p.n1235 vss 4.56fF $ **FLOATING
C3147 out_p.n1236 vss 4.56fF $ **FLOATING
C3148 out_p.n1237 vss 4.56fF $ **FLOATING
C3149 out_p.n1238 vss 4.56fF $ **FLOATING
C3150 out_p.n1239 vss 4.56fF $ **FLOATING
C3151 out_p.n1240 vss 4.56fF $ **FLOATING
C3152 out_p.n1241 vss 4.56fF $ **FLOATING
C3153 out_p.n1242 vss 4.56fF $ **FLOATING
C3154 out_p.n1243 vss 4.56fF $ **FLOATING
C3155 out_p.n1244 vss 4.56fF $ **FLOATING
C3156 out_p.n1245 vss 4.56fF $ **FLOATING
C3157 out_p.n1246 vss 4.56fF $ **FLOATING
C3158 out_p.n1247 vss 4.56fF $ **FLOATING
C3159 out_p.n1248 vss 4.56fF $ **FLOATING
C3160 out_p.n1249 vss 4.56fF $ **FLOATING
C3161 out_p.n1250 vss 4.56fF $ **FLOATING
C3162 out_p.n1251 vss 4.56fF $ **FLOATING
C3163 out_p.n1252 vss 4.27fF $ **FLOATING
C3164 out_p.n1253 vss 4.37fF $ **FLOATING
C3165 out_p.n1254 vss 4.53fF $ **FLOATING
C3166 out_p.n1255 vss 4.53fF $ **FLOATING
C3167 out_p.n1256 vss 4.26fF $ **FLOATING
C3168 out_p.n1257 vss 4.40fF $ **FLOATING
C3169 out_p.n1258 vss 4.56fF $ **FLOATING
C3170 out_p.n1259 vss 4.56fF $ **FLOATING
C3171 out_p.n1260 vss 4.56fF $ **FLOATING
C3172 out_p.n1261 vss 4.56fF $ **FLOATING
C3173 out_p.n1262 vss 4.56fF $ **FLOATING
C3174 out_p.n1263 vss 4.56fF $ **FLOATING
C3175 out_p.n1264 vss 4.56fF $ **FLOATING
C3176 out_p.n1265 vss 4.56fF $ **FLOATING
C3177 out_p.n1266 vss 4.56fF $ **FLOATING
C3178 out_p.n1267 vss 4.56fF $ **FLOATING
C3179 out_p.n1268 vss 4.56fF $ **FLOATING
C3180 out_p.n1269 vss 4.56fF $ **FLOATING
C3181 out_p.n1270 vss 4.56fF $ **FLOATING
C3182 out_p.n1271 vss 4.56fF $ **FLOATING
C3183 out_p.n1272 vss 4.56fF $ **FLOATING
C3184 out_p.n1273 vss 4.56fF $ **FLOATING
C3185 out_p.n1274 vss 4.56fF $ **FLOATING
C3186 out_p.n1275 vss 4.56fF $ **FLOATING
C3187 out_p.n1276 vss 4.27fF $ **FLOATING
C3188 out_p.n1277 vss 4.37fF $ **FLOATING
C3189 out_p.n1278 vss 4.53fF $ **FLOATING
C3190 out_p.n1279 vss 4.53fF $ **FLOATING
C3191 out_p.n1280 vss 4.26fF $ **FLOATING
C3192 out_p.n1281 vss 4.40fF $ **FLOATING
C3193 out_p.n1282 vss 4.56fF $ **FLOATING
C3194 out_p.n1283 vss 4.56fF $ **FLOATING
C3195 out_p.n1284 vss 4.56fF $ **FLOATING
C3196 out_p.n1285 vss 4.56fF $ **FLOATING
C3197 out_p.n1286 vss 4.56fF $ **FLOATING
C3198 out_p.n1287 vss 4.56fF $ **FLOATING
C3199 out_p.n1288 vss 4.56fF $ **FLOATING
C3200 out_p.n1289 vss 4.56fF $ **FLOATING
C3201 out_p.n1290 vss 4.56fF $ **FLOATING
C3202 out_p.n1291 vss 4.56fF $ **FLOATING
C3203 out_p.n1292 vss 4.56fF $ **FLOATING
C3204 out_p.n1293 vss 4.56fF $ **FLOATING
C3205 out_p.n1294 vss 4.56fF $ **FLOATING
C3206 out_p.n1295 vss 4.56fF $ **FLOATING
C3207 out_p.n1296 vss 4.56fF $ **FLOATING
C3208 out_p.n1297 vss 4.56fF $ **FLOATING
C3209 out_p.n1298 vss 4.56fF $ **FLOATING
C3210 out_p.n1299 vss 4.56fF $ **FLOATING
C3211 out_p.n1300 vss 4.27fF $ **FLOATING
C3212 out_p.n1301 vss 4.37fF $ **FLOATING
C3213 out_p.n1302 vss 4.53fF $ **FLOATING
C3214 out_p.n1303 vss 4.53fF $ **FLOATING
C3215 out_p.n1304 vss 4.26fF $ **FLOATING
C3216 out_p.n1305 vss 4.40fF $ **FLOATING
C3217 out_p.n1306 vss 4.56fF $ **FLOATING
C3218 out_p.n1307 vss 4.56fF $ **FLOATING
C3219 out_p.n1308 vss 4.56fF $ **FLOATING
C3220 out_p.n1309 vss 4.56fF $ **FLOATING
C3221 out_p.n1310 vss 4.56fF $ **FLOATING
C3222 out_p.n1311 vss 4.56fF $ **FLOATING
C3223 out_p.n1312 vss 4.56fF $ **FLOATING
C3224 out_p.n1313 vss 4.56fF $ **FLOATING
C3225 out_p.n1314 vss 4.56fF $ **FLOATING
C3226 out_p.n1315 vss 4.56fF $ **FLOATING
C3227 out_p.n1316 vss 4.56fF $ **FLOATING
C3228 out_p.n1317 vss 4.56fF $ **FLOATING
C3229 out_p.n1318 vss 4.56fF $ **FLOATING
C3230 out_p.n1319 vss 4.56fF $ **FLOATING
C3231 out_p.n1320 vss 4.56fF $ **FLOATING
C3232 out_p.n1321 vss 4.56fF $ **FLOATING
C3233 out_p.n1322 vss 4.56fF $ **FLOATING
C3234 out_p.n1323 vss 4.56fF $ **FLOATING
C3235 out_p.n1324 vss 4.27fF $ **FLOATING
C3236 out_p.n1325 vss 4.37fF $ **FLOATING
C3237 out_p.n1326 vss 4.53fF $ **FLOATING
C3238 out_p.n1327 vss 4.53fF $ **FLOATING
C3239 out_p.n1328 vss 4.26fF $ **FLOATING
C3240 out_p.n1329 vss 4.40fF $ **FLOATING
C3241 out_p.n1330 vss 4.56fF $ **FLOATING
C3242 out_p.n1331 vss 4.56fF $ **FLOATING
C3243 out_p.n1332 vss 4.56fF $ **FLOATING
C3244 out_p.n1333 vss 4.56fF $ **FLOATING
C3245 out_p.n1334 vss 4.56fF $ **FLOATING
C3246 out_p.n1335 vss 4.56fF $ **FLOATING
C3247 out_p.n1336 vss 4.56fF $ **FLOATING
C3248 out_p.n1337 vss 4.56fF $ **FLOATING
C3249 out_p.n1338 vss 4.56fF $ **FLOATING
C3250 out_p.n1339 vss 4.56fF $ **FLOATING
C3251 out_p.n1340 vss 4.56fF $ **FLOATING
C3252 out_p.n1341 vss 4.56fF $ **FLOATING
C3253 out_p.n1342 vss 4.56fF $ **FLOATING
C3254 out_p.n1343 vss 4.56fF $ **FLOATING
C3255 out_p.n1344 vss 4.56fF $ **FLOATING
C3256 out_p.n1345 vss 4.56fF $ **FLOATING
C3257 out_p.n1346 vss 4.56fF $ **FLOATING
C3258 out_p.n1347 vss 4.56fF $ **FLOATING
C3259 out_p.n1348 vss 4.27fF $ **FLOATING
C3260 out_p.n1349 vss 4.37fF $ **FLOATING
C3261 out_p.n1350 vss 4.53fF $ **FLOATING
C3262 out_p.n1351 vss 4.53fF $ **FLOATING
C3263 out_p.n1352 vss 4.26fF $ **FLOATING
C3264 out_p.n1353 vss 4.40fF $ **FLOATING
C3265 out_p.n1354 vss 4.56fF $ **FLOATING
C3266 out_p.n1355 vss 4.56fF $ **FLOATING
C3267 out_p.n1356 vss 4.56fF $ **FLOATING
C3268 out_p.n1357 vss 4.56fF $ **FLOATING
C3269 out_p.n1358 vss 4.56fF $ **FLOATING
C3270 out_p.n1359 vss 4.56fF $ **FLOATING
C3271 out_p.n1360 vss 4.56fF $ **FLOATING
C3272 out_p.n1361 vss 4.56fF $ **FLOATING
C3273 out_p.n1362 vss 4.56fF $ **FLOATING
C3274 out_p.n1363 vss 4.56fF $ **FLOATING
C3275 out_p.n1364 vss 4.56fF $ **FLOATING
C3276 out_p.n1365 vss 4.56fF $ **FLOATING
C3277 out_p.n1366 vss 4.56fF $ **FLOATING
C3278 out_p.n1367 vss 4.56fF $ **FLOATING
C3279 out_p.n1368 vss 4.56fF $ **FLOATING
C3280 out_p.n1369 vss 4.56fF $ **FLOATING
C3281 out_p.n1370 vss 4.56fF $ **FLOATING
C3282 out_p.n1371 vss 4.56fF $ **FLOATING
C3283 out_p.n1372 vss 4.27fF $ **FLOATING
C3284 out_p.n1373 vss 4.37fF $ **FLOATING
C3285 out_p.n1374 vss 4.53fF $ **FLOATING
C3286 out_p.n1375 vss 4.53fF $ **FLOATING
C3287 out_p.n1376 vss 4.26fF $ **FLOATING
C3288 out_p.n1377 vss 4.40fF $ **FLOATING
C3289 out_p.n1378 vss 4.56fF $ **FLOATING
C3290 out_p.n1379 vss 4.56fF $ **FLOATING
C3291 out_p.n1380 vss 4.56fF $ **FLOATING
C3292 out_p.n1381 vss 4.56fF $ **FLOATING
C3293 out_p.n1382 vss 4.56fF $ **FLOATING
C3294 out_p.n1383 vss 4.56fF $ **FLOATING
C3295 out_p.n1384 vss 4.56fF $ **FLOATING
C3296 out_p.n1385 vss 4.56fF $ **FLOATING
C3297 out_p.n1386 vss 4.56fF $ **FLOATING
C3298 out_p.n1387 vss 4.56fF $ **FLOATING
C3299 out_p.n1388 vss 4.56fF $ **FLOATING
C3300 out_p.n1389 vss 4.56fF $ **FLOATING
C3301 out_p.n1390 vss 4.56fF $ **FLOATING
C3302 out_p.n1391 vss 4.56fF $ **FLOATING
C3303 out_p.n1392 vss 4.56fF $ **FLOATING
C3304 out_p.n1393 vss 4.56fF $ **FLOATING
C3305 out_p.n1394 vss 4.56fF $ **FLOATING
C3306 out_p.n1395 vss 4.56fF $ **FLOATING
C3307 out_p.n1396 vss 4.27fF $ **FLOATING
C3308 out_p.n1397 vss 4.37fF $ **FLOATING
C3309 out_p.n1398 vss 4.53fF $ **FLOATING
C3310 out_p.n1399 vss 4.53fF $ **FLOATING
C3311 out_p.n1400 vss 4.26fF $ **FLOATING
C3312 out_p.n1401 vss 4.40fF $ **FLOATING
C3313 out_p.n1402 vss 4.56fF $ **FLOATING
C3314 out_p.n1403 vss 4.56fF $ **FLOATING
C3315 out_p.n1404 vss 4.56fF $ **FLOATING
C3316 out_p.n1405 vss 4.56fF $ **FLOATING
C3317 out_p.n1406 vss 4.56fF $ **FLOATING
C3318 out_p.n1407 vss 4.56fF $ **FLOATING
C3319 out_p.n1408 vss 4.56fF $ **FLOATING
C3320 out_p.n1409 vss 4.56fF $ **FLOATING
C3321 out_p.n1410 vss 4.56fF $ **FLOATING
C3322 out_p.n1411 vss 4.56fF $ **FLOATING
C3323 out_p.n1412 vss 4.56fF $ **FLOATING
C3324 out_p.n1413 vss 4.56fF $ **FLOATING
C3325 out_p.n1414 vss 4.56fF $ **FLOATING
C3326 out_p.n1415 vss 4.56fF $ **FLOATING
C3327 out_p.n1416 vss 4.56fF $ **FLOATING
C3328 out_p.n1417 vss 4.56fF $ **FLOATING
C3329 out_p.n1418 vss 4.56fF $ **FLOATING
C3330 out_p.n1419 vss 4.56fF $ **FLOATING
C3331 out_p.n1420 vss 4.27fF $ **FLOATING
C3332 out_p.n1421 vss 4.37fF $ **FLOATING
C3333 out_p.n1422 vss 4.53fF $ **FLOATING
C3334 out_p.n1423 vss 4.53fF $ **FLOATING
C3335 out_p.n1424 vss 4.26fF $ **FLOATING
C3336 out_p.n1425 vss 4.40fF $ **FLOATING
C3337 out_p.n1426 vss 4.56fF $ **FLOATING
C3338 out_p.n1427 vss 4.56fF $ **FLOATING
C3339 out_p.n1428 vss 4.56fF $ **FLOATING
C3340 out_p.n1429 vss 4.56fF $ **FLOATING
C3341 out_p.n1430 vss 4.56fF $ **FLOATING
C3342 out_p.n1431 vss 4.56fF $ **FLOATING
C3343 out_p.n1432 vss 4.56fF $ **FLOATING
C3344 out_p.n1433 vss 4.56fF $ **FLOATING
C3345 out_p.n1434 vss 4.56fF $ **FLOATING
C3346 out_p.n1435 vss 4.56fF $ **FLOATING
C3347 out_p.n1436 vss 4.56fF $ **FLOATING
C3348 out_p.n1437 vss 4.56fF $ **FLOATING
C3349 out_p.n1438 vss 4.56fF $ **FLOATING
C3350 out_p.n1439 vss 4.56fF $ **FLOATING
C3351 out_p.n1440 vss 4.56fF $ **FLOATING
C3352 out_p.n1441 vss 4.56fF $ **FLOATING
C3353 out_p.n1442 vss 4.56fF $ **FLOATING
C3354 out_p.n1443 vss 4.56fF $ **FLOATING
C3355 out_p.n1444 vss 4.27fF $ **FLOATING
C3356 out_p.n1445 vss 4.37fF $ **FLOATING
C3357 out_p.n1446 vss 4.53fF $ **FLOATING
C3358 out_p.n1447 vss 4.53fF $ **FLOATING
C3359 out_p.n1448 vss 4.26fF $ **FLOATING
C3360 out_p.n1449 vss 4.40fF $ **FLOATING
C3361 out_p.n1450 vss 4.56fF $ **FLOATING
C3362 out_p.n1451 vss 4.56fF $ **FLOATING
C3363 out_p.n1452 vss 4.56fF $ **FLOATING
C3364 out_p.n1453 vss 4.56fF $ **FLOATING
C3365 out_p.n1454 vss 4.56fF $ **FLOATING
C3366 out_p.n1455 vss 4.56fF $ **FLOATING
C3367 out_p.n1456 vss 4.56fF $ **FLOATING
C3368 out_p.n1457 vss 4.56fF $ **FLOATING
C3369 out_p.n1458 vss 4.56fF $ **FLOATING
C3370 out_p.n1459 vss 4.56fF $ **FLOATING
C3371 out_p.n1460 vss 4.56fF $ **FLOATING
C3372 out_p.n1461 vss 4.56fF $ **FLOATING
C3373 out_p.n1462 vss 4.56fF $ **FLOATING
C3374 out_p.n1463 vss 4.56fF $ **FLOATING
C3375 out_p.n1464 vss 4.56fF $ **FLOATING
C3376 out_p.n1465 vss 4.56fF $ **FLOATING
C3377 out_p.n1466 vss 4.56fF $ **FLOATING
C3378 out_p.n1467 vss 4.56fF $ **FLOATING
C3379 out_p.n1468 vss 4.27fF $ **FLOATING
C3380 out_p.n1469 vss 4.37fF $ **FLOATING
C3381 out_p.n1470 vss 4.53fF $ **FLOATING
C3382 out_p.n1471 vss 4.53fF $ **FLOATING
C3383 out_p.n1472 vss 4.26fF $ **FLOATING
C3384 out_p.n1473 vss 4.40fF $ **FLOATING
C3385 out_p.n1474 vss 4.56fF $ **FLOATING
C3386 out_p.n1475 vss 4.56fF $ **FLOATING
C3387 out_p.n1476 vss 4.56fF $ **FLOATING
C3388 out_p.n1477 vss 4.56fF $ **FLOATING
C3389 out_p.n1478 vss 4.56fF $ **FLOATING
C3390 out_p.n1479 vss 4.56fF $ **FLOATING
C3391 out_p.n1480 vss 4.56fF $ **FLOATING
C3392 out_p.n1481 vss 4.56fF $ **FLOATING
C3393 out_p.n1482 vss 4.56fF $ **FLOATING
C3394 out_p.n1483 vss 4.56fF $ **FLOATING
C3395 out_p.n1484 vss 4.56fF $ **FLOATING
C3396 out_p.n1485 vss 4.56fF $ **FLOATING
C3397 out_p.n1486 vss 4.56fF $ **FLOATING
C3398 out_p.n1487 vss 4.56fF $ **FLOATING
C3399 out_p.n1488 vss 4.56fF $ **FLOATING
C3400 out_p.n1489 vss 4.56fF $ **FLOATING
C3401 out_p.n1490 vss 4.56fF $ **FLOATING
C3402 out_p.n1491 vss 4.56fF $ **FLOATING
C3403 out_p.n1492 vss 4.27fF $ **FLOATING
C3404 out_p.n1493 vss 4.37fF $ **FLOATING
C3405 out_p.n1494 vss 4.53fF $ **FLOATING
C3406 out_p.n1495 vss 4.53fF $ **FLOATING
C3407 out_p.n1496 vss 4.26fF $ **FLOATING
C3408 out_p.n1497 vss 4.40fF $ **FLOATING
C3409 out_p.n1498 vss 4.56fF $ **FLOATING
C3410 out_p.n1499 vss 4.56fF $ **FLOATING
C3411 out_p.n1500 vss 4.56fF $ **FLOATING
C3412 out_p.n1501 vss 4.56fF $ **FLOATING
C3413 out_p.n1502 vss 4.56fF $ **FLOATING
C3414 out_p.n1503 vss 4.56fF $ **FLOATING
C3415 out_p.n1504 vss 4.56fF $ **FLOATING
C3416 out_p.n1505 vss 4.56fF $ **FLOATING
C3417 out_p.n1506 vss 4.56fF $ **FLOATING
C3418 out_p.n1507 vss 4.56fF $ **FLOATING
C3419 out_p.n1508 vss 4.56fF $ **FLOATING
C3420 out_p.n1509 vss 4.56fF $ **FLOATING
C3421 out_p.n1510 vss 4.56fF $ **FLOATING
C3422 out_p.n1511 vss 4.56fF $ **FLOATING
C3423 out_p.n1512 vss 4.56fF $ **FLOATING
C3424 out_p.n1513 vss 4.56fF $ **FLOATING
C3425 out_p.n1514 vss 4.56fF $ **FLOATING
C3426 out_p.n1515 vss 4.56fF $ **FLOATING
C3427 out_p.n1516 vss 4.27fF $ **FLOATING
C3428 out_p.n1517 vss 4.37fF $ **FLOATING
C3429 out_p.n1518 vss 4.53fF $ **FLOATING
C3430 out_p.n1519 vss 4.53fF $ **FLOATING
C3431 out_p.n1520 vss 4.26fF $ **FLOATING
C3432 out_p.n1521 vss 4.40fF $ **FLOATING
C3433 out_p.n1522 vss 4.56fF $ **FLOATING
C3434 out_p.n1523 vss 4.56fF $ **FLOATING
C3435 out_p.n1524 vss 4.56fF $ **FLOATING
C3436 out_p.n1525 vss 4.56fF $ **FLOATING
C3437 out_p.n1526 vss 4.56fF $ **FLOATING
C3438 out_p.n1527 vss 4.56fF $ **FLOATING
C3439 out_p.n1528 vss 4.56fF $ **FLOATING
C3440 out_p.n1529 vss 4.56fF $ **FLOATING
C3441 out_p.n1530 vss 4.56fF $ **FLOATING
C3442 out_p.n1531 vss 4.56fF $ **FLOATING
C3443 out_p.n1532 vss 4.56fF $ **FLOATING
C3444 out_p.n1533 vss 4.56fF $ **FLOATING
C3445 out_p.n1534 vss 4.56fF $ **FLOATING
C3446 out_p.n1535 vss 4.56fF $ **FLOATING
C3447 out_p.n1536 vss 4.56fF $ **FLOATING
C3448 out_p.n1537 vss 4.56fF $ **FLOATING
C3449 out_p.n1538 vss 4.56fF $ **FLOATING
C3450 out_p.n1539 vss 4.56fF $ **FLOATING
C3451 out_p.n1540 vss 4.27fF $ **FLOATING
C3452 out_p.n1541 vss 4.37fF $ **FLOATING
C3453 out_p.n1542 vss 4.53fF $ **FLOATING
C3454 out_p.n1543 vss 4.53fF $ **FLOATING
C3455 out_p.n1544 vss 4.26fF $ **FLOATING
C3456 out_p.n1545 vss 4.40fF $ **FLOATING
C3457 out_p.n1546 vss 4.56fF $ **FLOATING
C3458 out_p.n1547 vss 4.56fF $ **FLOATING
C3459 out_p.n1548 vss 4.56fF $ **FLOATING
C3460 out_p.n1549 vss 4.56fF $ **FLOATING
C3461 out_p.n1550 vss 4.56fF $ **FLOATING
C3462 out_p.n1551 vss 4.56fF $ **FLOATING
C3463 out_p.n1552 vss 4.56fF $ **FLOATING
C3464 out_p.n1553 vss 4.56fF $ **FLOATING
C3465 out_p.n1554 vss 4.56fF $ **FLOATING
C3466 out_p.n1555 vss 4.56fF $ **FLOATING
C3467 out_p.n1556 vss 4.56fF $ **FLOATING
C3468 out_p.n1557 vss 4.56fF $ **FLOATING
C3469 out_p.n1558 vss 4.56fF $ **FLOATING
C3470 out_p.n1559 vss 4.56fF $ **FLOATING
C3471 out_p.n1560 vss 4.56fF $ **FLOATING
C3472 out_p.n1561 vss 4.56fF $ **FLOATING
C3473 out_p.n1562 vss 4.56fF $ **FLOATING
C3474 out_p.n1563 vss 4.56fF $ **FLOATING
C3475 out_p.n1564 vss 4.27fF $ **FLOATING
C3476 out_p.n1565 vss 4.37fF $ **FLOATING
C3477 out_p.n1566 vss 4.53fF $ **FLOATING
C3478 out_p.n1567 vss 4.53fF $ **FLOATING
C3479 out_p.n1568 vss 4.26fF $ **FLOATING
C3480 out_p.n1569 vss 4.40fF $ **FLOATING
C3481 out_p.n1570 vss 4.56fF $ **FLOATING
C3482 out_p.n1571 vss 4.56fF $ **FLOATING
C3483 out_p.n1572 vss 4.56fF $ **FLOATING
C3484 out_p.n1573 vss 4.56fF $ **FLOATING
C3485 out_p.n1574 vss 4.56fF $ **FLOATING
C3486 out_p.n1575 vss 4.56fF $ **FLOATING
C3487 out_p.n1576 vss 4.56fF $ **FLOATING
C3488 out_p.n1577 vss 4.56fF $ **FLOATING
C3489 out_p.n1578 vss 4.56fF $ **FLOATING
C3490 out_p.n1579 vss 4.56fF $ **FLOATING
C3491 out_p.n1580 vss 4.56fF $ **FLOATING
C3492 out_p.n1581 vss 4.56fF $ **FLOATING
C3493 out_p.n1582 vss 4.56fF $ **FLOATING
C3494 out_p.n1583 vss 4.56fF $ **FLOATING
C3495 out_p.n1584 vss 4.56fF $ **FLOATING
C3496 out_p.n1585 vss 4.56fF $ **FLOATING
C3497 out_p.n1586 vss 4.56fF $ **FLOATING
C3498 out_p.n1587 vss 4.56fF $ **FLOATING
C3499 out_p.n1588 vss 4.27fF $ **FLOATING
C3500 out_p.n1589 vss 4.37fF $ **FLOATING
C3501 out_p.n1590 vss 4.53fF $ **FLOATING
C3502 out_p.n1591 vss 4.53fF $ **FLOATING
C3503 out_p.n1592 vss 4.26fF $ **FLOATING
C3504 out_p.n1593 vss 4.40fF $ **FLOATING
C3505 out_p.n1594 vss 4.56fF $ **FLOATING
C3506 out_p.n1595 vss 4.56fF $ **FLOATING
C3507 out_p.n1596 vss 4.56fF $ **FLOATING
C3508 out_p.n1597 vss 4.56fF $ **FLOATING
C3509 out_p.n1598 vss 4.56fF $ **FLOATING
C3510 out_p.n1599 vss 4.56fF $ **FLOATING
C3511 out_p.n1600 vss 4.56fF $ **FLOATING
C3512 out_p.n1601 vss 4.56fF $ **FLOATING
C3513 out_p.n1602 vss 4.56fF $ **FLOATING
C3514 out_p.n1603 vss 4.56fF $ **FLOATING
C3515 out_p.n1604 vss 4.56fF $ **FLOATING
C3516 out_p.n1605 vss 4.56fF $ **FLOATING
C3517 out_p.n1606 vss 4.56fF $ **FLOATING
C3518 out_p.n1607 vss 4.56fF $ **FLOATING
C3519 out_p.n1608 vss 4.56fF $ **FLOATING
C3520 out_p.n1609 vss 4.56fF $ **FLOATING
C3521 out_p.n1610 vss 4.56fF $ **FLOATING
C3522 out_p.n1611 vss 4.56fF $ **FLOATING
C3523 out_p.n1612 vss 4.27fF $ **FLOATING
C3524 out_p.n1613 vss 4.37fF $ **FLOATING
C3525 out_p.n1614 vss 4.53fF $ **FLOATING
C3526 out_p.n1615 vss 4.53fF $ **FLOATING
C3527 out_p.n1616 vss 4.26fF $ **FLOATING
C3528 out_p.n1617 vss 4.40fF $ **FLOATING
C3529 out_p.n1618 vss 4.56fF $ **FLOATING
C3530 out_p.n1619 vss 4.56fF $ **FLOATING
C3531 out_p.n1620 vss 4.56fF $ **FLOATING
C3532 out_p.n1621 vss 4.56fF $ **FLOATING
C3533 out_p.n1622 vss 4.56fF $ **FLOATING
C3534 out_p.n1623 vss 4.56fF $ **FLOATING
C3535 out_p.n1624 vss 4.56fF $ **FLOATING
C3536 out_p.n1625 vss 4.56fF $ **FLOATING
C3537 out_p.n1626 vss 4.56fF $ **FLOATING
C3538 out_p.n1627 vss 4.56fF $ **FLOATING
C3539 out_p.n1628 vss 4.56fF $ **FLOATING
C3540 out_p.n1629 vss 4.56fF $ **FLOATING
C3541 out_p.n1630 vss 4.56fF $ **FLOATING
C3542 out_p.n1631 vss 4.56fF $ **FLOATING
C3543 out_p.n1632 vss 4.56fF $ **FLOATING
C3544 out_p.n1633 vss 4.56fF $ **FLOATING
C3545 out_p.n1634 vss 4.56fF $ **FLOATING
C3546 out_p.n1635 vss 4.56fF $ **FLOATING
C3547 out_p.n1636 vss 4.27fF $ **FLOATING
C3548 out_p.n1637 vss 4.37fF $ **FLOATING
C3549 out_p.n1638 vss 4.53fF $ **FLOATING
C3550 out_p.n1639 vss 4.53fF $ **FLOATING
C3551 out_p.n1640 vss 4.26fF $ **FLOATING
C3552 out_p.n1641 vss 4.40fF $ **FLOATING
C3553 out_p.n1642 vss 4.56fF $ **FLOATING
C3554 out_p.n1643 vss 4.56fF $ **FLOATING
C3555 out_p.n1644 vss 4.56fF $ **FLOATING
C3556 out_p.n1645 vss 4.56fF $ **FLOATING
C3557 out_p.n1646 vss 4.56fF $ **FLOATING
C3558 out_p.n1647 vss 4.56fF $ **FLOATING
C3559 out_p.n1648 vss 4.56fF $ **FLOATING
C3560 out_p.n1649 vss 4.56fF $ **FLOATING
C3561 out_p.n1650 vss 4.56fF $ **FLOATING
C3562 out_p.n1651 vss 4.56fF $ **FLOATING
C3563 out_p.n1652 vss 4.56fF $ **FLOATING
C3564 out_p.n1653 vss 4.56fF $ **FLOATING
C3565 out_p.n1654 vss 4.56fF $ **FLOATING
C3566 out_p.n1655 vss 4.56fF $ **FLOATING
C3567 out_p.n1656 vss 4.56fF $ **FLOATING
C3568 out_p.n1657 vss 4.56fF $ **FLOATING
C3569 out_p.n1658 vss 4.56fF $ **FLOATING
C3570 out_p.n1659 vss 4.56fF $ **FLOATING
C3571 out_p.n1660 vss 4.27fF $ **FLOATING
C3572 out_p.n1661 vss 4.37fF $ **FLOATING
C3573 out_p.n1662 vss 4.53fF $ **FLOATING
C3574 out_p.n1663 vss 4.53fF $ **FLOATING
C3575 out_p.n1664 vss 4.26fF $ **FLOATING
C3576 out_p.n1665 vss 4.40fF $ **FLOATING
C3577 out_p.n1666 vss 4.56fF $ **FLOATING
C3578 out_p.n1667 vss 4.56fF $ **FLOATING
C3579 out_p.n1668 vss 4.56fF $ **FLOATING
C3580 out_p.n1669 vss 4.56fF $ **FLOATING
C3581 out_p.n1670 vss 4.56fF $ **FLOATING
C3582 out_p.n1671 vss 4.56fF $ **FLOATING
C3583 out_p.n1672 vss 4.56fF $ **FLOATING
C3584 out_p.n1673 vss 4.56fF $ **FLOATING
C3585 out_p.n1674 vss 4.56fF $ **FLOATING
C3586 out_p.n1675 vss 4.56fF $ **FLOATING
C3587 out_p.n1676 vss 4.56fF $ **FLOATING
C3588 out_p.n1677 vss 4.56fF $ **FLOATING
C3589 out_p.n1678 vss 4.56fF $ **FLOATING
C3590 out_p.n1679 vss 4.56fF $ **FLOATING
C3591 out_p.n1680 vss 4.56fF $ **FLOATING
C3592 out_p.n1681 vss 4.56fF $ **FLOATING
C3593 out_p.n1682 vss 4.56fF $ **FLOATING
C3594 out_p.n1683 vss 4.56fF $ **FLOATING
C3595 out_p.n1684 vss 4.27fF $ **FLOATING
C3596 out_p.n1685 vss 4.37fF $ **FLOATING
C3597 out_p.n1686 vss 4.53fF $ **FLOATING
C3598 out_p.n1687 vss 4.53fF $ **FLOATING
C3599 out_p.n1688 vss 4.26fF $ **FLOATING
C3600 out_p.n1689 vss 4.40fF $ **FLOATING
C3601 out_p.n1690 vss 4.56fF $ **FLOATING
C3602 out_p.n1691 vss 4.56fF $ **FLOATING
C3603 out_p.n1692 vss 4.56fF $ **FLOATING
C3604 out_p.n1693 vss 4.56fF $ **FLOATING
C3605 out_p.n1694 vss 4.56fF $ **FLOATING
C3606 out_p.n1695 vss 4.56fF $ **FLOATING
C3607 out_p.n1696 vss 4.56fF $ **FLOATING
C3608 out_p.n1697 vss 4.56fF $ **FLOATING
C3609 out_p.n1698 vss 4.56fF $ **FLOATING
C3610 out_p.n1699 vss 4.56fF $ **FLOATING
C3611 out_p.n1700 vss 4.56fF $ **FLOATING
C3612 out_p.n1701 vss 4.56fF $ **FLOATING
C3613 out_p.n1702 vss 4.56fF $ **FLOATING
C3614 out_p.n1703 vss 4.56fF $ **FLOATING
C3615 out_p.n1704 vss 4.56fF $ **FLOATING
C3616 out_p.n1705 vss 4.56fF $ **FLOATING
C3617 out_p.n1706 vss 4.56fF $ **FLOATING
C3618 out_p.n1707 vss 4.56fF $ **FLOATING
C3619 out_p.n1708 vss 4.27fF $ **FLOATING
C3620 out_p.n1709 vss 4.37fF $ **FLOATING
C3621 out_p.n1710 vss 4.53fF $ **FLOATING
C3622 out_p.n1711 vss 4.53fF $ **FLOATING
C3623 out_p.n1712 vss 4.26fF $ **FLOATING
C3624 out_p.n1713 vss 4.40fF $ **FLOATING
C3625 out_p.n1714 vss 4.56fF $ **FLOATING
C3626 out_p.n1715 vss 4.56fF $ **FLOATING
C3627 out_p.n1716 vss 4.56fF $ **FLOATING
C3628 out_p.n1717 vss 4.56fF $ **FLOATING
C3629 out_p.n1718 vss 4.56fF $ **FLOATING
C3630 out_p.n1719 vss 4.56fF $ **FLOATING
C3631 out_p.n1720 vss 4.56fF $ **FLOATING
C3632 out_p.n1721 vss 4.56fF $ **FLOATING
C3633 out_p.n1722 vss 4.56fF $ **FLOATING
C3634 out_p.n1723 vss 4.56fF $ **FLOATING
C3635 out_p.n1724 vss 4.56fF $ **FLOATING
C3636 out_p.n1725 vss 4.56fF $ **FLOATING
C3637 out_p.n1726 vss 4.56fF $ **FLOATING
C3638 out_p.n1727 vss 4.56fF $ **FLOATING
C3639 out_p.n1728 vss 4.56fF $ **FLOATING
C3640 out_p.n1729 vss 4.56fF $ **FLOATING
C3641 out_p.n1730 vss 4.56fF $ **FLOATING
C3642 out_p.n1731 vss 4.56fF $ **FLOATING
C3643 out_p.n1732 vss 4.27fF $ **FLOATING
C3644 out_p.n1733 vss 4.37fF $ **FLOATING
C3645 out_p.n1734 vss 4.53fF $ **FLOATING
C3646 out_p.n1735 vss 4.53fF $ **FLOATING
C3647 out_p.n1736 vss 4.26fF $ **FLOATING
C3648 out_p.n1737 vss 4.40fF $ **FLOATING
C3649 out_p.n1738 vss 4.56fF $ **FLOATING
C3650 out_p.n1739 vss 4.56fF $ **FLOATING
C3651 out_p.n1740 vss 4.56fF $ **FLOATING
C3652 out_p.n1741 vss 4.56fF $ **FLOATING
C3653 out_p.n1742 vss 4.56fF $ **FLOATING
C3654 out_p.n1743 vss 4.56fF $ **FLOATING
C3655 out_p.n1744 vss 4.56fF $ **FLOATING
C3656 out_p.n1745 vss 4.56fF $ **FLOATING
C3657 out_p.n1746 vss 4.56fF $ **FLOATING
C3658 out_p.n1747 vss 4.56fF $ **FLOATING
C3659 out_p.n1748 vss 4.56fF $ **FLOATING
C3660 out_p.n1749 vss 4.56fF $ **FLOATING
C3661 out_p.n1750 vss 4.56fF $ **FLOATING
C3662 out_p.n1751 vss 4.56fF $ **FLOATING
C3663 out_p.n1752 vss 4.56fF $ **FLOATING
C3664 out_p.n1753 vss 4.56fF $ **FLOATING
C3665 out_p.n1754 vss 4.56fF $ **FLOATING
C3666 out_p.n1755 vss 4.56fF $ **FLOATING
C3667 out_p.n1756 vss 4.27fF $ **FLOATING
C3668 out_p.n1757 vss 4.37fF $ **FLOATING
C3669 out_p.n1758 vss 4.53fF $ **FLOATING
C3670 out_p.n1759 vss 4.53fF $ **FLOATING
C3671 out_p.n1760 vss 4.26fF $ **FLOATING
C3672 out_p.n1761 vss 4.40fF $ **FLOATING
C3673 out_p.n1762 vss 4.56fF $ **FLOATING
C3674 out_p.n1763 vss 4.56fF $ **FLOATING
C3675 out_p.n1764 vss 4.56fF $ **FLOATING
C3676 out_p.n1765 vss 4.56fF $ **FLOATING
C3677 out_p.n1766 vss 4.56fF $ **FLOATING
C3678 out_p.n1767 vss 4.56fF $ **FLOATING
C3679 out_p.n1768 vss 4.56fF $ **FLOATING
C3680 out_p.n1769 vss 4.56fF $ **FLOATING
C3681 out_p.n1770 vss 4.56fF $ **FLOATING
C3682 out_p.n1771 vss 4.56fF $ **FLOATING
C3683 out_p.n1772 vss 4.56fF $ **FLOATING
C3684 out_p.n1773 vss 4.56fF $ **FLOATING
C3685 out_p.n1774 vss 4.56fF $ **FLOATING
C3686 out_p.n1775 vss 4.56fF $ **FLOATING
C3687 out_p.n1776 vss 4.56fF $ **FLOATING
C3688 out_p.n1777 vss 4.56fF $ **FLOATING
C3689 out_p.n1778 vss 4.56fF $ **FLOATING
C3690 out_p.n1779 vss 4.56fF $ **FLOATING
C3691 out_p.n1780 vss 4.27fF $ **FLOATING
C3692 out_p.n1781 vss 4.37fF $ **FLOATING
C3693 out_p.n1782 vss 4.53fF $ **FLOATING
C3694 out_p.n1783 vss 4.53fF $ **FLOATING
C3695 out_p.n1784 vss 4.26fF $ **FLOATING
C3696 out_p.n1785 vss 4.40fF $ **FLOATING
C3697 out_p.n1786 vss 4.56fF $ **FLOATING
C3698 out_p.n1787 vss 4.56fF $ **FLOATING
C3699 out_p.n1788 vss 4.56fF $ **FLOATING
C3700 out_p.n1789 vss 4.56fF $ **FLOATING
C3701 out_p.n1790 vss 4.56fF $ **FLOATING
C3702 out_p.n1791 vss 4.56fF $ **FLOATING
C3703 out_p.n1792 vss 4.56fF $ **FLOATING
C3704 out_p.n1793 vss 4.56fF $ **FLOATING
C3705 out_p.n1794 vss 4.56fF $ **FLOATING
C3706 out_p.n1795 vss 4.56fF $ **FLOATING
C3707 out_p.n1796 vss 4.56fF $ **FLOATING
C3708 out_p.n1797 vss 4.56fF $ **FLOATING
C3709 out_p.n1798 vss 4.56fF $ **FLOATING
C3710 out_p.n1799 vss 4.56fF $ **FLOATING
C3711 out_p.n1800 vss 4.56fF $ **FLOATING
C3712 out_p.n1801 vss 4.56fF $ **FLOATING
C3713 out_p.n1802 vss 4.56fF $ **FLOATING
C3714 out_p.n1803 vss 4.56fF $ **FLOATING
C3715 out_p.n1804 vss 4.27fF $ **FLOATING
C3716 out_p.n1805 vss 4.37fF $ **FLOATING
C3717 out_p.n1806 vss 4.53fF $ **FLOATING
C3718 out_p.n1807 vss 4.53fF $ **FLOATING
C3719 out_p.n1808 vss 4.26fF $ **FLOATING
C3720 out_p.n1809 vss 4.40fF $ **FLOATING
C3721 out_p.n1810 vss 4.56fF $ **FLOATING
C3722 out_p.n1811 vss 4.56fF $ **FLOATING
C3723 out_p.n1812 vss 4.56fF $ **FLOATING
C3724 out_p.n1813 vss 4.56fF $ **FLOATING
C3725 out_p.n1814 vss 4.56fF $ **FLOATING
C3726 out_p.n1815 vss 4.56fF $ **FLOATING
C3727 out_p.n1816 vss 4.56fF $ **FLOATING
C3728 out_p.n1817 vss 4.56fF $ **FLOATING
C3729 out_p.n1818 vss 4.56fF $ **FLOATING
C3730 out_p.n1819 vss 4.56fF $ **FLOATING
C3731 out_p.n1820 vss 4.56fF $ **FLOATING
C3732 out_p.n1821 vss 4.56fF $ **FLOATING
C3733 out_p.n1822 vss 4.56fF $ **FLOATING
C3734 out_p.n1823 vss 4.56fF $ **FLOATING
C3735 out_p.n1824 vss 4.56fF $ **FLOATING
C3736 out_p.n1825 vss 4.56fF $ **FLOATING
C3737 out_p.n1826 vss 4.56fF $ **FLOATING
C3738 out_p.n1827 vss 4.56fF $ **FLOATING
C3739 out_p.n1828 vss 4.27fF $ **FLOATING
C3740 out_p.n1829 vss 4.37fF $ **FLOATING
C3741 out_p.n1830 vss 4.53fF $ **FLOATING
C3742 out_p.n1831 vss 4.53fF $ **FLOATING
C3743 out_p.n1832 vss 4.26fF $ **FLOATING
C3744 out_p.n1833 vss 59.59fF $ **FLOATING
C3745 out_p.n1834 vss 85.93fF $ **FLOATING
C3746 out_p.n1835 vss 85.93fF $ **FLOATING
C3747 out_p.n1836 vss 85.93fF $ **FLOATING
C3748 out_p.n1837 vss 85.93fF $ **FLOATING
C3749 out_p.n1838 vss 85.93fF $ **FLOATING
C3750 out_p.n1839 vss 85.93fF $ **FLOATING
C3751 out_p.n1840 vss 85.93fF $ **FLOATING
C3752 out_p.n1841 vss 85.93fF $ **FLOATING
C3753 out_p.n1842 vss 85.93fF $ **FLOATING
C3754 out_p.n1843 vss 85.93fF $ **FLOATING
C3755 out_p.n1844 vss 85.93fF $ **FLOATING
C3756 out_p.n1845 vss 85.93fF $ **FLOATING
C3757 out_p.n1846 vss 85.93fF $ **FLOATING
C3758 out_p.n1847 vss 85.93fF $ **FLOATING
C3759 out_p.n1848 vss 85.93fF $ **FLOATING
C3760 out_p.n1849 vss 85.93fF $ **FLOATING
C3761 out_p.n1850 vss 85.93fF $ **FLOATING
C3762 out_p.n1851 vss 85.93fF $ **FLOATING
C3763 out_p.n1852 vss 85.93fF $ **FLOATING
C3764 out_p.n1853 vss 85.93fF $ **FLOATING
C3765 out_p.n1854 vss 85.93fF $ **FLOATING
C3766 out_p.n1855 vss 85.93fF $ **FLOATING
C3767 out_p.n1856 vss 85.93fF $ **FLOATING
C3768 out_p.n1857 vss 85.93fF $ **FLOATING
C3769 out_p.n1858 vss 85.93fF $ **FLOATING
C3770 out_p.n1859 vss 85.93fF $ **FLOATING
C3771 out_p.n1860 vss 85.93fF $ **FLOATING
C3772 out_p.n1861 vss 85.93fF $ **FLOATING
C3773 out_p.n1862 vss 85.93fF $ **FLOATING
C3774 out_p.n1863 vss 85.93fF $ **FLOATING
C3775 out_p.n1864 vss 85.93fF $ **FLOATING
C3776 out_p.n1865 vss 85.93fF $ **FLOATING
C3777 out_p.n1866 vss 85.93fF $ **FLOATING
C3778 out_p.n1867 vss 85.93fF $ **FLOATING
C3779 out_p.n1868 vss 85.93fF $ **FLOATING
C3780 out_p.n1869 vss 85.93fF $ **FLOATING
C3781 out_p.n1870 vss 85.93fF $ **FLOATING
C3782 out_p.n1871 vss 85.93fF $ **FLOATING
C3783 out_p.n1872 vss 85.93fF $ **FLOATING
C3784 out_p.n1873 vss 85.93fF $ **FLOATING
C3785 out_p.n1874 vss 74.13fF $ **FLOATING
C3786 vp_p.n451 vss 1.47fF $ **FLOATING
C3787 vp_p.n452 vss 15.99fF $ **FLOATING
C3788 vp_p.n453 vss 11.54fF $ **FLOATING
C3789 vp_p.n454 vss 11.54fF $ **FLOATING
C3790 vp_p.n455 vss 11.54fF $ **FLOATING
C3791 vp_p.n456 vss 11.54fF $ **FLOATING
C3792 vp_p.n457 vss 11.54fF $ **FLOATING
C3793 vp_p.n8727 vss 1.61fF $ **FLOATING
C3794 vp_p.n8728 vss 14.82fF $ **FLOATING
C3795 vp_p.n8729 vss 10.85fF $ **FLOATING
C3796 vp_p.n8730 vss 10.85fF $ **FLOATING
C3797 vp_p.n8731 vss 10.85fF $ **FLOATING
C3798 vp_p.n8732 vss 10.85fF $ **FLOATING
C3799 vp_p.n8733 vss 7.18fF $ **FLOATING
C3800 vp_p.n9190 vss 1.47fF $ **FLOATING
C3801 vp_p.n9191 vss 15.99fF $ **FLOATING
C3802 vp_p.n9192 vss 11.54fF $ **FLOATING
C3803 vp_p.n9193 vss 11.54fF $ **FLOATING
C3804 vp_p.n9194 vss 11.54fF $ **FLOATING
C3805 vp_p.n9195 vss 11.54fF $ **FLOATING
C3806 vp_p.n9196 vss 11.54fF $ **FLOATING
C3807 vp_p.n9197 vss 11.54fF $ **FLOATING
C3808 vp_p.n9198 vss 11.54fF $ **FLOATING
C3809 vp_p.n9199 vss 11.54fF $ **FLOATING
C3810 vp_p.n9200 vss 11.54fF $ **FLOATING
C3811 vp_p.n9201 vss 11.54fF $ **FLOATING
C3812 vp_p.n9202 vss 11.54fF $ **FLOATING
C3813 vp_p.n9203 vss 11.54fF $ **FLOATING
C3814 vp_p.n27425 vss 1.61fF $ **FLOATING
C3815 vp_p.n27426 vss 14.82fF $ **FLOATING
C3816 vp_p.n27427 vss 10.85fF $ **FLOATING
C3817 vp_p.n27428 vss 10.85fF $ **FLOATING
C3818 vp_p.n27429 vss 10.85fF $ **FLOATING
C3819 vp_p.n27430 vss 10.85fF $ **FLOATING
C3820 vp_p.n27431 vss 10.85fF $ **FLOATING
C3821 vp_p.n27432 vss 10.85fF $ **FLOATING
C3822 vp_p.n27433 vss 10.85fF $ **FLOATING
C3823 vp_p.n27434 vss 10.85fF $ **FLOATING
C3824 vp_p.n27435 vss 10.85fF $ **FLOATING
C3825 vp_p.n27436 vss 10.85fF $ **FLOATING
C3826 vp_p.n27437 vss 10.85fF $ **FLOATING
C3827 vp_p.n27438 vss 9.30fF $ **FLOATING
.ends
